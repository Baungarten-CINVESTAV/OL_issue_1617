magic
tech sky130A
magscale 1 2
timestamp 1674175363
<< viali >>
rect 14565 37349 14599 37383
rect 2053 37281 2087 37315
rect 3985 37281 4019 37315
rect 9137 37281 9171 37315
rect 12633 37281 12667 37315
rect 22661 37281 22695 37315
rect 37473 37281 37507 37315
rect 2329 37213 2363 37247
rect 4261 37213 4295 37247
rect 5457 37213 5491 37247
rect 6745 37213 6779 37247
rect 7389 37213 7423 37247
rect 9413 37213 9447 37247
rect 10425 37213 10459 37247
rect 11897 37213 11931 37247
rect 12449 37213 12483 37247
rect 14381 37213 14415 37247
rect 15209 37213 15243 37247
rect 16037 37213 16071 37247
rect 16865 37213 16899 37247
rect 18337 37213 18371 37247
rect 20085 37213 20119 37247
rect 21189 37213 21223 37247
rect 22937 37213 22971 37247
rect 24777 37213 24811 37247
rect 26065 37213 26099 37247
rect 27169 37213 27203 37247
rect 28089 37213 28123 37247
rect 29929 37213 29963 37247
rect 30573 37213 30607 37247
rect 31033 37213 31067 37247
rect 32505 37213 32539 37247
rect 32965 37213 32999 37247
rect 34897 37213 34931 37247
rect 36185 37213 36219 37247
rect 37749 37213 37783 37247
rect 5273 37077 5307 37111
rect 6561 37077 6595 37111
rect 7205 37077 7239 37111
rect 10609 37077 10643 37111
rect 11713 37077 11747 37111
rect 15025 37077 15059 37111
rect 16221 37077 16255 37111
rect 17049 37077 17083 37111
rect 18153 37077 18187 37111
rect 20269 37077 20303 37111
rect 21373 37077 21407 37111
rect 24593 37077 24627 37111
rect 25881 37077 25915 37111
rect 27353 37077 27387 37111
rect 27905 37077 27939 37111
rect 29745 37077 29779 37111
rect 30389 37077 30423 37111
rect 31217 37077 31251 37111
rect 32321 37077 32355 37111
rect 33149 37077 33183 37111
rect 35081 37077 35115 37111
rect 36369 37077 36403 37111
rect 10425 36873 10459 36907
rect 19625 36873 19659 36907
rect 23489 36873 23523 36907
rect 27169 36873 27203 36907
rect 36093 36873 36127 36907
rect 36829 36873 36863 36907
rect 37657 36873 37691 36907
rect 1685 36805 1719 36839
rect 2881 36737 2915 36771
rect 3525 36737 3559 36771
rect 9321 36737 9355 36771
rect 10609 36737 10643 36771
rect 19441 36737 19475 36771
rect 23305 36737 23339 36771
rect 27353 36737 27387 36771
rect 35449 36737 35483 36771
rect 35909 36737 35943 36771
rect 36645 36737 36679 36771
rect 37473 36737 37507 36771
rect 38025 36737 38059 36771
rect 1869 36601 1903 36635
rect 2697 36533 2731 36567
rect 3341 36533 3375 36567
rect 9137 36533 9171 36567
rect 35265 36533 35299 36567
rect 1777 36329 1811 36363
rect 36645 36329 36679 36363
rect 1593 36125 1627 36159
rect 2513 36125 2547 36159
rect 36829 36125 36863 36159
rect 37381 36125 37415 36159
rect 38025 36125 38059 36159
rect 2329 35989 2363 36023
rect 37473 35989 37507 36023
rect 38209 35989 38243 36023
rect 35541 35785 35575 35819
rect 1777 35649 1811 35683
rect 35449 35649 35483 35683
rect 38025 35649 38059 35683
rect 1593 35445 1627 35479
rect 38209 35445 38243 35479
rect 14749 35241 14783 35275
rect 14933 35037 14967 35071
rect 1593 34561 1627 34595
rect 6561 34561 6595 34595
rect 38025 34561 38059 34595
rect 6653 34493 6687 34527
rect 1777 34357 1811 34391
rect 38209 34357 38243 34391
rect 22109 33609 22143 33643
rect 15393 33473 15427 33507
rect 22293 33473 22327 33507
rect 15485 33269 15519 33303
rect 32137 33065 32171 33099
rect 1593 32861 1627 32895
rect 2513 32861 2547 32895
rect 32321 32861 32355 32895
rect 37473 32861 37507 32895
rect 37749 32861 37783 32895
rect 1777 32725 1811 32759
rect 2329 32725 2363 32759
rect 29653 32521 29687 32555
rect 1593 32385 1627 32419
rect 29837 32385 29871 32419
rect 38301 32385 38335 32419
rect 1777 32181 1811 32215
rect 38117 32181 38151 32215
rect 22293 31977 22327 32011
rect 27997 31977 28031 32011
rect 31125 31977 31159 32011
rect 36921 31977 36955 32011
rect 25789 31841 25823 31875
rect 27445 31841 27479 31875
rect 7941 31773 7975 31807
rect 8033 31773 8067 31807
rect 22477 31773 22511 31807
rect 25697 31773 25731 31807
rect 27353 31773 27387 31807
rect 28181 31773 28215 31807
rect 31033 31773 31067 31807
rect 37105 31773 37139 31807
rect 32505 31433 32539 31467
rect 6561 31297 6595 31331
rect 7205 31297 7239 31331
rect 16865 31297 16899 31331
rect 32689 31297 32723 31331
rect 6653 31093 6687 31127
rect 7297 31093 7331 31127
rect 16957 31093 16991 31127
rect 3985 30889 4019 30923
rect 36277 30889 36311 30923
rect 1593 30685 1627 30719
rect 4169 30685 4203 30719
rect 10425 30685 10459 30719
rect 21833 30685 21867 30719
rect 22661 30685 22695 30719
rect 27997 30685 28031 30719
rect 36185 30685 36219 30719
rect 38301 30685 38335 30719
rect 22753 30617 22787 30651
rect 1777 30549 1811 30583
rect 10517 30549 10551 30583
rect 21925 30549 21959 30583
rect 28089 30549 28123 30583
rect 38117 30549 38151 30583
rect 13921 30277 13955 30311
rect 29653 30277 29687 30311
rect 6561 30209 6595 30243
rect 13829 30209 13863 30243
rect 14473 30209 14507 30243
rect 23397 30209 23431 30243
rect 26249 30209 26283 30243
rect 29561 30209 29595 30243
rect 38025 30209 38059 30243
rect 26341 30073 26375 30107
rect 37841 30073 37875 30107
rect 6653 30005 6687 30039
rect 14565 30005 14599 30039
rect 23489 30005 23523 30039
rect 21557 29801 21591 29835
rect 29837 29801 29871 29835
rect 1593 29597 1627 29631
rect 11437 29597 11471 29631
rect 21465 29597 21499 29631
rect 29745 29597 29779 29631
rect 38117 29529 38151 29563
rect 1777 29461 1811 29495
rect 11529 29461 11563 29495
rect 38209 29461 38243 29495
rect 22017 29257 22051 29291
rect 1777 29121 1811 29155
rect 11989 29121 12023 29155
rect 22201 29121 22235 29155
rect 38301 29121 38335 29155
rect 1593 28985 1627 29019
rect 12081 28985 12115 29019
rect 38117 28985 38151 29019
rect 6285 28713 6319 28747
rect 6469 28509 6503 28543
rect 11713 28509 11747 28543
rect 27537 28509 27571 28543
rect 11529 28373 11563 28407
rect 27629 28373 27663 28407
rect 10333 28169 10367 28203
rect 9137 28033 9171 28067
rect 10517 28033 10551 28067
rect 11161 28033 11195 28067
rect 11805 28033 11839 28067
rect 12633 28033 12667 28067
rect 13461 28033 13495 28067
rect 10977 27897 11011 27931
rect 9229 27829 9263 27863
rect 11897 27829 11931 27863
rect 12725 27829 12759 27863
rect 13277 27829 13311 27863
rect 10425 27557 10459 27591
rect 13461 27557 13495 27591
rect 11897 27489 11931 27523
rect 13001 27489 13035 27523
rect 1593 27421 1627 27455
rect 1869 27421 1903 27455
rect 10609 27421 10643 27455
rect 11069 27421 11103 27455
rect 11161 27421 11195 27455
rect 11713 27421 11747 27455
rect 12357 27421 12391 27455
rect 12817 27421 12851 27455
rect 38301 27421 38335 27455
rect 14749 27285 14783 27319
rect 38117 27285 38151 27319
rect 12449 27081 12483 27115
rect 13553 27081 13587 27115
rect 22477 27081 22511 27115
rect 10977 27013 11011 27047
rect 10425 26945 10459 26979
rect 11989 26945 12023 26979
rect 13093 26945 13127 26979
rect 14749 26945 14783 26979
rect 15393 26945 15427 26979
rect 22661 26945 22695 26979
rect 23305 26945 23339 26979
rect 11805 26877 11839 26911
rect 12909 26877 12943 26911
rect 10241 26809 10275 26843
rect 11069 26741 11103 26775
rect 14565 26741 14599 26775
rect 15209 26741 15243 26775
rect 23121 26741 23155 26775
rect 9413 26537 9447 26571
rect 10057 26537 10091 26571
rect 13461 26537 13495 26571
rect 14657 26537 14691 26571
rect 21281 26537 21315 26571
rect 1869 26469 1903 26503
rect 38117 26469 38151 26503
rect 11989 26401 12023 26435
rect 13277 26401 13311 26435
rect 15485 26401 15519 26435
rect 16497 26401 16531 26435
rect 9321 26333 9355 26367
rect 10241 26333 10275 26367
rect 10701 26333 10735 26367
rect 11529 26333 11563 26367
rect 12173 26333 12207 26367
rect 13093 26333 13127 26367
rect 14841 26333 14875 26367
rect 15301 26333 15335 26367
rect 16405 26333 16439 26367
rect 20821 26333 20855 26367
rect 21465 26333 21499 26367
rect 22661 26333 22695 26367
rect 38301 26333 38335 26367
rect 1685 26265 1719 26299
rect 10793 26265 10827 26299
rect 11345 26197 11379 26231
rect 12633 26197 12667 26231
rect 15945 26197 15979 26231
rect 20637 26197 20671 26231
rect 22477 26197 22511 26231
rect 23121 26197 23155 26231
rect 14013 25993 14047 26027
rect 15301 25993 15335 26027
rect 20269 25993 20303 26027
rect 8401 25925 8435 25959
rect 12081 25925 12115 25959
rect 18429 25925 18463 25959
rect 18521 25925 18555 25959
rect 20177 25925 20211 25959
rect 8309 25857 8343 25891
rect 10517 25857 10551 25891
rect 14197 25857 14231 25891
rect 14657 25857 14691 25891
rect 14841 25857 14875 25891
rect 20821 25857 20855 25891
rect 22017 25857 22051 25891
rect 23121 25857 23155 25891
rect 23305 25857 23339 25891
rect 30389 25857 30423 25891
rect 11989 25789 12023 25823
rect 13001 25789 13035 25823
rect 19257 25789 19291 25823
rect 22201 25789 22235 25823
rect 10609 25653 10643 25687
rect 20913 25653 20947 25687
rect 22661 25653 22695 25687
rect 23765 25653 23799 25687
rect 30481 25653 30515 25687
rect 10793 25449 10827 25483
rect 12633 25449 12667 25483
rect 13461 25449 13495 25483
rect 19533 25449 19567 25483
rect 24685 25449 24719 25483
rect 6377 25381 6411 25415
rect 11989 25313 12023 25347
rect 13277 25313 13311 25347
rect 21189 25313 21223 25347
rect 21465 25313 21499 25347
rect 6285 25245 6319 25279
rect 10701 25245 10735 25279
rect 12173 25245 12207 25279
rect 13093 25245 13127 25279
rect 14289 25245 14323 25279
rect 15117 25245 15151 25279
rect 15761 25245 15795 25279
rect 16681 25245 16715 25279
rect 19441 25245 19475 25279
rect 23121 25245 23155 25279
rect 24593 25245 24627 25279
rect 31125 25245 31159 25279
rect 38025 25245 38059 25279
rect 11345 25177 11379 25211
rect 15853 25177 15887 25211
rect 21281 25177 21315 25211
rect 14381 25109 14415 25143
rect 15209 25109 15243 25143
rect 16773 25109 16807 25143
rect 22937 25109 22971 25143
rect 31217 25109 31251 25143
rect 38209 25109 38243 25143
rect 22109 24905 22143 24939
rect 24225 24905 24259 24939
rect 13185 24837 13219 24871
rect 14749 24837 14783 24871
rect 18061 24837 18095 24871
rect 22937 24837 22971 24871
rect 1593 24769 1627 24803
rect 10609 24769 10643 24803
rect 11713 24769 11747 24803
rect 11805 24769 11839 24803
rect 12357 24769 12391 24803
rect 16129 24769 16163 24803
rect 17233 24769 17267 24803
rect 17325 24769 17359 24803
rect 19625 24769 19659 24803
rect 22017 24769 22051 24803
rect 24409 24769 24443 24803
rect 25053 24769 25087 24803
rect 25789 24769 25823 24803
rect 25881 24769 25915 24803
rect 30665 24769 30699 24803
rect 13093 24701 13127 24735
rect 14105 24701 14139 24735
rect 14657 24701 14691 24735
rect 15301 24701 15335 24735
rect 16221 24701 16255 24735
rect 17969 24689 18003 24723
rect 18245 24701 18279 24735
rect 22845 24701 22879 24735
rect 23397 24633 23431 24667
rect 1777 24565 1811 24599
rect 10701 24565 10735 24599
rect 12449 24565 12483 24599
rect 19441 24565 19475 24599
rect 24869 24565 24903 24599
rect 30757 24565 30791 24599
rect 14749 24361 14783 24395
rect 17693 24293 17727 24327
rect 24961 24293 24995 24327
rect 12541 24225 12575 24259
rect 14565 24225 14599 24259
rect 22753 24225 22787 24259
rect 24593 24225 24627 24259
rect 24777 24225 24811 24259
rect 37749 24225 37783 24259
rect 1593 24157 1627 24191
rect 1869 24157 1903 24191
rect 14381 24157 14415 24191
rect 15577 24157 15611 24191
rect 16773 24157 16807 24191
rect 16865 24157 16899 24191
rect 18337 24157 18371 24191
rect 29745 24157 29779 24191
rect 37473 24157 37507 24191
rect 12633 24089 12667 24123
rect 13185 24089 13219 24123
rect 17509 24089 17543 24123
rect 22845 24089 22879 24123
rect 23765 24089 23799 24123
rect 15669 24021 15703 24055
rect 18429 24021 18463 24055
rect 20085 24021 20119 24055
rect 29837 24021 29871 24055
rect 19257 23817 19291 23851
rect 20729 23817 20763 23851
rect 30481 23817 30515 23851
rect 13001 23749 13035 23783
rect 15393 23749 15427 23783
rect 16957 23749 16991 23783
rect 22201 23749 22235 23783
rect 23397 23749 23431 23783
rect 2145 23681 2179 23715
rect 4721 23681 4755 23715
rect 10149 23681 10183 23715
rect 11897 23681 11931 23715
rect 14565 23681 14599 23715
rect 16865 23681 16899 23715
rect 17785 23681 17819 23715
rect 18613 23681 18647 23715
rect 18797 23681 18831 23715
rect 20085 23681 20119 23715
rect 20269 23681 20303 23715
rect 29745 23681 29779 23715
rect 30389 23681 30423 23715
rect 12909 23613 12943 23647
rect 15301 23613 15335 23647
rect 15577 23613 15611 23647
rect 22109 23613 22143 23647
rect 22385 23613 22419 23647
rect 23305 23613 23339 23647
rect 23581 23613 23615 23647
rect 4537 23545 4571 23579
rect 13461 23545 13495 23579
rect 1961 23477 1995 23511
rect 10241 23477 10275 23511
rect 11989 23477 12023 23511
rect 14657 23477 14691 23511
rect 17877 23477 17911 23511
rect 29837 23477 29871 23511
rect 17969 23273 18003 23307
rect 10241 23137 10275 23171
rect 11253 23137 11287 23171
rect 15025 23137 15059 23171
rect 16957 23137 16991 23171
rect 20177 23137 20211 23171
rect 21097 23137 21131 23171
rect 24777 23137 24811 23171
rect 12265 23069 12299 23103
rect 15853 23069 15887 23103
rect 16773 23069 16807 23103
rect 17877 23069 17911 23103
rect 10333 23001 10367 23035
rect 14749 23001 14783 23035
rect 14841 23001 14875 23035
rect 19901 23001 19935 23035
rect 19993 23001 20027 23035
rect 21189 23001 21223 23035
rect 22109 23001 22143 23035
rect 24869 23001 24903 23035
rect 25421 23001 25455 23035
rect 9505 22933 9539 22967
rect 12357 22933 12391 22967
rect 15945 22933 15979 22967
rect 17417 22933 17451 22967
rect 9045 22729 9079 22763
rect 11897 22729 11931 22763
rect 15209 22729 15243 22763
rect 20361 22729 20395 22763
rect 22109 22729 22143 22763
rect 25053 22729 25087 22763
rect 30757 22729 30791 22763
rect 7297 22661 7331 22695
rect 7849 22661 7883 22695
rect 9781 22661 9815 22695
rect 9873 22661 9907 22695
rect 13461 22661 13495 22695
rect 17233 22661 17267 22695
rect 27261 22661 27295 22695
rect 27353 22661 27387 22695
rect 1777 22593 1811 22627
rect 9229 22593 9263 22627
rect 10885 22593 10919 22627
rect 11805 22593 11839 22627
rect 14749 22593 14783 22627
rect 16129 22593 16163 22627
rect 18613 22593 18647 22627
rect 22017 22593 22051 22627
rect 24961 22593 24995 22627
rect 26157 22593 26191 22627
rect 30481 22593 30515 22627
rect 30941 22593 30975 22627
rect 38025 22593 38059 22627
rect 7205 22525 7239 22559
rect 10425 22525 10459 22559
rect 13369 22525 13403 22559
rect 13829 22525 13863 22559
rect 14565 22525 14599 22559
rect 17141 22525 17175 22559
rect 17969 22525 18003 22559
rect 27537 22525 27571 22559
rect 38209 22457 38243 22491
rect 1593 22389 1627 22423
rect 10977 22389 11011 22423
rect 16221 22389 16255 22423
rect 18705 22389 18739 22423
rect 26249 22389 26283 22423
rect 26341 22185 26375 22219
rect 27537 22117 27571 22151
rect 7021 22049 7055 22083
rect 11713 22049 11747 22083
rect 14381 22049 14415 22083
rect 17601 22049 17635 22083
rect 17969 22049 18003 22083
rect 6929 21981 6963 22015
rect 8033 21981 8067 22015
rect 9137 21981 9171 22015
rect 14289 21981 14323 22015
rect 15393 21981 15427 22015
rect 15853 21981 15887 22015
rect 16865 21981 16899 22015
rect 19533 21981 19567 22015
rect 24593 21981 24627 22015
rect 26249 21981 26283 22015
rect 34897 21981 34931 22015
rect 34989 21981 35023 22015
rect 37565 21981 37599 22015
rect 38025 21981 38059 22015
rect 9229 21913 9263 21947
rect 10057 21913 10091 21947
rect 10149 21913 10183 21947
rect 10701 21913 10735 21947
rect 11437 21913 11471 21947
rect 11529 21913 11563 21947
rect 15209 21913 15243 21947
rect 15945 21913 15979 21947
rect 17693 21913 17727 21947
rect 26985 21913 27019 21947
rect 27077 21913 27111 21947
rect 8125 21845 8159 21879
rect 16957 21845 16991 21879
rect 19625 21845 19659 21879
rect 24685 21845 24719 21879
rect 37381 21845 37415 21879
rect 38209 21845 38243 21879
rect 8585 21641 8619 21675
rect 22385 21641 22419 21675
rect 28273 21641 28307 21675
rect 5457 21573 5491 21607
rect 7389 21573 7423 21607
rect 7481 21573 7515 21607
rect 12817 21573 12851 21607
rect 14197 21573 14231 21607
rect 15393 21573 15427 21607
rect 16957 21573 16991 21607
rect 18429 21573 18463 21607
rect 18981 21573 19015 21607
rect 19625 21573 19659 21607
rect 23581 21573 23615 21607
rect 1685 21505 1719 21539
rect 6009 21505 6043 21539
rect 8493 21505 8527 21539
rect 9137 21505 9171 21539
rect 14105 21505 14139 21539
rect 17601 21505 17635 21539
rect 20637 21505 20671 21539
rect 22569 21505 22603 21539
rect 24777 21505 24811 21539
rect 28181 21505 28215 21539
rect 5365 21437 5399 21471
rect 12725 21437 12759 21471
rect 13369 21437 13403 21471
rect 15301 21437 15335 21471
rect 16313 21437 16347 21471
rect 18337 21437 18371 21471
rect 19533 21437 19567 21471
rect 23489 21437 23523 21471
rect 1869 21369 1903 21403
rect 7941 21369 7975 21403
rect 20085 21369 20119 21403
rect 24041 21369 24075 21403
rect 9229 21301 9263 21335
rect 17049 21301 17083 21335
rect 17693 21301 17727 21335
rect 20729 21301 20763 21335
rect 24593 21301 24627 21335
rect 37841 21097 37875 21131
rect 23765 21029 23799 21063
rect 4813 20961 4847 20995
rect 5641 20961 5675 20995
rect 10425 20961 10459 20995
rect 12265 20961 12299 20995
rect 13277 20961 13311 20995
rect 16589 20961 16623 20995
rect 16957 20961 16991 20995
rect 18889 20961 18923 20995
rect 19625 20961 19659 20995
rect 20361 20961 20395 20995
rect 23213 20961 23247 20995
rect 1593 20893 1627 20927
rect 1869 20893 1903 20927
rect 6285 20893 6319 20927
rect 8401 20893 8435 20927
rect 9137 20893 9171 20927
rect 21005 20893 21039 20927
rect 22477 20893 22511 20927
rect 22569 20893 22603 20927
rect 25237 20893 25271 20927
rect 38025 20893 38059 20927
rect 4537 20825 4571 20859
rect 4629 20825 4663 20859
rect 10149 20825 10183 20859
rect 10241 20825 10275 20859
rect 12357 20825 12391 20859
rect 14657 20825 14691 20859
rect 14749 20825 14783 20859
rect 15669 20825 15703 20859
rect 16681 20825 16715 20859
rect 18245 20825 18279 20859
rect 18337 20825 18371 20859
rect 20453 20825 20487 20859
rect 23305 20825 23339 20859
rect 6377 20757 6411 20791
rect 8493 20757 8527 20791
rect 9229 20757 9263 20791
rect 25053 20757 25087 20791
rect 7757 20553 7791 20587
rect 14381 20553 14415 20587
rect 26433 20553 26467 20587
rect 8401 20485 8435 20519
rect 8493 20485 8527 20519
rect 10333 20485 10367 20519
rect 10425 20485 10459 20519
rect 11897 20485 11931 20519
rect 13277 20485 13311 20519
rect 15393 20485 15427 20519
rect 17325 20485 17359 20519
rect 18429 20485 18463 20519
rect 19349 20485 19383 20519
rect 19441 20485 19475 20519
rect 22201 20485 22235 20519
rect 23397 20485 23431 20519
rect 7665 20417 7699 20451
rect 14289 20417 14323 20451
rect 18337 20417 18371 20451
rect 24409 20417 24443 20451
rect 24593 20417 24627 20451
rect 25789 20417 25823 20451
rect 27169 20417 27203 20451
rect 38301 20417 38335 20451
rect 9229 20349 9263 20383
rect 10977 20349 11011 20383
rect 11805 20349 11839 20383
rect 12081 20349 12115 20383
rect 13185 20349 13219 20383
rect 13461 20349 13495 20383
rect 15301 20349 15335 20383
rect 16313 20349 16347 20383
rect 17233 20349 17267 20383
rect 20177 20349 20211 20383
rect 22109 20349 22143 20383
rect 23305 20349 23339 20383
rect 25973 20349 26007 20383
rect 27261 20349 27295 20383
rect 17785 20281 17819 20315
rect 22661 20281 22695 20315
rect 23857 20281 23891 20315
rect 25053 20213 25087 20247
rect 38117 20213 38151 20247
rect 9229 20009 9263 20043
rect 10793 20009 10827 20043
rect 25697 20009 25731 20043
rect 6929 19941 6963 19975
rect 25145 19941 25179 19975
rect 5273 19873 5307 19907
rect 6377 19873 6411 19907
rect 14381 19873 14415 19907
rect 17601 19873 17635 19907
rect 19901 19873 19935 19907
rect 21281 19873 21315 19907
rect 22293 19873 22327 19907
rect 24593 19873 24627 19907
rect 9137 19805 9171 19839
rect 9781 19805 9815 19839
rect 10701 19805 10735 19839
rect 11529 19805 11563 19839
rect 16221 19805 16255 19839
rect 17049 19805 17083 19839
rect 19809 19805 19843 19839
rect 24777 19805 24811 19839
rect 25881 19805 25915 19839
rect 26341 19805 26375 19839
rect 26985 19805 27019 19839
rect 29929 19805 29963 19839
rect 4261 19737 4295 19771
rect 4353 19737 4387 19771
rect 6469 19737 6503 19771
rect 7573 19737 7607 19771
rect 7665 19737 7699 19771
rect 8585 19737 8619 19771
rect 12449 19737 12483 19771
rect 12541 19737 12575 19771
rect 13461 19737 13495 19771
rect 14473 19737 14507 19771
rect 15393 19737 15427 19771
rect 16313 19737 16347 19771
rect 17693 19737 17727 19771
rect 18613 19737 18647 19771
rect 21373 19737 21407 19771
rect 23397 19737 23431 19771
rect 9873 19669 9907 19703
rect 11621 19669 11655 19703
rect 16865 19669 16899 19703
rect 23489 19669 23523 19703
rect 26433 19669 26467 19703
rect 27077 19669 27111 19703
rect 29745 19669 29779 19703
rect 1777 19465 1811 19499
rect 5089 19465 5123 19499
rect 10425 19465 10459 19499
rect 14565 19465 14599 19499
rect 15301 19465 15335 19499
rect 16037 19465 16071 19499
rect 17877 19465 17911 19499
rect 20269 19465 20303 19499
rect 23029 19465 23063 19499
rect 23673 19465 23707 19499
rect 24685 19465 24719 19499
rect 25329 19465 25363 19499
rect 26525 19465 26559 19499
rect 28641 19465 28675 19499
rect 29929 19465 29963 19499
rect 6837 19397 6871 19431
rect 8401 19397 8435 19431
rect 9321 19397 9355 19431
rect 11069 19397 11103 19431
rect 13093 19397 13127 19431
rect 14013 19397 14047 19431
rect 1961 19329 1995 19363
rect 4997 19329 5031 19363
rect 5641 19329 5675 19363
rect 10333 19329 10367 19363
rect 10977 19329 11011 19363
rect 12265 19329 12299 19363
rect 14749 19329 14783 19363
rect 15209 19329 15243 19363
rect 15945 19329 15979 19363
rect 17233 19329 17267 19363
rect 17325 19329 17359 19363
rect 18061 19329 18095 19363
rect 19625 19329 19659 19363
rect 21281 19329 21315 19363
rect 21373 19329 21407 19363
rect 23213 19329 23247 19363
rect 23857 19329 23891 19363
rect 24593 19329 24627 19363
rect 25237 19329 25271 19363
rect 25881 19329 25915 19363
rect 27353 19329 27387 19363
rect 28825 19329 28859 19363
rect 29285 19329 29319 19363
rect 30113 19329 30147 19363
rect 38025 19329 38059 19363
rect 6745 19261 6779 19295
rect 7113 19261 7147 19295
rect 8309 19261 8343 19295
rect 13001 19261 13035 19295
rect 19809 19261 19843 19295
rect 26065 19261 26099 19295
rect 5733 19125 5767 19159
rect 12357 19125 12391 19159
rect 27169 19125 27203 19159
rect 29377 19125 29411 19159
rect 38209 19125 38243 19159
rect 7849 18921 7883 18955
rect 8493 18921 8527 18955
rect 11161 18921 11195 18955
rect 17233 18921 17267 18955
rect 20637 18921 20671 18955
rect 27353 18921 27387 18955
rect 34989 18921 35023 18955
rect 1593 18853 1627 18887
rect 11805 18853 11839 18887
rect 31585 18853 31619 18887
rect 12449 18785 12483 18819
rect 16037 18785 16071 18819
rect 16681 18785 16715 18819
rect 25605 18785 25639 18819
rect 26249 18785 26283 18819
rect 29101 18785 29135 18819
rect 29929 18785 29963 18819
rect 1777 18717 1811 18751
rect 5825 18717 5859 18751
rect 6469 18717 6503 18751
rect 7113 18717 7147 18751
rect 7757 18717 7791 18751
rect 8401 18717 8435 18751
rect 9137 18717 9171 18751
rect 9781 18717 9815 18751
rect 10425 18717 10459 18751
rect 11069 18717 11103 18751
rect 11713 18717 11747 18751
rect 17141 18717 17175 18751
rect 17969 18717 18003 18751
rect 20545 18717 20579 18751
rect 23857 18717 23891 18751
rect 27537 18717 27571 18751
rect 29009 18717 29043 18751
rect 29745 18717 29779 18751
rect 31493 18717 31527 18751
rect 33517 18717 33551 18751
rect 35173 18717 35207 18751
rect 9873 18649 9907 18683
rect 12541 18649 12575 18683
rect 13461 18649 13495 18683
rect 14749 18649 14783 18683
rect 14841 18649 14875 18683
rect 15393 18649 15427 18683
rect 16129 18649 16163 18683
rect 24685 18649 24719 18683
rect 24777 18649 24811 18683
rect 26341 18649 26375 18683
rect 26893 18649 26927 18683
rect 5917 18581 5951 18615
rect 6561 18581 6595 18615
rect 7205 18581 7239 18615
rect 9229 18581 9263 18615
rect 10517 18581 10551 18615
rect 17785 18581 17819 18615
rect 23949 18581 23983 18615
rect 30389 18581 30423 18615
rect 33609 18581 33643 18615
rect 13553 18377 13587 18411
rect 18153 18377 18187 18411
rect 18797 18377 18831 18411
rect 29561 18377 29595 18411
rect 30297 18377 30331 18411
rect 4261 18309 4295 18343
rect 4813 18309 4847 18343
rect 5457 18309 5491 18343
rect 6929 18309 6963 18343
rect 7021 18309 7055 18343
rect 11897 18309 11931 18343
rect 12817 18309 12851 18343
rect 14933 18309 14967 18343
rect 17049 18309 17083 18343
rect 19441 18309 19475 18343
rect 24685 18309 24719 18343
rect 24869 18309 24903 18343
rect 27813 18309 27847 18343
rect 27905 18309 27939 18343
rect 1869 18241 1903 18275
rect 8401 18241 8435 18275
rect 9045 18241 9079 18275
rect 9689 18241 9723 18275
rect 10333 18241 10367 18275
rect 11001 18241 11035 18275
rect 13461 18241 13495 18275
rect 14105 18241 14139 18275
rect 18061 18241 18095 18275
rect 18705 18241 18739 18275
rect 20545 18241 20579 18275
rect 20637 18241 20671 18275
rect 25513 18241 25547 18275
rect 28917 18241 28951 18275
rect 29745 18241 29779 18275
rect 30205 18241 30239 18275
rect 1593 18173 1627 18207
rect 4169 18173 4203 18207
rect 5365 18173 5399 18207
rect 6009 18173 6043 18207
rect 7941 18173 7975 18207
rect 10425 18173 10459 18207
rect 11805 18173 11839 18207
rect 14841 18173 14875 18207
rect 15393 18173 15427 18207
rect 16957 18173 16991 18207
rect 19625 18173 19659 18207
rect 25329 18173 25363 18207
rect 28089 18173 28123 18207
rect 8493 18105 8527 18139
rect 9781 18105 9815 18139
rect 11069 18105 11103 18139
rect 14197 18105 14231 18139
rect 17509 18105 17543 18139
rect 9137 18037 9171 18071
rect 25697 18037 25731 18071
rect 29009 18037 29043 18071
rect 4353 17833 4387 17867
rect 18521 17833 18555 17867
rect 21281 17833 21315 17867
rect 21925 17833 21959 17867
rect 9413 17765 9447 17799
rect 8493 17697 8527 17731
rect 11345 17697 11379 17731
rect 12357 17697 12391 17731
rect 15209 17697 15243 17731
rect 16773 17697 16807 17731
rect 17877 17697 17911 17731
rect 18061 17697 18095 17731
rect 25881 17697 25915 17731
rect 4261 17629 4295 17663
rect 4905 17629 4939 17663
rect 7757 17629 7791 17663
rect 8401 17629 8435 17663
rect 9321 17629 9355 17663
rect 9965 17629 9999 17663
rect 10609 17629 10643 17663
rect 12817 17629 12851 17663
rect 14473 17629 14507 17663
rect 20085 17629 20119 17663
rect 21189 17629 21223 17663
rect 21833 17629 21867 17663
rect 28549 17629 28583 17663
rect 10057 17561 10091 17595
rect 11437 17561 11471 17595
rect 13093 17561 13127 17595
rect 15301 17561 15335 17595
rect 15853 17561 15887 17595
rect 16405 17561 16439 17595
rect 16497 17561 16531 17595
rect 25973 17561 26007 17595
rect 26893 17561 26927 17595
rect 4997 17493 5031 17527
rect 7849 17493 7883 17527
rect 10701 17493 10735 17527
rect 14565 17493 14599 17527
rect 19441 17493 19475 17527
rect 20177 17493 20211 17527
rect 22477 17493 22511 17527
rect 27905 17493 27939 17527
rect 28641 17493 28675 17527
rect 7941 17289 7975 17323
rect 15209 17289 15243 17323
rect 16221 17289 16255 17323
rect 28825 17289 28859 17323
rect 4261 17221 4295 17255
rect 5181 17221 5215 17255
rect 10609 17221 10643 17255
rect 13185 17221 13219 17255
rect 14105 17221 14139 17255
rect 17141 17221 17175 17255
rect 18889 17221 18923 17255
rect 18981 17221 19015 17255
rect 20821 17221 20855 17255
rect 20913 17221 20947 17255
rect 22201 17221 22235 17255
rect 22293 17221 22327 17255
rect 23213 17221 23247 17255
rect 24225 17221 24259 17255
rect 1777 17153 1811 17187
rect 6561 17153 6595 17187
rect 7205 17153 7239 17187
rect 7849 17153 7883 17187
rect 8493 17153 8527 17187
rect 9137 17153 9171 17187
rect 9781 17153 9815 17187
rect 11897 17153 11931 17187
rect 15117 17153 15151 17187
rect 16129 17153 16163 17187
rect 19993 17153 20027 17187
rect 28181 17153 28215 17187
rect 28365 17153 28399 17187
rect 32965 17153 32999 17187
rect 38025 17153 38059 17187
rect 4169 17085 4203 17119
rect 6653 17085 6687 17119
rect 10517 17085 10551 17119
rect 12081 17085 12115 17119
rect 13093 17085 13127 17119
rect 17049 17085 17083 17119
rect 17877 17085 17911 17119
rect 19533 17085 19567 17119
rect 21097 17085 21131 17119
rect 24133 17085 24167 17119
rect 24409 17085 24443 17119
rect 29285 17085 29319 17119
rect 9229 17017 9263 17051
rect 11069 17017 11103 17051
rect 32781 17017 32815 17051
rect 38209 17017 38243 17051
rect 1593 16949 1627 16983
rect 7297 16949 7331 16983
rect 8585 16949 8619 16983
rect 9873 16949 9907 16983
rect 20085 16949 20119 16983
rect 17049 16745 17083 16779
rect 18613 16745 18647 16779
rect 23489 16745 23523 16779
rect 14933 16677 14967 16711
rect 7021 16609 7055 16643
rect 10241 16609 10275 16643
rect 10885 16609 10919 16643
rect 12633 16609 12667 16643
rect 28733 16609 28767 16643
rect 29837 16609 29871 16643
rect 30113 16609 30147 16643
rect 6285 16541 6319 16575
rect 11437 16541 11471 16575
rect 15485 16541 15519 16575
rect 16957 16541 16991 16575
rect 17601 16541 17635 16575
rect 18521 16541 18555 16575
rect 20177 16541 20211 16575
rect 21741 16541 21775 16575
rect 22477 16541 22511 16575
rect 22569 16541 22603 16575
rect 23397 16541 23431 16575
rect 24593 16541 24627 16575
rect 27537 16541 27571 16575
rect 7113 16473 7147 16507
rect 8033 16473 8067 16507
rect 10333 16473 10367 16507
rect 11805 16473 11839 16507
rect 12725 16473 12759 16507
rect 13645 16473 13679 16507
rect 14381 16473 14415 16507
rect 14473 16473 14507 16507
rect 15761 16473 15795 16507
rect 19533 16473 19567 16507
rect 19625 16473 19659 16507
rect 21833 16473 21867 16507
rect 28457 16473 28491 16507
rect 28549 16473 28583 16507
rect 29929 16473 29963 16507
rect 6377 16405 6411 16439
rect 9505 16405 9539 16439
rect 17693 16405 17727 16439
rect 24685 16405 24719 16439
rect 27353 16405 27387 16439
rect 3893 16201 3927 16235
rect 5181 16201 5215 16235
rect 25697 16201 25731 16235
rect 28181 16201 28215 16235
rect 8493 16133 8527 16167
rect 8585 16133 8619 16167
rect 9689 16133 9723 16167
rect 9781 16133 9815 16167
rect 12265 16133 12299 16167
rect 13461 16133 13495 16167
rect 14381 16133 14415 16167
rect 15669 16133 15703 16167
rect 18521 16133 18555 16167
rect 20085 16133 20119 16167
rect 21189 16133 21223 16167
rect 22845 16133 22879 16167
rect 1593 16065 1627 16099
rect 2513 16065 2547 16099
rect 4077 16065 4111 16099
rect 5089 16065 5123 16099
rect 5825 16065 5859 16099
rect 7113 16065 7147 16099
rect 7757 16065 7791 16099
rect 9137 16065 9171 16099
rect 14841 16065 14875 16099
rect 17049 16065 17083 16099
rect 17693 16065 17727 16099
rect 21097 16065 21131 16099
rect 22017 16065 22051 16099
rect 25237 16065 25271 16099
rect 27537 16065 27571 16099
rect 28825 16065 28859 16099
rect 30297 16065 30331 16099
rect 30941 16065 30975 16099
rect 38025 16065 38059 16099
rect 7849 15997 7883 16031
rect 10701 15997 10735 16031
rect 12173 15997 12207 16031
rect 12817 15997 12851 16031
rect 13369 15997 13403 16031
rect 15577 15997 15611 16031
rect 18429 15997 18463 16031
rect 18705 15997 18739 16031
rect 19993 15997 20027 16031
rect 22753 15997 22787 16031
rect 23121 15997 23155 16031
rect 25053 15997 25087 16031
rect 27721 15997 27755 16031
rect 29285 15997 29319 16031
rect 16129 15929 16163 15963
rect 20545 15929 20579 15963
rect 30113 15929 30147 15963
rect 1777 15861 1811 15895
rect 2329 15861 2363 15895
rect 5917 15861 5951 15895
rect 7205 15861 7239 15895
rect 14933 15861 14967 15895
rect 17141 15861 17175 15895
rect 17785 15861 17819 15895
rect 22109 15861 22143 15895
rect 28641 15861 28675 15895
rect 30757 15861 30791 15895
rect 38209 15861 38243 15895
rect 1777 15657 1811 15691
rect 27997 15657 28031 15691
rect 28549 15657 28583 15691
rect 6561 15521 6595 15555
rect 9229 15521 9263 15555
rect 9781 15521 9815 15555
rect 11897 15521 11931 15555
rect 12725 15521 12759 15555
rect 14565 15521 14599 15555
rect 15577 15521 15611 15555
rect 18153 15521 18187 15555
rect 20453 15521 20487 15555
rect 24593 15521 24627 15555
rect 25237 15521 25271 15555
rect 27537 15521 27571 15555
rect 1961 15453 1995 15487
rect 4537 15453 4571 15487
rect 5181 15453 5215 15487
rect 5825 15453 5859 15487
rect 6469 15453 6503 15487
rect 7297 15453 7331 15487
rect 7757 15453 7791 15487
rect 8401 15453 8435 15487
rect 17509 15453 17543 15487
rect 17693 15453 17727 15487
rect 18705 15453 18739 15487
rect 19717 15453 19751 15487
rect 21925 15453 21959 15487
rect 22569 15453 22603 15487
rect 23857 15453 23891 15487
rect 24777 15453 24811 15487
rect 26525 15453 26559 15487
rect 27353 15453 27387 15487
rect 28457 15453 28491 15487
rect 29929 15453 29963 15487
rect 7849 15385 7883 15419
rect 9321 15385 9355 15419
rect 10885 15385 10919 15419
rect 10977 15385 11011 15419
rect 12817 15385 12851 15419
rect 13737 15385 13771 15419
rect 14657 15385 14691 15419
rect 16129 15385 16163 15419
rect 16957 15385 16991 15419
rect 20545 15385 20579 15419
rect 21465 15385 21499 15419
rect 25697 15385 25731 15419
rect 38117 15385 38151 15419
rect 2421 15317 2455 15351
rect 4629 15317 4663 15351
rect 5273 15317 5307 15351
rect 5917 15317 5951 15351
rect 7113 15317 7147 15351
rect 8493 15317 8527 15351
rect 18797 15317 18831 15351
rect 19809 15317 19843 15351
rect 22017 15317 22051 15351
rect 22661 15317 22695 15351
rect 23949 15317 23983 15351
rect 26341 15317 26375 15351
rect 29745 15317 29779 15351
rect 38209 15317 38243 15351
rect 6929 15113 6963 15147
rect 26065 15113 26099 15147
rect 5273 15045 5307 15079
rect 8861 15045 8895 15079
rect 10609 15045 10643 15079
rect 12725 15045 12759 15079
rect 13369 15045 13403 15079
rect 13461 15045 13495 15079
rect 17601 15045 17635 15079
rect 19809 15045 19843 15079
rect 22201 15045 22235 15079
rect 24685 15045 24719 15079
rect 1777 14977 1811 15011
rect 2421 14977 2455 15011
rect 2605 14977 2639 15011
rect 3893 14977 3927 15011
rect 5181 14977 5215 15011
rect 5825 14977 5859 15011
rect 6653 14977 6687 15011
rect 8033 14977 8067 15011
rect 12173 14977 12207 15011
rect 14933 14977 14967 15011
rect 16129 14977 16163 15011
rect 18981 14977 19015 15011
rect 26249 14977 26283 15011
rect 27169 14977 27203 15011
rect 28641 14977 28675 15011
rect 29745 14977 29779 15011
rect 31217 14977 31251 15011
rect 33149 14977 33183 15011
rect 4537 14909 4571 14943
rect 8770 14909 8804 14943
rect 9137 14909 9171 14943
rect 10517 14909 10551 14943
rect 14381 14909 14415 14943
rect 15209 14909 15243 14943
rect 17509 14909 17543 14943
rect 18153 14909 18187 14943
rect 19717 14909 19751 14943
rect 20085 14909 20119 14943
rect 22109 14909 22143 14943
rect 23121 14909 23155 14943
rect 24593 14909 24627 14943
rect 24869 14909 24903 14943
rect 27353 14909 27387 14943
rect 28457 14909 28491 14943
rect 11069 14841 11103 14875
rect 1869 14773 1903 14807
rect 3065 14773 3099 14807
rect 3985 14773 4019 14807
rect 5917 14773 5951 14807
rect 8125 14773 8159 14807
rect 16221 14773 16255 14807
rect 19073 14773 19107 14807
rect 27813 14773 27847 14807
rect 28825 14773 28859 14807
rect 29561 14773 29595 14807
rect 31033 14773 31067 14807
rect 32965 14773 32999 14807
rect 1593 14569 1627 14603
rect 3065 14569 3099 14603
rect 6285 14569 6319 14603
rect 12817 14569 12851 14603
rect 20545 14569 20579 14603
rect 23213 14501 23247 14535
rect 28825 14501 28859 14535
rect 2697 14433 2731 14467
rect 7849 14433 7883 14467
rect 13553 14433 13587 14467
rect 16037 14433 16071 14467
rect 21465 14433 21499 14467
rect 22109 14433 22143 14467
rect 25697 14433 25731 14467
rect 1777 14365 1811 14399
rect 2513 14365 2547 14399
rect 3985 14365 4019 14399
rect 4905 14365 4939 14399
rect 5549 14365 5583 14399
rect 6193 14365 6227 14399
rect 6837 14365 6871 14399
rect 6929 14365 6963 14399
rect 9137 14365 9171 14399
rect 11069 14365 11103 14399
rect 13277 14365 13311 14399
rect 14289 14365 14323 14399
rect 15301 14365 15335 14399
rect 18061 14365 18095 14399
rect 18705 14365 18739 14399
rect 19809 14365 19843 14399
rect 20453 14365 20487 14399
rect 23765 14365 23799 14399
rect 24593 14365 24627 14399
rect 28733 14365 28767 14399
rect 29745 14365 29779 14399
rect 29837 14365 29871 14399
rect 35081 14365 35115 14399
rect 4997 14297 5031 14331
rect 7573 14297 7607 14331
rect 7665 14297 7699 14331
rect 9873 14297 9907 14331
rect 11345 14297 11379 14331
rect 14565 14297 14599 14331
rect 16129 14297 16163 14331
rect 17049 14297 17083 14331
rect 21557 14297 21591 14331
rect 22661 14297 22695 14331
rect 22753 14297 22787 14331
rect 25789 14297 25823 14331
rect 26709 14297 26743 14331
rect 27261 14297 27295 14331
rect 27353 14297 27387 14331
rect 28273 14297 28307 14331
rect 4077 14229 4111 14263
rect 5641 14229 5675 14263
rect 15393 14229 15427 14263
rect 18153 14229 18187 14263
rect 18797 14229 18831 14263
rect 19901 14229 19935 14263
rect 23857 14229 23891 14263
rect 24685 14229 24719 14263
rect 34897 14229 34931 14263
rect 2973 14025 3007 14059
rect 3709 14025 3743 14059
rect 6929 14025 6963 14059
rect 9229 14025 9263 14059
rect 18245 14025 18279 14059
rect 20545 14025 20579 14059
rect 21189 14025 21223 14059
rect 25697 14025 25731 14059
rect 26341 14025 26375 14059
rect 27813 14025 27847 14059
rect 4353 13957 4387 13991
rect 7757 13957 7791 13991
rect 11989 13957 12023 13991
rect 14933 13957 14967 13991
rect 22477 13957 22511 13991
rect 23397 13957 23431 13991
rect 24041 13957 24075 13991
rect 24961 13957 24995 13991
rect 1593 13889 1627 13923
rect 3157 13889 3191 13923
rect 3617 13889 3651 13923
rect 4261 13889 4295 13923
rect 4905 13889 4939 13923
rect 5825 13889 5859 13923
rect 6837 13889 6871 13923
rect 10241 13889 10275 13923
rect 11897 13889 11931 13923
rect 16865 13889 16899 13923
rect 18153 13889 18187 13923
rect 21097 13889 21131 13923
rect 25605 13889 25639 13923
rect 26249 13889 26283 13923
rect 27169 13889 27203 13923
rect 27261 13889 27295 13923
rect 28733 13889 28767 13923
rect 29837 13889 29871 13923
rect 31493 13889 31527 13923
rect 38025 13889 38059 13923
rect 4997 13821 5031 13855
rect 5917 13821 5951 13855
rect 7481 13821 7515 13855
rect 11069 13821 11103 13855
rect 12541 13821 12575 13855
rect 15669 13821 15703 13855
rect 17141 13821 17175 13855
rect 18797 13821 18831 13855
rect 19073 13821 19107 13855
rect 22385 13821 22419 13855
rect 23949 13821 23983 13855
rect 28917 13821 28951 13855
rect 1777 13685 1811 13719
rect 12798 13685 12832 13719
rect 14289 13685 14323 13719
rect 29101 13685 29135 13719
rect 31309 13685 31343 13719
rect 38209 13685 38243 13719
rect 18337 13481 18371 13515
rect 21833 13481 21867 13515
rect 27353 13481 27387 13515
rect 29745 13481 29779 13515
rect 8585 13413 8619 13447
rect 13645 13413 13679 13447
rect 6837 13345 6871 13379
rect 9137 13345 9171 13379
rect 10885 13345 10919 13379
rect 12173 13345 12207 13379
rect 14565 13345 14599 13379
rect 21189 13345 21223 13379
rect 23213 13345 23247 13379
rect 23489 13345 23523 13379
rect 24685 13345 24719 13379
rect 24961 13345 24995 13379
rect 26893 13345 26927 13379
rect 27905 13345 27939 13379
rect 28549 13345 28583 13379
rect 4721 13277 4755 13311
rect 5181 13277 5215 13311
rect 5825 13277 5859 13311
rect 5917 13277 5951 13311
rect 11897 13277 11931 13311
rect 14289 13277 14323 13311
rect 16589 13277 16623 13311
rect 19441 13277 19475 13311
rect 21741 13277 21775 13311
rect 22385 13277 22419 13311
rect 26709 13277 26743 13311
rect 27813 13277 27847 13311
rect 28733 13277 28767 13311
rect 29929 13277 29963 13311
rect 5273 13209 5307 13243
rect 7113 13209 7147 13243
rect 9413 13209 9447 13243
rect 16865 13209 16899 13243
rect 19717 13209 19751 13243
rect 23305 13209 23339 13243
rect 24777 13209 24811 13243
rect 4537 13141 4571 13175
rect 16037 13141 16071 13175
rect 22477 13141 22511 13175
rect 29193 13141 29227 13175
rect 30757 13141 30791 13175
rect 4077 12937 4111 12971
rect 5917 12937 5951 12971
rect 16221 12937 16255 12971
rect 22477 12937 22511 12971
rect 23121 12937 23155 12971
rect 26341 12937 26375 12971
rect 29193 12937 29227 12971
rect 17141 12869 17175 12903
rect 24317 12869 24351 12903
rect 1593 12801 1627 12835
rect 3985 12801 4019 12835
rect 5181 12801 5215 12835
rect 5825 12801 5859 12835
rect 7113 12801 7147 12835
rect 7757 12801 7791 12835
rect 10149 12801 10183 12835
rect 12081 12801 12115 12835
rect 14473 12801 14507 12835
rect 19441 12801 19475 12835
rect 22385 12801 22419 12835
rect 23029 12801 23063 12835
rect 25697 12801 25731 12835
rect 29101 12801 29135 12835
rect 30665 12801 30699 12835
rect 30849 12801 30883 12835
rect 38025 12801 38059 12835
rect 5273 12733 5307 12767
rect 8033 12733 8067 12767
rect 10333 12733 10367 12767
rect 12357 12733 12391 12767
rect 14749 12733 14783 12767
rect 16865 12733 16899 12767
rect 18613 12733 18647 12767
rect 19717 12733 19751 12767
rect 21465 12733 21499 12767
rect 24225 12733 24259 12767
rect 25881 12733 25915 12767
rect 27997 12733 28031 12767
rect 28181 12733 28215 12767
rect 24777 12665 24811 12699
rect 31033 12665 31067 12699
rect 1777 12597 1811 12631
rect 7205 12597 7239 12631
rect 9505 12597 9539 12631
rect 13829 12597 13863 12631
rect 28641 12597 28675 12631
rect 38209 12597 38243 12631
rect 9873 12393 9907 12427
rect 10682 12393 10716 12427
rect 13645 12393 13679 12427
rect 18521 12393 18555 12427
rect 26433 12393 26467 12427
rect 28457 12393 28491 12427
rect 24961 12325 24995 12359
rect 6745 12257 6779 12291
rect 7021 12257 7055 12291
rect 12449 12257 12483 12291
rect 14933 12257 14967 12291
rect 15945 12257 15979 12291
rect 17969 12257 18003 12291
rect 19993 12257 20027 12291
rect 20269 12257 20303 12291
rect 22017 12257 22051 12291
rect 22937 12257 22971 12291
rect 23489 12257 23523 12291
rect 9137 12189 9171 12223
rect 9781 12189 9815 12223
rect 10425 12189 10459 12223
rect 12909 12189 12943 12223
rect 13553 12189 13587 12223
rect 14759 12189 14793 12223
rect 18429 12189 18463 12223
rect 24593 12189 24627 12223
rect 24777 12189 24811 12223
rect 25697 12189 25731 12223
rect 26341 12189 26375 12223
rect 28365 12189 28399 12223
rect 30113 12189 30147 12223
rect 16221 12121 16255 12155
rect 23029 12121 23063 12155
rect 8493 12053 8527 12087
rect 9229 12053 9263 12087
rect 13001 12053 13035 12087
rect 25789 12053 25823 12087
rect 29929 12053 29963 12087
rect 18889 11849 18923 11883
rect 22385 11849 22419 11883
rect 24777 11849 24811 11883
rect 30481 11849 30515 11883
rect 32413 11849 32447 11883
rect 11989 11781 12023 11815
rect 14289 11781 14323 11815
rect 17417 11781 17451 11815
rect 23305 11781 23339 11815
rect 25513 11781 25547 11815
rect 27261 11781 27295 11815
rect 27353 11781 27387 11815
rect 29377 11781 29411 11815
rect 29469 11781 29503 11815
rect 7941 11713 7975 11747
rect 9965 11713 9999 11747
rect 10977 11713 11011 11747
rect 11713 11713 11747 11747
rect 17141 11713 17175 11747
rect 19441 11713 19475 11747
rect 22293 11713 22327 11747
rect 24685 11713 24719 11747
rect 30665 11713 30699 11747
rect 32321 11713 32355 11747
rect 8217 11645 8251 11679
rect 14013 11645 14047 11679
rect 19717 11645 19751 11679
rect 21465 11645 21499 11679
rect 23213 11645 23247 11679
rect 24225 11645 24259 11679
rect 25421 11645 25455 11679
rect 26341 11645 26375 11679
rect 27629 11645 27663 11679
rect 29653 11645 29687 11679
rect 11069 11509 11103 11543
rect 13461 11509 13495 11543
rect 15761 11509 15795 11543
rect 11976 11305 12010 11339
rect 23213 11305 23247 11339
rect 23857 11305 23891 11339
rect 27905 11305 27939 11339
rect 38209 11237 38243 11271
rect 6837 11169 6871 11203
rect 7113 11169 7147 11203
rect 8585 11169 8619 11203
rect 9781 11169 9815 11203
rect 11713 11169 11747 11203
rect 13737 11169 13771 11203
rect 14289 11169 14323 11203
rect 16773 11169 16807 11203
rect 17049 11169 17083 11203
rect 18521 11169 18555 11203
rect 20177 11169 20211 11203
rect 26249 11169 26283 11203
rect 28457 11169 28491 11203
rect 1777 11101 1811 11135
rect 2513 11101 2547 11135
rect 9505 11101 9539 11135
rect 23121 11101 23155 11135
rect 23765 11101 23799 11135
rect 27813 11101 27847 11135
rect 28641 11101 28675 11135
rect 29929 11101 29963 11135
rect 37381 11101 37415 11135
rect 38025 11101 38059 11135
rect 14565 11033 14599 11067
rect 16313 11033 16347 11067
rect 19441 11033 19475 11067
rect 25145 11033 25179 11067
rect 25237 11033 25271 11067
rect 25789 11033 25823 11067
rect 29101 11033 29135 11067
rect 1593 10965 1627 10999
rect 2329 10965 2363 10999
rect 11253 10965 11287 10999
rect 29745 10965 29779 10999
rect 37473 10965 37507 10999
rect 1593 10761 1627 10795
rect 3801 10761 3835 10795
rect 9045 10761 9079 10795
rect 12173 10761 12207 10795
rect 12817 10761 12851 10795
rect 15117 10761 15151 10795
rect 25605 10761 25639 10795
rect 29285 10761 29319 10795
rect 35173 10761 35207 10795
rect 23765 10693 23799 10727
rect 1777 10625 1811 10659
rect 2605 10625 2639 10659
rect 3709 10625 3743 10659
rect 10149 10625 10183 10659
rect 10793 10625 10827 10659
rect 10885 10625 10919 10659
rect 12081 10625 12115 10659
rect 12725 10625 12759 10659
rect 13369 10625 13403 10659
rect 19257 10625 19291 10659
rect 22569 10625 22603 10659
rect 25513 10625 25547 10659
rect 29469 10625 29503 10659
rect 34529 10625 34563 10659
rect 35357 10625 35391 10659
rect 38025 10625 38059 10659
rect 7297 10557 7331 10591
rect 7573 10557 7607 10591
rect 13645 10557 13679 10591
rect 16957 10557 16991 10591
rect 17233 10557 17267 10591
rect 18705 10557 18739 10591
rect 19533 10557 19567 10591
rect 23673 10557 23707 10591
rect 23949 10557 23983 10591
rect 10241 10489 10275 10523
rect 2697 10421 2731 10455
rect 21005 10421 21039 10455
rect 22661 10421 22695 10455
rect 34345 10421 34379 10455
rect 38209 10421 38243 10455
rect 3985 10217 4019 10251
rect 8585 10217 8619 10251
rect 11437 10217 11471 10251
rect 18613 10217 18647 10251
rect 23121 10217 23155 10251
rect 37841 10217 37875 10251
rect 2697 10149 2731 10183
rect 13645 10149 13679 10183
rect 3341 10081 3375 10115
rect 7113 10081 7147 10115
rect 18061 10081 18095 10115
rect 21557 10081 21591 10115
rect 24685 10081 24719 10115
rect 1961 10013 1995 10047
rect 2605 10013 2639 10047
rect 3249 10013 3283 10047
rect 4169 10013 4203 10047
rect 6837 10013 6871 10047
rect 9689 10013 9723 10047
rect 11897 10013 11931 10047
rect 14933 10013 14967 10047
rect 16037 10013 16071 10047
rect 18521 10013 18555 10047
rect 19809 10013 19843 10047
rect 23029 10013 23063 10047
rect 38025 10013 38059 10047
rect 2053 9945 2087 9979
rect 9965 9945 9999 9979
rect 12173 9945 12207 9979
rect 16313 9945 16347 9979
rect 20085 9945 20119 9979
rect 24777 9945 24811 9979
rect 25697 9945 25731 9979
rect 15025 9877 15059 9911
rect 4537 9673 4571 9707
rect 10977 9605 11011 9639
rect 15485 9605 15519 9639
rect 23765 9605 23799 9639
rect 30205 9605 30239 9639
rect 1685 9537 1719 9571
rect 2329 9537 2363 9571
rect 3249 9537 3283 9571
rect 3893 9537 3927 9571
rect 4713 9537 4747 9571
rect 5365 9537 5399 9571
rect 10241 9537 10275 9571
rect 11713 9537 11747 9571
rect 14657 9537 14691 9571
rect 16037 9537 16071 9571
rect 17233 9537 17267 9571
rect 30113 9537 30147 9571
rect 30941 9537 30975 9571
rect 31585 9537 31619 9571
rect 2421 9469 2455 9503
rect 5457 9469 5491 9503
rect 7757 9469 7791 9503
rect 8033 9469 8067 9503
rect 12357 9469 12391 9503
rect 12633 9469 12667 9503
rect 17509 9469 17543 9503
rect 18981 9469 19015 9503
rect 19441 9469 19475 9503
rect 19717 9469 19751 9503
rect 21189 9469 21223 9503
rect 23673 9469 23707 9503
rect 24041 9469 24075 9503
rect 29377 9469 29411 9503
rect 3341 9401 3375 9435
rect 3985 9401 4019 9435
rect 30757 9401 30791 9435
rect 1777 9333 1811 9367
rect 9505 9333 9539 9367
rect 11805 9333 11839 9367
rect 14105 9333 14139 9367
rect 16129 9333 16163 9367
rect 31401 9333 31435 9367
rect 7100 9129 7134 9163
rect 10885 9129 10919 9163
rect 23029 9129 23063 9163
rect 23673 9129 23707 9163
rect 4169 9061 4203 9095
rect 13093 9061 13127 9095
rect 9137 8993 9171 9027
rect 9413 8993 9447 9027
rect 11345 8993 11379 9027
rect 14381 8993 14415 9027
rect 18705 8993 18739 9027
rect 19625 8993 19659 9027
rect 29929 8993 29963 9027
rect 30941 8993 30975 9027
rect 1593 8925 1627 8959
rect 2329 8925 2363 8959
rect 3249 8925 3283 8959
rect 4353 8925 4387 8959
rect 4997 8925 5031 8959
rect 6837 8925 6871 8959
rect 16589 8925 16623 8959
rect 21649 8925 21683 8959
rect 22937 8925 22971 8959
rect 23581 8925 23615 8959
rect 28641 8925 28675 8959
rect 29745 8925 29779 8959
rect 30849 8925 30883 8959
rect 38301 8925 38335 8959
rect 2421 8857 2455 8891
rect 5457 8857 5491 8891
rect 6285 8857 6319 8891
rect 11621 8857 11655 8891
rect 14657 8857 14691 8891
rect 17969 8857 18003 8891
rect 19901 8857 19935 8891
rect 24961 8857 24995 8891
rect 25053 8857 25087 8891
rect 25973 8857 26007 8891
rect 1777 8789 1811 8823
rect 3065 8789 3099 8823
rect 4813 8789 4847 8823
rect 8585 8789 8619 8823
rect 16129 8789 16163 8823
rect 16681 8789 16715 8823
rect 28733 8789 28767 8823
rect 30389 8789 30423 8823
rect 38117 8789 38151 8823
rect 1593 8585 1627 8619
rect 2237 8585 2271 8619
rect 22937 8585 22971 8619
rect 23765 8585 23799 8619
rect 24409 8585 24443 8619
rect 25053 8585 25087 8619
rect 25973 8585 26007 8619
rect 29929 8585 29963 8619
rect 4537 8517 4571 8551
rect 6653 8517 6687 8551
rect 7941 8517 7975 8551
rect 12357 8517 12391 8551
rect 13185 8517 13219 8551
rect 14933 8517 14967 8551
rect 15393 8517 15427 8551
rect 17141 8517 17175 8551
rect 1777 8449 1811 8483
rect 2421 8449 2455 8483
rect 3065 8449 3099 8483
rect 3801 8449 3835 8483
rect 4261 8449 4295 8483
rect 6561 8449 6595 8483
rect 7205 8449 7239 8483
rect 10977 8449 11011 8483
rect 12265 8449 12299 8483
rect 12909 8449 12943 8483
rect 16865 8449 16899 8483
rect 19073 8449 19107 8483
rect 22845 8449 22879 8483
rect 23673 8449 23707 8483
rect 24317 8449 24351 8483
rect 24961 8449 24995 8483
rect 25881 8449 25915 8483
rect 27353 8449 27387 8483
rect 28457 8449 28491 8483
rect 29285 8449 29319 8483
rect 29469 8449 29503 8483
rect 30389 8449 30423 8483
rect 8585 8381 8619 8415
rect 8861 8381 8895 8415
rect 10333 8381 10367 8415
rect 11069 8381 11103 8415
rect 16129 8381 16163 8415
rect 19349 8381 19383 8415
rect 21097 8381 21131 8415
rect 2881 8313 2915 8347
rect 6009 8313 6043 8347
rect 18613 8313 18647 8347
rect 27169 8313 27203 8347
rect 28641 8313 28675 8347
rect 30481 8313 30515 8347
rect 3617 8245 3651 8279
rect 1961 8041 1995 8075
rect 5457 8041 5491 8075
rect 14920 8041 14954 8075
rect 18889 8041 18923 8075
rect 23305 8041 23339 8075
rect 24685 8041 24719 8075
rect 4077 7973 4111 8007
rect 8493 7973 8527 8007
rect 10885 7973 10919 8007
rect 16405 7973 16439 8007
rect 21741 7973 21775 8007
rect 25329 7973 25363 8007
rect 6745 7905 6779 7939
rect 9137 7905 9171 7939
rect 9413 7905 9447 7939
rect 14657 7905 14691 7939
rect 17141 7905 17175 7939
rect 17417 7905 17451 7939
rect 23949 7905 23983 7939
rect 27261 7905 27295 7939
rect 37749 7905 37783 7939
rect 2145 7837 2179 7871
rect 2605 7837 2639 7871
rect 3249 7837 3283 7871
rect 3985 7837 4019 7871
rect 4721 7837 4755 7871
rect 5365 7837 5399 7871
rect 6009 7837 6043 7871
rect 13553 7837 13587 7871
rect 19993 7837 20027 7871
rect 23213 7837 23247 7871
rect 23857 7837 23891 7871
rect 24593 7837 24627 7871
rect 25237 7837 25271 7871
rect 27721 7837 27755 7871
rect 37473 7837 37507 7871
rect 4813 7769 4847 7803
rect 7021 7769 7055 7803
rect 11989 7769 12023 7803
rect 20269 7769 20303 7803
rect 26249 7769 26283 7803
rect 26341 7769 26375 7803
rect 27813 7769 27847 7803
rect 2697 7701 2731 7735
rect 3341 7701 3375 7735
rect 6101 7701 6135 7735
rect 2605 7497 2639 7531
rect 13645 7497 13679 7531
rect 15945 7497 15979 7531
rect 25145 7497 25179 7531
rect 25789 7497 25823 7531
rect 27813 7497 27847 7531
rect 38117 7497 38151 7531
rect 17785 7429 17819 7463
rect 22753 7429 22787 7463
rect 23949 7429 23983 7463
rect 24041 7429 24075 7463
rect 26433 7429 26467 7463
rect 3249 7361 3283 7395
rect 3341 7361 3375 7395
rect 4077 7361 4111 7395
rect 4537 7361 4571 7395
rect 5181 7361 5215 7395
rect 5825 7361 5859 7395
rect 7113 7361 7147 7395
rect 14197 7361 14231 7395
rect 16865 7361 16899 7395
rect 17509 7361 17543 7395
rect 19717 7361 19751 7395
rect 22017 7361 22051 7395
rect 25053 7361 25087 7395
rect 25697 7361 25731 7395
rect 26341 7361 26375 7395
rect 27169 7361 27203 7395
rect 34253 7361 34287 7395
rect 38301 7361 38335 7395
rect 1961 7293 1995 7327
rect 2145 7293 2179 7327
rect 7389 7293 7423 7327
rect 8861 7293 8895 7327
rect 9321 7293 9355 7327
rect 9597 7293 9631 7327
rect 11897 7293 11931 7327
rect 12173 7293 12207 7327
rect 14473 7293 14507 7327
rect 19993 7293 20027 7327
rect 24225 7293 24259 7327
rect 4629 7225 4663 7259
rect 5273 7225 5307 7259
rect 5917 7225 5951 7259
rect 3893 7157 3927 7191
rect 11069 7157 11103 7191
rect 16957 7157 16991 7191
rect 19257 7157 19291 7191
rect 21465 7157 21499 7191
rect 27261 7157 27295 7191
rect 34345 7157 34379 7191
rect 2697 6953 2731 6987
rect 11976 6953 12010 6987
rect 17128 6953 17162 6987
rect 2421 6817 2455 6851
rect 4997 6817 5031 6851
rect 5641 6817 5675 6851
rect 6837 6817 6871 6851
rect 8585 6817 8619 6851
rect 14473 6817 14507 6851
rect 14749 6817 14783 6851
rect 16221 6817 16255 6851
rect 16865 6817 16899 6851
rect 18889 6817 18923 6851
rect 19717 6817 19751 6851
rect 22017 6817 22051 6851
rect 25237 6817 25271 6851
rect 26525 6817 26559 6851
rect 26801 6817 26835 6851
rect 1777 6749 1811 6783
rect 2237 6749 2271 6783
rect 4261 6749 4295 6783
rect 4353 6749 4387 6783
rect 4905 6749 4939 6783
rect 5549 6749 5583 6783
rect 6193 6749 6227 6783
rect 6285 6749 6319 6783
rect 9689 6749 9723 6783
rect 10333 6749 10367 6783
rect 11161 6749 11195 6783
rect 11713 6749 11747 6783
rect 21925 6749 21959 6783
rect 22569 6749 22603 6783
rect 23213 6749 23247 6783
rect 24041 6749 24075 6783
rect 27997 6749 28031 6783
rect 28641 6749 28675 6783
rect 7113 6681 7147 6715
rect 19993 6681 20027 6715
rect 24961 6681 24995 6715
rect 25053 6681 25087 6715
rect 26594 6681 26628 6715
rect 1593 6613 1627 6647
rect 9781 6613 9815 6647
rect 13461 6613 13495 6647
rect 21465 6613 21499 6647
rect 22661 6613 22695 6647
rect 23305 6613 23339 6647
rect 23857 6613 23891 6647
rect 28089 6613 28123 6647
rect 28733 6613 28767 6647
rect 5917 6409 5951 6443
rect 15761 6409 15795 6443
rect 27997 6409 28031 6443
rect 2973 6341 3007 6375
rect 3893 6341 3927 6375
rect 6561 6341 6595 6375
rect 8125 6341 8159 6375
rect 11989 6341 12023 6375
rect 14289 6341 14323 6375
rect 17509 6341 17543 6375
rect 23765 6341 23799 6375
rect 25329 6341 25363 6375
rect 25421 6341 25455 6375
rect 2145 6273 2179 6307
rect 4537 6273 4571 6307
rect 5181 6273 5215 6307
rect 5825 6273 5859 6307
rect 8033 6273 8067 6307
rect 8677 6273 8711 6307
rect 10977 6273 11011 6307
rect 14013 6273 14047 6307
rect 17233 6273 17267 6307
rect 19717 6273 19751 6307
rect 22385 6273 22419 6307
rect 27169 6273 27203 6307
rect 27445 6273 27479 6307
rect 27905 6273 27939 6307
rect 28549 6273 28583 6307
rect 30205 6273 30239 6307
rect 36829 6273 36863 6307
rect 2881 6205 2915 6239
rect 5273 6205 5307 6239
rect 7297 6205 7331 6239
rect 10425 6205 10459 6239
rect 11713 6205 11747 6239
rect 18981 6205 19015 6239
rect 19993 6205 20027 6239
rect 23673 6205 23707 6239
rect 23949 6205 23983 6239
rect 25605 6205 25639 6239
rect 4629 6137 4663 6171
rect 11069 6137 11103 6171
rect 13461 6137 13495 6171
rect 21465 6137 21499 6171
rect 28641 6137 28675 6171
rect 2237 6069 2271 6103
rect 8934 6069 8968 6103
rect 22569 6069 22603 6103
rect 30021 6069 30055 6103
rect 36645 6069 36679 6103
rect 2697 5865 2731 5899
rect 4800 5865 4834 5899
rect 6285 5865 6319 5899
rect 22385 5865 22419 5899
rect 26893 5865 26927 5899
rect 27537 5865 27571 5899
rect 1961 5797 1995 5831
rect 8493 5797 8527 5831
rect 11069 5797 11103 5831
rect 6745 5729 6779 5763
rect 9321 5729 9355 5763
rect 12265 5729 12299 5763
rect 13737 5729 13771 5763
rect 14381 5729 14415 5763
rect 16129 5729 16163 5763
rect 17141 5729 17175 5763
rect 18889 5729 18923 5763
rect 19809 5729 19843 5763
rect 23029 5729 23063 5763
rect 24685 5729 24719 5763
rect 2145 5661 2179 5695
rect 2605 5661 2639 5695
rect 3249 5661 3283 5695
rect 4537 5661 4571 5695
rect 11989 5661 12023 5695
rect 22293 5661 22327 5695
rect 26157 5661 26191 5695
rect 26249 5661 26283 5695
rect 26801 5661 26835 5695
rect 27445 5661 27479 5695
rect 28089 5661 28123 5695
rect 29745 5661 29779 5695
rect 38025 5661 38059 5695
rect 7021 5593 7055 5627
rect 9597 5593 9631 5627
rect 14657 5593 14691 5627
rect 17417 5593 17451 5627
rect 20085 5593 20119 5627
rect 23121 5593 23155 5627
rect 23673 5593 23707 5627
rect 24777 5593 24811 5627
rect 25697 5593 25731 5627
rect 3341 5525 3375 5559
rect 21557 5525 21591 5559
rect 28181 5525 28215 5559
rect 28733 5525 28767 5559
rect 29837 5525 29871 5559
rect 38209 5525 38243 5559
rect 1685 5321 1719 5355
rect 2421 5321 2455 5355
rect 3709 5321 3743 5355
rect 15945 5321 15979 5355
rect 28549 5321 28583 5355
rect 7481 5253 7515 5287
rect 9689 5253 9723 5287
rect 13737 5253 13771 5287
rect 17233 5253 17267 5287
rect 23305 5253 23339 5287
rect 25697 5253 25731 5287
rect 1593 5185 1627 5219
rect 2329 5185 2363 5219
rect 3157 5185 3191 5219
rect 3617 5185 3651 5219
rect 4261 5185 4295 5219
rect 6561 5185 6595 5219
rect 9413 5185 9447 5219
rect 19533 5185 19567 5219
rect 22477 5185 22511 5219
rect 24685 5185 24719 5219
rect 27169 5185 27203 5219
rect 27813 5185 27847 5219
rect 28457 5185 28491 5219
rect 29101 5185 29135 5219
rect 29745 5185 29779 5219
rect 30389 5185 30423 5219
rect 4537 5117 4571 5151
rect 7205 5117 7239 5151
rect 11161 5117 11195 5151
rect 11713 5117 11747 5151
rect 11989 5117 12023 5151
rect 14197 5117 14231 5151
rect 14473 5117 14507 5151
rect 16957 5117 16991 5151
rect 18705 5117 18739 5151
rect 19809 5117 19843 5151
rect 23213 5117 23247 5151
rect 24041 5117 24075 5151
rect 25605 5117 25639 5151
rect 25881 5117 25915 5151
rect 6009 5049 6043 5083
rect 27905 5049 27939 5083
rect 2973 4981 3007 5015
rect 6653 4981 6687 5015
rect 8953 4981 8987 5015
rect 21281 4981 21315 5015
rect 22569 4981 22603 5015
rect 24777 4981 24811 5015
rect 27261 4981 27295 5015
rect 29193 4981 29227 5015
rect 29837 4981 29871 5015
rect 30481 4981 30515 5015
rect 19796 4777 19830 4811
rect 30481 4777 30515 4811
rect 31769 4777 31803 4811
rect 38209 4777 38243 4811
rect 6285 4709 6319 4743
rect 11345 4709 11379 4743
rect 16313 4709 16347 4743
rect 21281 4709 21315 4743
rect 28825 4709 28859 4743
rect 2697 4641 2731 4675
rect 4813 4641 4847 4675
rect 6745 4641 6779 4675
rect 7021 4641 7055 4675
rect 9597 4641 9631 4675
rect 9873 4641 9907 4675
rect 11805 4641 11839 4675
rect 18797 4641 18831 4675
rect 19533 4641 19567 4675
rect 24961 4641 24995 4675
rect 25789 4641 25823 4675
rect 26985 4641 27019 4675
rect 1593 4573 1627 4607
rect 2605 4573 2639 4607
rect 3249 4573 3283 4607
rect 4537 4573 4571 4607
rect 14565 4573 14599 4607
rect 17049 4573 17083 4607
rect 21741 4573 21775 4607
rect 28089 4573 28123 4607
rect 28733 4573 28767 4607
rect 29745 4573 29779 4607
rect 30389 4573 30423 4607
rect 31217 4573 31251 4607
rect 31677 4573 31711 4607
rect 32321 4573 32355 4607
rect 33517 4573 33551 4607
rect 12081 4505 12115 4539
rect 14841 4505 14875 4539
rect 17325 4505 17359 4539
rect 22017 4505 22051 4539
rect 25046 4505 25080 4539
rect 26617 4505 26651 4539
rect 26709 4505 26743 4539
rect 38117 4505 38151 4539
rect 1777 4437 1811 4471
rect 3341 4437 3375 4471
rect 8493 4437 8527 4471
rect 13553 4437 13587 4471
rect 23489 4437 23523 4471
rect 28181 4437 28215 4471
rect 29837 4437 29871 4471
rect 31033 4437 31067 4471
rect 32413 4437 32447 4471
rect 33609 4437 33643 4471
rect 9873 4165 9907 4199
rect 16957 4165 16991 4199
rect 23305 4165 23339 4199
rect 24869 4165 24903 4199
rect 26074 4165 26108 4199
rect 28549 4165 28583 4199
rect 2053 4097 2087 4131
rect 2697 4097 2731 4131
rect 3341 4097 3375 4131
rect 4169 4097 4203 4131
rect 4629 4097 4663 4131
rect 5273 4097 5307 4131
rect 7113 4097 7147 4131
rect 9137 4097 9171 4131
rect 11989 4097 12023 4131
rect 20637 4097 20671 4131
rect 20729 4097 20763 4131
rect 21281 4097 21315 4131
rect 21373 4097 21407 4131
rect 22477 4097 22511 4131
rect 22569 4097 22603 4131
rect 27169 4097 27203 4131
rect 27813 4097 27847 4131
rect 28457 4097 28491 4131
rect 29101 4097 29135 4131
rect 29745 4097 29779 4131
rect 30389 4097 30423 4131
rect 30481 4097 30515 4131
rect 31033 4097 31067 4131
rect 32505 4097 32539 4131
rect 33885 4097 33919 4131
rect 2145 4029 2179 4063
rect 7389 4029 7423 4063
rect 10609 4029 10643 4063
rect 12265 4029 12299 4063
rect 14565 4029 14599 4063
rect 14841 4029 14875 4063
rect 16313 4029 16347 4063
rect 17693 4029 17727 4063
rect 18337 4029 18371 4063
rect 18613 4029 18647 4063
rect 23213 4029 23247 4063
rect 24133 4029 24167 4063
rect 24777 4029 24811 4063
rect 25053 4029 25087 4063
rect 25973 4029 26007 4063
rect 27261 4029 27295 4063
rect 29193 4029 29227 4063
rect 4721 3961 4755 3995
rect 26525 3961 26559 3995
rect 29837 3961 29871 3995
rect 2789 3893 2823 3927
rect 3433 3893 3467 3927
rect 3985 3893 4019 3927
rect 5457 3893 5491 3927
rect 13737 3893 13771 3927
rect 20085 3893 20119 3927
rect 27905 3893 27939 3927
rect 31125 3893 31159 3927
rect 32321 3893 32355 3927
rect 33701 3893 33735 3927
rect 38301 3893 38335 3927
rect 4077 3689 4111 3723
rect 7100 3689 7134 3723
rect 8585 3689 8619 3723
rect 10314 3689 10348 3723
rect 11805 3689 11839 3723
rect 16037 3689 16071 3723
rect 16497 3689 16531 3723
rect 23857 3689 23891 3723
rect 32965 3689 32999 3723
rect 6377 3621 6411 3655
rect 33609 3621 33643 3655
rect 2237 3553 2271 3587
rect 2697 3553 2731 3587
rect 4629 3553 4663 3587
rect 6837 3553 6871 3587
rect 17141 3553 17175 3587
rect 19441 3553 19475 3587
rect 19717 3553 19751 3587
rect 22661 3553 22695 3587
rect 27077 3553 27111 3587
rect 1593 3485 1627 3519
rect 2605 3485 2639 3519
rect 3249 3485 3283 3519
rect 3985 3485 4019 3519
rect 10057 3485 10091 3519
rect 12819 3485 12853 3519
rect 14289 3485 14323 3519
rect 16681 3485 16715 3519
rect 21925 3485 21959 3519
rect 23305 3485 23339 3519
rect 23765 3485 23799 3519
rect 25329 3485 25363 3519
rect 28549 3485 28583 3519
rect 29745 3485 29779 3519
rect 30389 3485 30423 3519
rect 31033 3485 31067 3519
rect 31861 3485 31895 3519
rect 33149 3485 33183 3519
rect 33793 3485 33827 3519
rect 38025 3485 38059 3519
rect 3341 3417 3375 3451
rect 4905 3417 4939 3451
rect 9229 3417 9263 3451
rect 9413 3417 9447 3451
rect 13645 3417 13679 3451
rect 14565 3417 14599 3451
rect 17417 3417 17451 3451
rect 21465 3417 21499 3451
rect 22753 3417 22787 3451
rect 24685 3417 24719 3451
rect 24777 3417 24811 3451
rect 25881 3417 25915 3451
rect 25973 3417 26007 3451
rect 26525 3417 26559 3451
rect 27169 3417 27203 3451
rect 28089 3417 28123 3451
rect 1777 3349 1811 3383
rect 18889 3349 18923 3383
rect 22017 3349 22051 3383
rect 28641 3349 28675 3383
rect 29837 3349 29871 3383
rect 30481 3349 30515 3383
rect 31125 3349 31159 3383
rect 31677 3349 31711 3383
rect 32321 3349 32355 3383
rect 38209 3349 38243 3383
rect 3065 3145 3099 3179
rect 6009 3145 6043 3179
rect 23765 3145 23799 3179
rect 32413 3145 32447 3179
rect 33057 3145 33091 3179
rect 36737 3145 36771 3179
rect 2421 3077 2455 3111
rect 8125 3077 8159 3111
rect 13645 3077 13679 3111
rect 16313 3077 16347 3111
rect 24317 3077 24351 3111
rect 24409 3077 24443 3111
rect 25973 3077 26007 3111
rect 27346 3077 27380 3111
rect 33701 3077 33735 3111
rect 1593 3009 1627 3043
rect 2329 3009 2363 3043
rect 2973 3009 3007 3043
rect 3801 3009 3835 3043
rect 4261 3009 4295 3043
rect 6561 3009 6595 3043
rect 7849 3009 7883 3043
rect 10333 3009 10367 3043
rect 10977 3009 11011 3043
rect 12173 3009 12207 3043
rect 12725 3009 12759 3043
rect 12909 3009 12943 3043
rect 13369 3009 13403 3043
rect 16129 3009 16163 3043
rect 17049 3009 17083 3043
rect 19257 3009 19291 3043
rect 22017 3009 22051 3043
rect 28365 3009 28399 3043
rect 29009 3009 29043 3043
rect 29653 3009 29687 3043
rect 30297 3009 30331 3043
rect 30941 3009 30975 3043
rect 31585 3009 31619 3043
rect 32321 3009 32355 3043
rect 32965 3009 32999 3043
rect 33609 3009 33643 3043
rect 35725 3009 35759 3043
rect 36921 3009 36955 3043
rect 38025 3009 38059 3043
rect 4537 2941 4571 2975
rect 9873 2941 9907 2975
rect 10425 2941 10459 2975
rect 11069 2941 11103 2975
rect 15117 2941 15151 2975
rect 17325 2941 17359 2975
rect 19533 2941 19567 2975
rect 22293 2941 22327 2975
rect 25145 2941 25179 2975
rect 25881 2941 25915 2975
rect 27261 2941 27295 2975
rect 27537 2941 27571 2975
rect 11989 2873 12023 2907
rect 26433 2873 26467 2907
rect 29101 2873 29135 2907
rect 35541 2873 35575 2907
rect 1777 2805 1811 2839
rect 3617 2805 3651 2839
rect 6745 2805 6779 2839
rect 18797 2805 18831 2839
rect 21005 2805 21039 2839
rect 28457 2805 28491 2839
rect 29745 2805 29779 2839
rect 30389 2805 30423 2839
rect 31033 2805 31067 2839
rect 31677 2805 31711 2839
rect 38209 2805 38243 2839
rect 6009 2601 6043 2635
rect 13737 2601 13771 2635
rect 18889 2601 18923 2635
rect 27261 2601 27295 2635
rect 28549 2601 28583 2635
rect 2605 2533 2639 2567
rect 16313 2533 16347 2567
rect 22017 2533 22051 2567
rect 36093 2533 36127 2567
rect 4261 2465 4295 2499
rect 6745 2465 6779 2499
rect 9413 2465 9447 2499
rect 9689 2465 9723 2499
rect 11989 2465 12023 2499
rect 14565 2465 14599 2499
rect 14841 2465 14875 2499
rect 17141 2465 17175 2499
rect 17417 2465 17451 2499
rect 19441 2465 19475 2499
rect 23029 2465 23063 2499
rect 24041 2465 24075 2499
rect 25973 2465 26007 2499
rect 26433 2465 26467 2499
rect 32597 2465 32631 2499
rect 37749 2465 37783 2499
rect 1685 2397 1719 2431
rect 2421 2397 2455 2431
rect 3157 2397 3191 2431
rect 22201 2397 22235 2431
rect 24593 2397 24627 2431
rect 24869 2397 24903 2431
rect 27169 2397 27203 2431
rect 27813 2397 27847 2431
rect 28733 2397 28767 2431
rect 29745 2397 29779 2431
rect 30481 2397 30515 2431
rect 31217 2397 31251 2431
rect 32321 2397 32355 2431
rect 33609 2397 33643 2431
rect 34897 2397 34931 2431
rect 35909 2397 35943 2431
rect 36645 2397 36679 2431
rect 37473 2397 37507 2431
rect 4537 2329 4571 2363
rect 7021 2329 7055 2363
rect 12265 2329 12299 2363
rect 19717 2329 19751 2363
rect 23121 2329 23155 2363
rect 26065 2329 26099 2363
rect 1869 2261 1903 2295
rect 3341 2261 3375 2295
rect 8493 2261 8527 2295
rect 11161 2261 11195 2295
rect 21189 2261 21223 2295
rect 27997 2261 28031 2295
rect 29929 2261 29963 2295
rect 30665 2261 30699 2295
rect 31309 2261 31343 2295
rect 33793 2261 33827 2295
rect 35081 2261 35115 2295
rect 36829 2261 36863 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 14553 37383 14611 37389
rect 14553 37349 14565 37383
rect 14599 37380 14611 37383
rect 20162 37380 20168 37392
rect 14599 37352 20168 37380
rect 14599 37349 14611 37352
rect 14553 37343 14611 37349
rect 20162 37340 20168 37352
rect 20220 37340 20226 37392
rect 36814 37340 36820 37392
rect 36872 37380 36878 37392
rect 39298 37380 39304 37392
rect 36872 37352 39304 37380
rect 36872 37340 36878 37352
rect 39298 37340 39304 37352
rect 39356 37340 39362 37392
rect 1946 37272 1952 37324
rect 2004 37312 2010 37324
rect 2041 37315 2099 37321
rect 2041 37312 2053 37315
rect 2004 37284 2053 37312
rect 2004 37272 2010 37284
rect 2041 37281 2053 37284
rect 2087 37281 2099 37315
rect 2041 37275 2099 37281
rect 3878 37272 3884 37324
rect 3936 37312 3942 37324
rect 3973 37315 4031 37321
rect 3973 37312 3985 37315
rect 3936 37284 3985 37312
rect 3936 37272 3942 37284
rect 3973 37281 3985 37284
rect 4019 37281 4031 37315
rect 3973 37275 4031 37281
rect 8386 37272 8392 37324
rect 8444 37312 8450 37324
rect 9125 37315 9183 37321
rect 9125 37312 9137 37315
rect 8444 37284 9137 37312
rect 8444 37272 8450 37284
rect 9125 37281 9137 37284
rect 9171 37281 9183 37315
rect 9125 37275 9183 37281
rect 12621 37315 12679 37321
rect 12621 37281 12633 37315
rect 12667 37312 12679 37315
rect 22462 37312 22468 37324
rect 12667 37284 22468 37312
rect 12667 37281 12679 37284
rect 12621 37275 12679 37281
rect 22462 37272 22468 37284
rect 22520 37272 22526 37324
rect 22554 37272 22560 37324
rect 22612 37312 22618 37324
rect 22649 37315 22707 37321
rect 22649 37312 22661 37315
rect 22612 37284 22661 37312
rect 22612 37272 22618 37284
rect 22649 37281 22661 37284
rect 22695 37281 22707 37315
rect 22649 37275 22707 37281
rect 29638 37272 29644 37324
rect 29696 37312 29702 37324
rect 37461 37315 37519 37321
rect 29696 37284 30236 37312
rect 29696 37272 29702 37284
rect 2317 37247 2375 37253
rect 2317 37213 2329 37247
rect 2363 37244 2375 37247
rect 2498 37244 2504 37256
rect 2363 37216 2504 37244
rect 2363 37213 2375 37216
rect 2317 37207 2375 37213
rect 2498 37204 2504 37216
rect 2556 37204 2562 37256
rect 4249 37247 4307 37253
rect 4249 37213 4261 37247
rect 4295 37213 4307 37247
rect 4249 37207 4307 37213
rect 4264 37176 4292 37207
rect 5166 37204 5172 37256
rect 5224 37244 5230 37256
rect 5445 37247 5503 37253
rect 5445 37244 5457 37247
rect 5224 37216 5457 37244
rect 5224 37204 5230 37216
rect 5445 37213 5457 37216
rect 5491 37213 5503 37247
rect 5445 37207 5503 37213
rect 5810 37204 5816 37256
rect 5868 37244 5874 37256
rect 6733 37247 6791 37253
rect 6733 37244 6745 37247
rect 5868 37216 6745 37244
rect 5868 37204 5874 37216
rect 6733 37213 6745 37216
rect 6779 37213 6791 37247
rect 6733 37207 6791 37213
rect 7098 37204 7104 37256
rect 7156 37244 7162 37256
rect 7377 37247 7435 37253
rect 7377 37244 7389 37247
rect 7156 37216 7389 37244
rect 7156 37204 7162 37216
rect 7377 37213 7389 37216
rect 7423 37213 7435 37247
rect 7377 37207 7435 37213
rect 8294 37204 8300 37256
rect 8352 37244 8358 37256
rect 9401 37247 9459 37253
rect 9401 37244 9413 37247
rect 8352 37216 9413 37244
rect 8352 37204 8358 37216
rect 9401 37213 9413 37216
rect 9447 37213 9459 37247
rect 10410 37244 10416 37256
rect 10371 37216 10416 37244
rect 9401 37207 9459 37213
rect 10410 37204 10416 37216
rect 10468 37204 10474 37256
rect 11606 37204 11612 37256
rect 11664 37244 11670 37256
rect 11885 37247 11943 37253
rect 11885 37244 11897 37247
rect 11664 37216 11897 37244
rect 11664 37204 11670 37216
rect 11885 37213 11897 37216
rect 11931 37213 11943 37247
rect 12434 37244 12440 37256
rect 12395 37216 12440 37244
rect 11885 37207 11943 37213
rect 12434 37204 12440 37216
rect 12492 37204 12498 37256
rect 13538 37204 13544 37256
rect 13596 37244 13602 37256
rect 14369 37247 14427 37253
rect 14369 37244 14381 37247
rect 13596 37216 14381 37244
rect 13596 37204 13602 37216
rect 14369 37213 14381 37216
rect 14415 37213 14427 37247
rect 15194 37244 15200 37256
rect 15155 37216 15200 37244
rect 14369 37207 14427 37213
rect 15194 37204 15200 37216
rect 15252 37204 15258 37256
rect 16022 37244 16028 37256
rect 15983 37216 16028 37244
rect 16022 37204 16028 37216
rect 16080 37204 16086 37256
rect 16853 37247 16911 37253
rect 16853 37213 16865 37247
rect 16899 37244 16911 37247
rect 16942 37244 16948 37256
rect 16899 37216 16948 37244
rect 16899 37213 16911 37216
rect 16853 37207 16911 37213
rect 16942 37204 16948 37216
rect 17000 37204 17006 37256
rect 18046 37204 18052 37256
rect 18104 37244 18110 37256
rect 18325 37247 18383 37253
rect 18325 37244 18337 37247
rect 18104 37216 18337 37244
rect 18104 37204 18110 37216
rect 18325 37213 18337 37216
rect 18371 37213 18383 37247
rect 20070 37244 20076 37256
rect 20031 37216 20076 37244
rect 18325 37207 18383 37213
rect 20070 37204 20076 37216
rect 20128 37204 20134 37256
rect 21174 37244 21180 37256
rect 21135 37216 21180 37244
rect 21174 37204 21180 37216
rect 21232 37204 21238 37256
rect 22922 37244 22928 37256
rect 22883 37216 22928 37244
rect 22922 37204 22928 37216
rect 22980 37204 22986 37256
rect 24486 37204 24492 37256
rect 24544 37244 24550 37256
rect 24765 37247 24823 37253
rect 24765 37244 24777 37247
rect 24544 37216 24777 37244
rect 24544 37204 24550 37216
rect 24765 37213 24777 37216
rect 24811 37213 24823 37247
rect 24765 37207 24823 37213
rect 25774 37204 25780 37256
rect 25832 37244 25838 37256
rect 26053 37247 26111 37253
rect 26053 37244 26065 37247
rect 25832 37216 26065 37244
rect 25832 37204 25838 37216
rect 26053 37213 26065 37216
rect 26099 37213 26111 37247
rect 27154 37244 27160 37256
rect 27115 37216 27160 37244
rect 26053 37207 26111 37213
rect 27154 37204 27160 37216
rect 27212 37204 27218 37256
rect 27706 37204 27712 37256
rect 27764 37244 27770 37256
rect 28077 37247 28135 37253
rect 28077 37244 28089 37247
rect 27764 37216 28089 37244
rect 27764 37204 27770 37216
rect 28077 37213 28089 37216
rect 28123 37213 28135 37247
rect 28077 37207 28135 37213
rect 28994 37204 29000 37256
rect 29052 37244 29058 37256
rect 29917 37247 29975 37253
rect 29917 37244 29929 37247
rect 29052 37216 29929 37244
rect 29052 37204 29058 37216
rect 29917 37213 29929 37216
rect 29963 37213 29975 37247
rect 30208 37244 30236 37284
rect 37461 37281 37473 37315
rect 37507 37312 37519 37315
rect 38654 37312 38660 37324
rect 37507 37284 38660 37312
rect 37507 37281 37519 37284
rect 37461 37275 37519 37281
rect 38654 37272 38660 37284
rect 38712 37272 38718 37324
rect 30561 37247 30619 37253
rect 30561 37244 30573 37247
rect 30208 37216 30573 37244
rect 29917 37207 29975 37213
rect 30561 37213 30573 37216
rect 30607 37213 30619 37247
rect 31018 37244 31024 37256
rect 30979 37216 31024 37244
rect 30561 37207 30619 37213
rect 31018 37204 31024 37216
rect 31076 37204 31082 37256
rect 32214 37204 32220 37256
rect 32272 37244 32278 37256
rect 32493 37247 32551 37253
rect 32493 37244 32505 37247
rect 32272 37216 32505 37244
rect 32272 37204 32278 37216
rect 32493 37213 32505 37216
rect 32539 37213 32551 37247
rect 32493 37207 32551 37213
rect 32953 37247 33011 37253
rect 32953 37213 32965 37247
rect 32999 37213 33011 37247
rect 32953 37207 33011 37213
rect 10502 37176 10508 37188
rect 4264 37148 10508 37176
rect 10502 37136 10508 37148
rect 10560 37136 10566 37188
rect 25498 37136 25504 37188
rect 25556 37176 25562 37188
rect 32968 37176 32996 37207
rect 33226 37204 33232 37256
rect 33284 37244 33290 37256
rect 34885 37247 34943 37253
rect 34885 37244 34897 37247
rect 33284 37216 34897 37244
rect 33284 37204 33290 37216
rect 34885 37213 34897 37216
rect 34931 37213 34943 37247
rect 34885 37207 34943 37213
rect 35986 37204 35992 37256
rect 36044 37244 36050 37256
rect 36173 37247 36231 37253
rect 36173 37244 36185 37247
rect 36044 37216 36185 37244
rect 36044 37204 36050 37216
rect 36173 37213 36185 37216
rect 36219 37213 36231 37247
rect 37734 37244 37740 37256
rect 37695 37216 37740 37244
rect 36173 37207 36231 37213
rect 37734 37204 37740 37216
rect 37792 37204 37798 37256
rect 25556 37148 32996 37176
rect 25556 37136 25562 37148
rect 5261 37111 5319 37117
rect 5261 37077 5273 37111
rect 5307 37108 5319 37111
rect 6178 37108 6184 37120
rect 5307 37080 6184 37108
rect 5307 37077 5319 37080
rect 5261 37071 5319 37077
rect 6178 37068 6184 37080
rect 6236 37068 6242 37120
rect 6546 37108 6552 37120
rect 6507 37080 6552 37108
rect 6546 37068 6552 37080
rect 6604 37068 6610 37120
rect 7193 37111 7251 37117
rect 7193 37077 7205 37111
rect 7239 37108 7251 37111
rect 7926 37108 7932 37120
rect 7239 37080 7932 37108
rect 7239 37077 7251 37080
rect 7193 37071 7251 37077
rect 7926 37068 7932 37080
rect 7984 37068 7990 37120
rect 10318 37068 10324 37120
rect 10376 37108 10382 37120
rect 10597 37111 10655 37117
rect 10597 37108 10609 37111
rect 10376 37080 10609 37108
rect 10376 37068 10382 37080
rect 10597 37077 10609 37080
rect 10643 37077 10655 37111
rect 11698 37108 11704 37120
rect 11659 37080 11704 37108
rect 10597 37071 10655 37077
rect 11698 37068 11704 37080
rect 11756 37068 11762 37120
rect 15010 37108 15016 37120
rect 14971 37080 15016 37108
rect 15010 37068 15016 37080
rect 15068 37068 15074 37120
rect 16114 37068 16120 37120
rect 16172 37108 16178 37120
rect 16209 37111 16267 37117
rect 16209 37108 16221 37111
rect 16172 37080 16221 37108
rect 16172 37068 16178 37080
rect 16209 37077 16221 37080
rect 16255 37077 16267 37111
rect 16209 37071 16267 37077
rect 16758 37068 16764 37120
rect 16816 37108 16822 37120
rect 17037 37111 17095 37117
rect 17037 37108 17049 37111
rect 16816 37080 17049 37108
rect 16816 37068 16822 37080
rect 17037 37077 17049 37080
rect 17083 37077 17095 37111
rect 17037 37071 17095 37077
rect 17126 37068 17132 37120
rect 17184 37108 17190 37120
rect 18141 37111 18199 37117
rect 18141 37108 18153 37111
rect 17184 37080 18153 37108
rect 17184 37068 17190 37080
rect 18141 37077 18153 37080
rect 18187 37077 18199 37111
rect 18141 37071 18199 37077
rect 19978 37068 19984 37120
rect 20036 37108 20042 37120
rect 20257 37111 20315 37117
rect 20257 37108 20269 37111
rect 20036 37080 20269 37108
rect 20036 37068 20042 37080
rect 20257 37077 20269 37080
rect 20303 37077 20315 37111
rect 20257 37071 20315 37077
rect 21266 37068 21272 37120
rect 21324 37108 21330 37120
rect 21361 37111 21419 37117
rect 21361 37108 21373 37111
rect 21324 37080 21373 37108
rect 21324 37068 21330 37080
rect 21361 37077 21373 37080
rect 21407 37077 21419 37111
rect 24578 37108 24584 37120
rect 24539 37080 24584 37108
rect 21361 37071 21419 37077
rect 24578 37068 24584 37080
rect 24636 37068 24642 37120
rect 25866 37108 25872 37120
rect 25827 37080 25872 37108
rect 25866 37068 25872 37080
rect 25924 37068 25930 37120
rect 26418 37068 26424 37120
rect 26476 37108 26482 37120
rect 27341 37111 27399 37117
rect 27341 37108 27353 37111
rect 26476 37080 27353 37108
rect 26476 37068 26482 37080
rect 27341 37077 27353 37080
rect 27387 37077 27399 37111
rect 27341 37071 27399 37077
rect 27430 37068 27436 37120
rect 27488 37108 27494 37120
rect 27893 37111 27951 37117
rect 27893 37108 27905 37111
rect 27488 37080 27905 37108
rect 27488 37068 27494 37080
rect 27893 37077 27905 37080
rect 27939 37077 27951 37111
rect 29730 37108 29736 37120
rect 29691 37080 29736 37108
rect 27893 37071 27951 37077
rect 29730 37068 29736 37080
rect 29788 37068 29794 37120
rect 30374 37108 30380 37120
rect 30335 37080 30380 37108
rect 30374 37068 30380 37080
rect 30432 37068 30438 37120
rect 30926 37068 30932 37120
rect 30984 37108 30990 37120
rect 31205 37111 31263 37117
rect 31205 37108 31217 37111
rect 30984 37080 31217 37108
rect 30984 37068 30990 37080
rect 31205 37077 31217 37080
rect 31251 37077 31263 37111
rect 31205 37071 31263 37077
rect 31294 37068 31300 37120
rect 31352 37108 31358 37120
rect 32309 37111 32367 37117
rect 32309 37108 32321 37111
rect 31352 37080 32321 37108
rect 31352 37068 31358 37080
rect 32309 37077 32321 37080
rect 32355 37077 32367 37111
rect 33134 37108 33140 37120
rect 33095 37080 33140 37108
rect 32309 37071 32367 37077
rect 33134 37068 33140 37080
rect 33192 37068 33198 37120
rect 34514 37068 34520 37120
rect 34572 37108 34578 37120
rect 35069 37111 35127 37117
rect 35069 37108 35081 37111
rect 34572 37080 35081 37108
rect 34572 37068 34578 37080
rect 35069 37077 35081 37080
rect 35115 37077 35127 37111
rect 35069 37071 35127 37077
rect 36078 37068 36084 37120
rect 36136 37108 36142 37120
rect 36357 37111 36415 37117
rect 36357 37108 36369 37111
rect 36136 37080 36369 37108
rect 36136 37068 36142 37080
rect 36357 37077 36369 37080
rect 36403 37077 36415 37111
rect 36357 37071 36415 37077
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 658 36864 664 36916
rect 716 36904 722 36916
rect 716 36876 3096 36904
rect 716 36864 722 36876
rect 1673 36839 1731 36845
rect 1673 36805 1685 36839
rect 1719 36836 1731 36839
rect 2958 36836 2964 36848
rect 1719 36808 2964 36836
rect 1719 36805 1731 36808
rect 1673 36799 1731 36805
rect 2958 36796 2964 36808
rect 3016 36796 3022 36848
rect 2774 36728 2780 36780
rect 2832 36768 2838 36780
rect 2869 36771 2927 36777
rect 2869 36768 2881 36771
rect 2832 36740 2881 36768
rect 2832 36728 2838 36740
rect 2869 36737 2881 36740
rect 2915 36737 2927 36771
rect 3068 36768 3096 36876
rect 6546 36864 6552 36916
rect 6604 36904 6610 36916
rect 9950 36904 9956 36916
rect 6604 36876 9956 36904
rect 6604 36864 6610 36876
rect 9950 36864 9956 36876
rect 10008 36864 10014 36916
rect 10410 36904 10416 36916
rect 10371 36876 10416 36904
rect 10410 36864 10416 36876
rect 10468 36864 10474 36916
rect 19334 36864 19340 36916
rect 19392 36904 19398 36916
rect 19613 36907 19671 36913
rect 19613 36904 19625 36907
rect 19392 36876 19625 36904
rect 19392 36864 19398 36876
rect 19613 36873 19625 36876
rect 19659 36873 19671 36907
rect 19613 36867 19671 36873
rect 23198 36864 23204 36916
rect 23256 36904 23262 36916
rect 23477 36907 23535 36913
rect 23477 36904 23489 36907
rect 23256 36876 23489 36904
rect 23256 36864 23262 36876
rect 23477 36873 23489 36876
rect 23523 36873 23535 36907
rect 27154 36904 27160 36916
rect 27115 36876 27160 36904
rect 23477 36867 23535 36873
rect 27154 36864 27160 36876
rect 27212 36864 27218 36916
rect 27982 36864 27988 36916
rect 28040 36904 28046 36916
rect 31018 36904 31024 36916
rect 28040 36876 31024 36904
rect 28040 36864 28046 36876
rect 31018 36864 31024 36876
rect 31076 36864 31082 36916
rect 36081 36907 36139 36913
rect 36081 36873 36093 36907
rect 36127 36904 36139 36907
rect 36170 36904 36176 36916
rect 36127 36876 36176 36904
rect 36127 36873 36139 36876
rect 36081 36867 36139 36873
rect 36170 36864 36176 36876
rect 36228 36864 36234 36916
rect 36814 36904 36820 36916
rect 36775 36876 36820 36904
rect 36814 36864 36820 36876
rect 36872 36864 36878 36916
rect 37366 36864 37372 36916
rect 37424 36904 37430 36916
rect 37645 36907 37703 36913
rect 37645 36904 37657 36907
rect 37424 36876 37657 36904
rect 37424 36864 37430 36876
rect 37645 36873 37657 36876
rect 37691 36873 37703 36907
rect 37645 36867 37703 36873
rect 3513 36771 3571 36777
rect 3513 36768 3525 36771
rect 3068 36740 3525 36768
rect 2869 36731 2927 36737
rect 3513 36737 3525 36740
rect 3559 36737 3571 36771
rect 3513 36731 3571 36737
rect 9030 36728 9036 36780
rect 9088 36768 9094 36780
rect 9309 36771 9367 36777
rect 9309 36768 9321 36771
rect 9088 36740 9321 36768
rect 9088 36728 9094 36740
rect 9309 36737 9321 36740
rect 9355 36737 9367 36771
rect 9309 36731 9367 36737
rect 10502 36728 10508 36780
rect 10560 36768 10566 36780
rect 10597 36771 10655 36777
rect 10597 36768 10609 36771
rect 10560 36740 10609 36768
rect 10560 36728 10566 36740
rect 10597 36737 10609 36740
rect 10643 36737 10655 36771
rect 19426 36768 19432 36780
rect 19387 36740 19432 36768
rect 10597 36731 10655 36737
rect 19426 36728 19432 36740
rect 19484 36728 19490 36780
rect 23290 36768 23296 36780
rect 23251 36740 23296 36768
rect 23290 36728 23296 36740
rect 23348 36728 23354 36780
rect 27341 36771 27399 36777
rect 27341 36737 27353 36771
rect 27387 36737 27399 36771
rect 35434 36768 35440 36780
rect 35395 36740 35440 36768
rect 27341 36731 27399 36737
rect 27356 36700 27384 36731
rect 35434 36728 35440 36740
rect 35492 36728 35498 36780
rect 35894 36728 35900 36780
rect 35952 36768 35958 36780
rect 36630 36768 36636 36780
rect 35952 36740 35997 36768
rect 36591 36740 36636 36768
rect 35952 36728 35958 36740
rect 36630 36728 36636 36740
rect 36688 36728 36694 36780
rect 37366 36728 37372 36780
rect 37424 36768 37430 36780
rect 37461 36771 37519 36777
rect 37461 36768 37473 36771
rect 37424 36740 37473 36768
rect 37424 36728 37430 36740
rect 37461 36737 37473 36740
rect 37507 36768 37519 36771
rect 38013 36771 38071 36777
rect 38013 36768 38025 36771
rect 37507 36740 38025 36768
rect 37507 36737 37519 36740
rect 37461 36731 37519 36737
rect 38013 36737 38025 36740
rect 38059 36737 38071 36771
rect 38013 36731 38071 36737
rect 27522 36700 27528 36712
rect 27356 36672 27528 36700
rect 27522 36660 27528 36672
rect 27580 36700 27586 36712
rect 37734 36700 37740 36712
rect 27580 36672 37740 36700
rect 27580 36660 27586 36672
rect 37734 36660 37740 36672
rect 37792 36660 37798 36712
rect 1854 36632 1860 36644
rect 1815 36604 1860 36632
rect 1854 36592 1860 36604
rect 1912 36592 1918 36644
rect 2685 36567 2743 36573
rect 2685 36533 2697 36567
rect 2731 36564 2743 36567
rect 3234 36564 3240 36576
rect 2731 36536 3240 36564
rect 2731 36533 2743 36536
rect 2685 36527 2743 36533
rect 3234 36524 3240 36536
rect 3292 36524 3298 36576
rect 3329 36567 3387 36573
rect 3329 36533 3341 36567
rect 3375 36564 3387 36567
rect 6546 36564 6552 36576
rect 3375 36536 6552 36564
rect 3375 36533 3387 36536
rect 3329 36527 3387 36533
rect 6546 36524 6552 36536
rect 6604 36524 6610 36576
rect 9125 36567 9183 36573
rect 9125 36533 9137 36567
rect 9171 36564 9183 36567
rect 9766 36564 9772 36576
rect 9171 36536 9772 36564
rect 9171 36533 9183 36536
rect 9125 36527 9183 36533
rect 9766 36524 9772 36536
rect 9824 36524 9830 36576
rect 32122 36524 32128 36576
rect 32180 36564 32186 36576
rect 35253 36567 35311 36573
rect 35253 36564 35265 36567
rect 32180 36536 35265 36564
rect 32180 36524 32186 36536
rect 35253 36533 35265 36536
rect 35299 36533 35311 36567
rect 35253 36527 35311 36533
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 1762 36360 1768 36372
rect 1723 36332 1768 36360
rect 1762 36320 1768 36332
rect 1820 36320 1826 36372
rect 36630 36360 36636 36372
rect 36591 36332 36636 36360
rect 36630 36320 36636 36332
rect 36688 36320 36694 36372
rect 1578 36156 1584 36168
rect 1539 36128 1584 36156
rect 1578 36116 1584 36128
rect 1636 36116 1642 36168
rect 2501 36159 2559 36165
rect 2501 36125 2513 36159
rect 2547 36156 2559 36159
rect 2866 36156 2872 36168
rect 2547 36128 2872 36156
rect 2547 36125 2559 36128
rect 2501 36119 2559 36125
rect 2866 36116 2872 36128
rect 2924 36116 2930 36168
rect 36814 36156 36820 36168
rect 36775 36128 36820 36156
rect 36814 36116 36820 36128
rect 36872 36116 36878 36168
rect 37182 36116 37188 36168
rect 37240 36156 37246 36168
rect 37369 36159 37427 36165
rect 37369 36156 37381 36159
rect 37240 36128 37381 36156
rect 37240 36116 37246 36128
rect 37369 36125 37381 36128
rect 37415 36125 37427 36159
rect 37369 36119 37427 36125
rect 37826 36116 37832 36168
rect 37884 36156 37890 36168
rect 38013 36159 38071 36165
rect 38013 36156 38025 36159
rect 37884 36128 38025 36156
rect 37884 36116 37890 36128
rect 38013 36125 38025 36128
rect 38059 36125 38071 36159
rect 38013 36119 38071 36125
rect 2317 36023 2375 36029
rect 2317 35989 2329 36023
rect 2363 36020 2375 36023
rect 6454 36020 6460 36032
rect 2363 35992 6460 36020
rect 2363 35989 2375 35992
rect 2317 35983 2375 35989
rect 6454 35980 6460 35992
rect 6512 35980 6518 36032
rect 37274 35980 37280 36032
rect 37332 36020 37338 36032
rect 37461 36023 37519 36029
rect 37461 36020 37473 36023
rect 37332 35992 37473 36020
rect 37332 35980 37338 35992
rect 37461 35989 37473 35992
rect 37507 35989 37519 36023
rect 38194 36020 38200 36032
rect 38155 35992 38200 36020
rect 37461 35983 37519 35989
rect 38194 35980 38200 35992
rect 38252 35980 38258 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 35529 35819 35587 35825
rect 35529 35785 35541 35819
rect 35575 35816 35587 35819
rect 36814 35816 36820 35828
rect 35575 35788 36820 35816
rect 35575 35785 35587 35788
rect 35529 35779 35587 35785
rect 36814 35776 36820 35788
rect 36872 35776 36878 35828
rect 1762 35680 1768 35692
rect 1723 35652 1768 35680
rect 1762 35640 1768 35652
rect 1820 35640 1826 35692
rect 14458 35640 14464 35692
rect 14516 35680 14522 35692
rect 35437 35683 35495 35689
rect 35437 35680 35449 35683
rect 14516 35652 35449 35680
rect 14516 35640 14522 35652
rect 35437 35649 35449 35652
rect 35483 35649 35495 35683
rect 38013 35683 38071 35689
rect 38013 35680 38025 35683
rect 35437 35643 35495 35649
rect 35866 35652 38025 35680
rect 32398 35572 32404 35624
rect 32456 35612 32462 35624
rect 35866 35612 35894 35652
rect 38013 35649 38025 35652
rect 38059 35649 38071 35683
rect 38013 35643 38071 35649
rect 32456 35584 35894 35612
rect 32456 35572 32462 35584
rect 1581 35479 1639 35485
rect 1581 35445 1593 35479
rect 1627 35476 1639 35479
rect 5534 35476 5540 35488
rect 1627 35448 5540 35476
rect 1627 35445 1639 35448
rect 1581 35439 1639 35445
rect 5534 35436 5540 35448
rect 5592 35436 5598 35488
rect 38194 35476 38200 35488
rect 38155 35448 38200 35476
rect 38194 35436 38200 35448
rect 38252 35436 38258 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 14737 35275 14795 35281
rect 14737 35241 14749 35275
rect 14783 35272 14795 35275
rect 16022 35272 16028 35284
rect 14783 35244 16028 35272
rect 14783 35241 14795 35244
rect 14737 35235 14795 35241
rect 16022 35232 16028 35244
rect 16080 35232 16086 35284
rect 13906 35028 13912 35080
rect 13964 35068 13970 35080
rect 14921 35071 14979 35077
rect 14921 35068 14933 35071
rect 13964 35040 14933 35068
rect 13964 35028 13970 35040
rect 14921 35037 14933 35040
rect 14967 35037 14979 35071
rect 14921 35031 14979 35037
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 1581 34595 1639 34601
rect 1581 34561 1593 34595
rect 1627 34592 1639 34595
rect 3050 34592 3056 34604
rect 1627 34564 3056 34592
rect 1627 34561 1639 34564
rect 1581 34555 1639 34561
rect 3050 34552 3056 34564
rect 3108 34552 3114 34604
rect 3234 34552 3240 34604
rect 3292 34592 3298 34604
rect 6549 34595 6607 34601
rect 6549 34592 6561 34595
rect 3292 34564 6561 34592
rect 3292 34552 3298 34564
rect 6549 34561 6561 34564
rect 6595 34561 6607 34595
rect 38010 34592 38016 34604
rect 37971 34564 38016 34592
rect 6549 34555 6607 34561
rect 38010 34552 38016 34564
rect 38068 34552 38074 34604
rect 6641 34527 6699 34533
rect 6641 34493 6653 34527
rect 6687 34524 6699 34527
rect 6730 34524 6736 34536
rect 6687 34496 6736 34524
rect 6687 34493 6699 34496
rect 6641 34487 6699 34493
rect 6730 34484 6736 34496
rect 6788 34484 6794 34536
rect 1762 34388 1768 34400
rect 1723 34360 1768 34388
rect 1762 34348 1768 34360
rect 1820 34348 1826 34400
rect 38194 34388 38200 34400
rect 38155 34360 38200 34388
rect 38194 34348 38200 34360
rect 38252 34348 38258 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 19426 33600 19432 33652
rect 19484 33640 19490 33652
rect 22097 33643 22155 33649
rect 22097 33640 22109 33643
rect 19484 33612 22109 33640
rect 19484 33600 19490 33612
rect 22097 33609 22109 33612
rect 22143 33609 22155 33643
rect 22097 33603 22155 33609
rect 11698 33464 11704 33516
rect 11756 33504 11762 33516
rect 15381 33507 15439 33513
rect 15381 33504 15393 33507
rect 11756 33476 15393 33504
rect 11756 33464 11762 33476
rect 15381 33473 15393 33476
rect 15427 33473 15439 33507
rect 15381 33467 15439 33473
rect 22281 33507 22339 33513
rect 22281 33473 22293 33507
rect 22327 33504 22339 33507
rect 24670 33504 24676 33516
rect 22327 33476 24676 33504
rect 22327 33473 22339 33476
rect 22281 33467 22339 33473
rect 24670 33464 24676 33476
rect 24728 33464 24734 33516
rect 15473 33303 15531 33309
rect 15473 33269 15485 33303
rect 15519 33300 15531 33303
rect 18598 33300 18604 33312
rect 15519 33272 18604 33300
rect 15519 33269 15531 33272
rect 15473 33263 15531 33269
rect 18598 33260 18604 33272
rect 18656 33260 18662 33312
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 32125 33099 32183 33105
rect 32125 33065 32137 33099
rect 32171 33096 32183 33099
rect 35986 33096 35992 33108
rect 32171 33068 35992 33096
rect 32171 33065 32183 33068
rect 32125 33059 32183 33065
rect 35986 33056 35992 33068
rect 36044 33056 36050 33108
rect 1581 32895 1639 32901
rect 1581 32861 1593 32895
rect 1627 32892 1639 32895
rect 2498 32892 2504 32904
rect 1627 32864 2360 32892
rect 2459 32864 2504 32892
rect 1627 32861 1639 32864
rect 1581 32855 1639 32861
rect 1762 32756 1768 32768
rect 1723 32728 1768 32756
rect 1762 32716 1768 32728
rect 1820 32716 1826 32768
rect 2332 32765 2360 32864
rect 2498 32852 2504 32864
rect 2556 32852 2562 32904
rect 31110 32852 31116 32904
rect 31168 32892 31174 32904
rect 32309 32895 32367 32901
rect 32309 32892 32321 32895
rect 31168 32864 32321 32892
rect 31168 32852 31174 32864
rect 32309 32861 32321 32864
rect 32355 32861 32367 32895
rect 37458 32892 37464 32904
rect 37419 32864 37464 32892
rect 32309 32855 32367 32861
rect 37458 32852 37464 32864
rect 37516 32852 37522 32904
rect 37737 32895 37795 32901
rect 37737 32861 37749 32895
rect 37783 32892 37795 32895
rect 38378 32892 38384 32904
rect 37783 32864 38384 32892
rect 37783 32861 37795 32864
rect 37737 32855 37795 32861
rect 38378 32852 38384 32864
rect 38436 32852 38442 32904
rect 2317 32759 2375 32765
rect 2317 32725 2329 32759
rect 2363 32725 2375 32759
rect 2317 32719 2375 32725
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 29641 32555 29699 32561
rect 29641 32521 29653 32555
rect 29687 32552 29699 32555
rect 33226 32552 33232 32564
rect 29687 32524 33232 32552
rect 29687 32521 29699 32524
rect 29641 32515 29699 32521
rect 33226 32512 33232 32524
rect 33284 32512 33290 32564
rect 1581 32419 1639 32425
rect 1581 32385 1593 32419
rect 1627 32416 1639 32419
rect 1854 32416 1860 32428
rect 1627 32388 1860 32416
rect 1627 32385 1639 32388
rect 1581 32379 1639 32385
rect 1854 32376 1860 32388
rect 1912 32376 1918 32428
rect 29638 32376 29644 32428
rect 29696 32416 29702 32428
rect 29825 32419 29883 32425
rect 29825 32416 29837 32419
rect 29696 32388 29837 32416
rect 29696 32376 29702 32388
rect 29825 32385 29837 32388
rect 29871 32385 29883 32419
rect 38286 32416 38292 32428
rect 38247 32388 38292 32416
rect 29825 32379 29883 32385
rect 38286 32376 38292 32388
rect 38344 32376 38350 32428
rect 25682 32240 25688 32292
rect 25740 32280 25746 32292
rect 29730 32280 29736 32292
rect 25740 32252 29736 32280
rect 25740 32240 25746 32252
rect 29730 32240 29736 32252
rect 29788 32240 29794 32292
rect 1762 32212 1768 32224
rect 1723 32184 1768 32212
rect 1762 32172 1768 32184
rect 1820 32172 1826 32224
rect 37642 32172 37648 32224
rect 37700 32212 37706 32224
rect 38105 32215 38163 32221
rect 38105 32212 38117 32215
rect 37700 32184 38117 32212
rect 37700 32172 37706 32184
rect 38105 32181 38117 32184
rect 38151 32181 38163 32215
rect 38105 32175 38163 32181
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 22281 32011 22339 32017
rect 22281 31977 22293 32011
rect 22327 32008 22339 32011
rect 23290 32008 23296 32020
rect 22327 31980 23296 32008
rect 22327 31977 22339 31980
rect 22281 31971 22339 31977
rect 23290 31968 23296 31980
rect 23348 31968 23354 32020
rect 27982 32008 27988 32020
rect 27943 31980 27988 32008
rect 27982 31968 27988 31980
rect 28040 31968 28046 32020
rect 31110 32008 31116 32020
rect 31071 31980 31116 32008
rect 31110 31968 31116 31980
rect 31168 31968 31174 32020
rect 36909 32011 36967 32017
rect 36909 31977 36921 32011
rect 36955 32008 36967 32011
rect 38010 32008 38016 32020
rect 36955 31980 38016 32008
rect 36955 31977 36967 31980
rect 36909 31971 36967 31977
rect 38010 31968 38016 31980
rect 38068 31968 38074 32020
rect 23198 31900 23204 31952
rect 23256 31940 23262 31952
rect 23256 31912 31064 31940
rect 23256 31900 23262 31912
rect 21266 31832 21272 31884
rect 21324 31872 21330 31884
rect 25777 31875 25835 31881
rect 25777 31872 25789 31875
rect 21324 31844 25789 31872
rect 21324 31832 21330 31844
rect 25777 31841 25789 31844
rect 25823 31841 25835 31875
rect 25777 31835 25835 31841
rect 27246 31832 27252 31884
rect 27304 31872 27310 31884
rect 27433 31875 27491 31881
rect 27433 31872 27445 31875
rect 27304 31844 27445 31872
rect 27304 31832 27310 31844
rect 27433 31841 27445 31844
rect 27479 31841 27491 31875
rect 30374 31872 30380 31884
rect 27433 31835 27491 31841
rect 28092 31844 30380 31872
rect 7926 31804 7932 31816
rect 7887 31776 7932 31804
rect 7926 31764 7932 31776
rect 7984 31764 7990 31816
rect 8021 31807 8079 31813
rect 8021 31773 8033 31807
rect 8067 31804 8079 31807
rect 8110 31804 8116 31816
rect 8067 31776 8116 31804
rect 8067 31773 8079 31776
rect 8021 31767 8079 31773
rect 8110 31764 8116 31776
rect 8168 31764 8174 31816
rect 21542 31764 21548 31816
rect 21600 31804 21606 31816
rect 22465 31807 22523 31813
rect 22465 31804 22477 31807
rect 21600 31776 22477 31804
rect 21600 31764 21606 31776
rect 22465 31773 22477 31776
rect 22511 31773 22523 31807
rect 25682 31804 25688 31816
rect 25643 31776 25688 31804
rect 22465 31767 22523 31773
rect 25682 31764 25688 31776
rect 25740 31764 25746 31816
rect 26878 31764 26884 31816
rect 26936 31804 26942 31816
rect 27341 31807 27399 31813
rect 26936 31776 27292 31804
rect 26936 31764 26942 31776
rect 27264 31736 27292 31776
rect 27341 31773 27353 31807
rect 27387 31804 27399 31807
rect 28092 31804 28120 31844
rect 30374 31832 30380 31844
rect 30432 31832 30438 31884
rect 31036 31813 31064 31912
rect 27387 31776 28120 31804
rect 28169 31807 28227 31813
rect 27387 31773 27399 31776
rect 27341 31767 27399 31773
rect 28169 31773 28181 31807
rect 28215 31773 28227 31807
rect 28169 31767 28227 31773
rect 31021 31807 31079 31813
rect 31021 31773 31033 31807
rect 31067 31773 31079 31807
rect 37090 31804 37096 31816
rect 37051 31776 37096 31804
rect 31021 31767 31079 31773
rect 28184 31736 28212 31767
rect 37090 31764 37096 31776
rect 37148 31764 37154 31816
rect 27264 31708 28212 31736
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 32493 31467 32551 31473
rect 32493 31433 32505 31467
rect 32539 31464 32551 31467
rect 35894 31464 35900 31476
rect 32539 31436 35900 31464
rect 32539 31433 32551 31436
rect 32493 31427 32551 31433
rect 35894 31424 35900 31436
rect 35952 31424 35958 31476
rect 6178 31356 6184 31408
rect 6236 31396 6242 31408
rect 6236 31368 7236 31396
rect 6236 31356 6242 31368
rect 6546 31328 6552 31340
rect 6507 31300 6552 31328
rect 6546 31288 6552 31300
rect 6604 31288 6610 31340
rect 7208 31337 7236 31368
rect 7193 31331 7251 31337
rect 7193 31297 7205 31331
rect 7239 31297 7251 31331
rect 7193 31291 7251 31297
rect 16853 31331 16911 31337
rect 16853 31297 16865 31331
rect 16899 31328 16911 31331
rect 17126 31328 17132 31340
rect 16899 31300 17132 31328
rect 16899 31297 16911 31300
rect 16853 31291 16911 31297
rect 17126 31288 17132 31300
rect 17184 31288 17190 31340
rect 30374 31288 30380 31340
rect 30432 31328 30438 31340
rect 32677 31331 32735 31337
rect 32677 31328 32689 31331
rect 30432 31300 32689 31328
rect 30432 31288 30438 31300
rect 32677 31297 32689 31300
rect 32723 31297 32735 31331
rect 32677 31291 32735 31297
rect 6641 31127 6699 31133
rect 6641 31093 6653 31127
rect 6687 31124 6699 31127
rect 6822 31124 6828 31136
rect 6687 31096 6828 31124
rect 6687 31093 6699 31096
rect 6641 31087 6699 31093
rect 6822 31084 6828 31096
rect 6880 31084 6886 31136
rect 7285 31127 7343 31133
rect 7285 31093 7297 31127
rect 7331 31124 7343 31127
rect 7374 31124 7380 31136
rect 7331 31096 7380 31124
rect 7331 31093 7343 31096
rect 7285 31087 7343 31093
rect 7374 31084 7380 31096
rect 7432 31084 7438 31136
rect 15470 31084 15476 31136
rect 15528 31124 15534 31136
rect 16945 31127 17003 31133
rect 16945 31124 16957 31127
rect 15528 31096 16957 31124
rect 15528 31084 15534 31096
rect 16945 31093 16957 31096
rect 16991 31093 17003 31127
rect 16945 31087 17003 31093
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 3050 30880 3056 30932
rect 3108 30920 3114 30932
rect 3973 30923 4031 30929
rect 3973 30920 3985 30923
rect 3108 30892 3985 30920
rect 3108 30880 3114 30892
rect 3973 30889 3985 30892
rect 4019 30889 4031 30923
rect 3973 30883 4031 30889
rect 36265 30923 36323 30929
rect 36265 30889 36277 30923
rect 36311 30920 36323 30923
rect 37090 30920 37096 30932
rect 36311 30892 37096 30920
rect 36311 30889 36323 30892
rect 36265 30883 36323 30889
rect 37090 30880 37096 30892
rect 37148 30880 37154 30932
rect 24578 30784 24584 30796
rect 22066 30756 24584 30784
rect 1581 30719 1639 30725
rect 1581 30685 1593 30719
rect 1627 30685 1639 30719
rect 1581 30679 1639 30685
rect 4157 30719 4215 30725
rect 4157 30685 4169 30719
rect 4203 30716 4215 30719
rect 8478 30716 8484 30728
rect 4203 30688 8484 30716
rect 4203 30685 4215 30688
rect 4157 30679 4215 30685
rect 1596 30648 1624 30679
rect 8478 30676 8484 30688
rect 8536 30676 8542 30728
rect 9950 30676 9956 30728
rect 10008 30716 10014 30728
rect 10413 30719 10471 30725
rect 10413 30716 10425 30719
rect 10008 30688 10425 30716
rect 10008 30676 10014 30688
rect 10413 30685 10425 30688
rect 10459 30685 10471 30719
rect 10413 30679 10471 30685
rect 21821 30719 21879 30725
rect 21821 30685 21833 30719
rect 21867 30716 21879 30719
rect 22066 30716 22094 30756
rect 24578 30744 24584 30756
rect 24636 30744 24642 30796
rect 21867 30688 22094 30716
rect 22649 30719 22707 30725
rect 21867 30685 21879 30688
rect 21821 30679 21879 30685
rect 22649 30685 22661 30719
rect 22695 30716 22707 30719
rect 25866 30716 25872 30728
rect 22695 30688 25872 30716
rect 22695 30685 22707 30688
rect 22649 30679 22707 30685
rect 25866 30676 25872 30688
rect 25924 30676 25930 30728
rect 27985 30719 28043 30725
rect 27985 30685 27997 30719
rect 28031 30716 28043 30719
rect 32122 30716 32128 30728
rect 28031 30688 32128 30716
rect 28031 30685 28043 30688
rect 27985 30679 28043 30685
rect 32122 30676 32128 30688
rect 32180 30676 32186 30728
rect 36170 30716 36176 30728
rect 36131 30688 36176 30716
rect 36170 30676 36176 30688
rect 36228 30676 36234 30728
rect 38286 30716 38292 30728
rect 38247 30688 38292 30716
rect 38286 30676 38292 30688
rect 38344 30676 38350 30728
rect 6270 30648 6276 30660
rect 1596 30620 6276 30648
rect 6270 30608 6276 30620
rect 6328 30608 6334 30660
rect 18414 30608 18420 30660
rect 18472 30648 18478 30660
rect 22741 30651 22799 30657
rect 22741 30648 22753 30651
rect 18472 30620 22753 30648
rect 18472 30608 18478 30620
rect 22741 30617 22753 30620
rect 22787 30617 22799 30651
rect 22741 30611 22799 30617
rect 1762 30580 1768 30592
rect 1723 30552 1768 30580
rect 1762 30540 1768 30552
rect 1820 30540 1826 30592
rect 10226 30540 10232 30592
rect 10284 30580 10290 30592
rect 10505 30583 10563 30589
rect 10505 30580 10517 30583
rect 10284 30552 10517 30580
rect 10284 30540 10290 30552
rect 10505 30549 10517 30552
rect 10551 30549 10563 30583
rect 21910 30580 21916 30592
rect 21871 30552 21916 30580
rect 10505 30543 10563 30549
rect 21910 30540 21916 30552
rect 21968 30540 21974 30592
rect 28074 30580 28080 30592
rect 28035 30552 28080 30580
rect 28074 30540 28080 30552
rect 28132 30540 28138 30592
rect 38010 30540 38016 30592
rect 38068 30580 38074 30592
rect 38105 30583 38163 30589
rect 38105 30580 38117 30583
rect 38068 30552 38117 30580
rect 38068 30540 38074 30552
rect 38105 30549 38117 30552
rect 38151 30549 38163 30583
rect 38105 30543 38163 30549
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 17954 30336 17960 30388
rect 18012 30376 18018 30388
rect 28074 30376 28080 30388
rect 18012 30348 28080 30376
rect 18012 30336 18018 30348
rect 28074 30336 28080 30348
rect 28132 30336 28138 30388
rect 13906 30308 13912 30320
rect 13867 30280 13912 30308
rect 13906 30268 13912 30280
rect 13964 30268 13970 30320
rect 27430 30308 27436 30320
rect 23400 30280 27436 30308
rect 6454 30200 6460 30252
rect 6512 30240 6518 30252
rect 6549 30243 6607 30249
rect 6549 30240 6561 30243
rect 6512 30212 6561 30240
rect 6512 30200 6518 30212
rect 6549 30209 6561 30212
rect 6595 30209 6607 30243
rect 6549 30203 6607 30209
rect 13446 30200 13452 30252
rect 13504 30240 13510 30252
rect 13817 30243 13875 30249
rect 13817 30240 13829 30243
rect 13504 30212 13829 30240
rect 13504 30200 13510 30212
rect 13817 30209 13829 30212
rect 13863 30209 13875 30243
rect 13817 30203 13875 30209
rect 14461 30243 14519 30249
rect 14461 30209 14473 30243
rect 14507 30240 14519 30243
rect 15010 30240 15016 30252
rect 14507 30212 15016 30240
rect 14507 30209 14519 30212
rect 14461 30203 14519 30209
rect 15010 30200 15016 30212
rect 15068 30200 15074 30252
rect 23400 30249 23428 30280
rect 27430 30268 27436 30280
rect 27488 30268 27494 30320
rect 29638 30308 29644 30320
rect 29599 30280 29644 30308
rect 29638 30268 29644 30280
rect 29696 30268 29702 30320
rect 23385 30243 23443 30249
rect 23385 30209 23397 30243
rect 23431 30209 23443 30243
rect 23385 30203 23443 30209
rect 26237 30243 26295 30249
rect 26237 30209 26249 30243
rect 26283 30209 26295 30243
rect 29546 30240 29552 30252
rect 29507 30212 29552 30240
rect 26237 30203 26295 30209
rect 26252 30172 26280 30203
rect 29546 30200 29552 30212
rect 29604 30200 29610 30252
rect 37734 30200 37740 30252
rect 37792 30240 37798 30252
rect 38013 30243 38071 30249
rect 38013 30240 38025 30243
rect 37792 30212 38025 30240
rect 37792 30200 37798 30212
rect 38013 30209 38025 30212
rect 38059 30209 38071 30243
rect 38013 30203 38071 30209
rect 31294 30172 31300 30184
rect 26252 30144 31300 30172
rect 31294 30132 31300 30144
rect 31352 30132 31358 30184
rect 15562 30064 15568 30116
rect 15620 30104 15626 30116
rect 26329 30107 26387 30113
rect 26329 30104 26341 30107
rect 15620 30076 26341 30104
rect 15620 30064 15626 30076
rect 26329 30073 26341 30076
rect 26375 30073 26387 30107
rect 37826 30104 37832 30116
rect 37787 30076 37832 30104
rect 26329 30067 26387 30073
rect 37826 30064 37832 30076
rect 37884 30064 37890 30116
rect 6638 30036 6644 30048
rect 6599 30008 6644 30036
rect 6638 29996 6644 30008
rect 6696 29996 6702 30048
rect 13078 29996 13084 30048
rect 13136 30036 13142 30048
rect 14553 30039 14611 30045
rect 14553 30036 14565 30039
rect 13136 30008 14565 30036
rect 13136 29996 13142 30008
rect 14553 30005 14565 30008
rect 14599 30005 14611 30039
rect 14553 29999 14611 30005
rect 23477 30039 23535 30045
rect 23477 30005 23489 30039
rect 23523 30036 23535 30039
rect 23566 30036 23572 30048
rect 23523 30008 23572 30036
rect 23523 30005 23535 30008
rect 23477 29999 23535 30005
rect 23566 29996 23572 30008
rect 23624 29996 23630 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 21542 29832 21548 29844
rect 21503 29804 21548 29832
rect 21542 29792 21548 29804
rect 21600 29792 21606 29844
rect 29825 29835 29883 29841
rect 29825 29801 29837 29835
rect 29871 29832 29883 29835
rect 30374 29832 30380 29844
rect 29871 29804 30380 29832
rect 29871 29801 29883 29804
rect 29825 29795 29883 29801
rect 30374 29792 30380 29804
rect 30432 29792 30438 29844
rect 1486 29588 1492 29640
rect 1544 29628 1550 29640
rect 1581 29631 1639 29637
rect 1581 29628 1593 29631
rect 1544 29600 1593 29628
rect 1544 29588 1550 29600
rect 1581 29597 1593 29600
rect 1627 29597 1639 29631
rect 1581 29591 1639 29597
rect 9766 29588 9772 29640
rect 9824 29628 9830 29640
rect 11425 29631 11483 29637
rect 11425 29628 11437 29631
rect 9824 29600 11437 29628
rect 9824 29588 9830 29600
rect 11425 29597 11437 29600
rect 11471 29597 11483 29631
rect 11425 29591 11483 29597
rect 15010 29588 15016 29640
rect 15068 29628 15074 29640
rect 21453 29631 21511 29637
rect 21453 29628 21465 29631
rect 15068 29600 21465 29628
rect 15068 29588 15074 29600
rect 21453 29597 21465 29600
rect 21499 29597 21511 29631
rect 21453 29591 21511 29597
rect 27154 29588 27160 29640
rect 27212 29628 27218 29640
rect 29733 29631 29791 29637
rect 29733 29628 29745 29631
rect 27212 29600 29745 29628
rect 27212 29588 27218 29600
rect 29733 29597 29745 29600
rect 29779 29597 29791 29631
rect 29733 29591 29791 29597
rect 38102 29560 38108 29572
rect 38063 29532 38108 29560
rect 38102 29520 38108 29532
rect 38160 29520 38166 29572
rect 1762 29492 1768 29504
rect 1723 29464 1768 29492
rect 1762 29452 1768 29464
rect 1820 29452 1826 29504
rect 11422 29452 11428 29504
rect 11480 29492 11486 29504
rect 11517 29495 11575 29501
rect 11517 29492 11529 29495
rect 11480 29464 11529 29492
rect 11480 29452 11486 29464
rect 11517 29461 11529 29464
rect 11563 29461 11575 29495
rect 38194 29492 38200 29504
rect 38155 29464 38200 29492
rect 11517 29455 11575 29461
rect 38194 29452 38200 29464
rect 38252 29452 38258 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 21174 29248 21180 29300
rect 21232 29288 21238 29300
rect 22005 29291 22063 29297
rect 22005 29288 22017 29291
rect 21232 29260 22017 29288
rect 21232 29248 21238 29260
rect 22005 29257 22017 29260
rect 22051 29257 22063 29291
rect 22005 29251 22063 29257
rect 1762 29152 1768 29164
rect 1723 29124 1768 29152
rect 1762 29112 1768 29124
rect 1820 29112 1826 29164
rect 10502 29112 10508 29164
rect 10560 29152 10566 29164
rect 11977 29155 12035 29161
rect 11977 29152 11989 29155
rect 10560 29124 11989 29152
rect 10560 29112 10566 29124
rect 11977 29121 11989 29124
rect 12023 29121 12035 29155
rect 11977 29115 12035 29121
rect 22094 29112 22100 29164
rect 22152 29152 22158 29164
rect 22189 29155 22247 29161
rect 22189 29152 22201 29155
rect 22152 29124 22201 29152
rect 22152 29112 22158 29124
rect 22189 29121 22201 29124
rect 22235 29121 22247 29155
rect 38286 29152 38292 29164
rect 38247 29124 38292 29152
rect 22189 29115 22247 29121
rect 38286 29112 38292 29124
rect 38344 29112 38350 29164
rect 1581 29019 1639 29025
rect 1581 28985 1593 29019
rect 1627 29016 1639 29019
rect 1946 29016 1952 29028
rect 1627 28988 1952 29016
rect 1627 28985 1639 28988
rect 1581 28979 1639 28985
rect 1946 28976 1952 28988
rect 2004 28976 2010 29028
rect 11330 28976 11336 29028
rect 11388 29016 11394 29028
rect 12069 29019 12127 29025
rect 12069 29016 12081 29019
rect 11388 28988 12081 29016
rect 11388 28976 11394 28988
rect 12069 28985 12081 28988
rect 12115 28985 12127 29019
rect 12069 28979 12127 28985
rect 17586 28976 17592 29028
rect 17644 29016 17650 29028
rect 21910 29016 21916 29028
rect 17644 28988 21916 29016
rect 17644 28976 17650 28988
rect 21910 28976 21916 28988
rect 21968 28976 21974 29028
rect 37918 28976 37924 29028
rect 37976 29016 37982 29028
rect 38105 29019 38163 29025
rect 38105 29016 38117 29019
rect 37976 28988 38117 29016
rect 37976 28976 37982 28988
rect 38105 28985 38117 28988
rect 38151 28985 38163 29019
rect 38105 28979 38163 28985
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 6270 28744 6276 28756
rect 6231 28716 6276 28744
rect 6270 28704 6276 28716
rect 6328 28704 6334 28756
rect 6457 28543 6515 28549
rect 6457 28509 6469 28543
rect 6503 28540 6515 28543
rect 8202 28540 8208 28552
rect 6503 28512 8208 28540
rect 6503 28509 6515 28512
rect 6457 28503 6515 28509
rect 8202 28500 8208 28512
rect 8260 28500 8266 28552
rect 10318 28500 10324 28552
rect 10376 28540 10382 28552
rect 11701 28543 11759 28549
rect 11701 28540 11713 28543
rect 10376 28512 11713 28540
rect 10376 28500 10382 28512
rect 11701 28509 11713 28512
rect 11747 28509 11759 28543
rect 27522 28540 27528 28552
rect 27483 28512 27528 28540
rect 11701 28503 11759 28509
rect 27522 28500 27528 28512
rect 27580 28500 27586 28552
rect 11514 28404 11520 28416
rect 11475 28376 11520 28404
rect 11514 28364 11520 28376
rect 11572 28364 11578 28416
rect 27617 28407 27675 28413
rect 27617 28373 27629 28407
rect 27663 28404 27675 28407
rect 27798 28404 27804 28416
rect 27663 28376 27804 28404
rect 27663 28373 27675 28376
rect 27617 28367 27675 28373
rect 27798 28364 27804 28376
rect 27856 28364 27862 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 10318 28200 10324 28212
rect 10279 28172 10324 28200
rect 10318 28160 10324 28172
rect 10376 28160 10382 28212
rect 5534 28024 5540 28076
rect 5592 28064 5598 28076
rect 9125 28067 9183 28073
rect 9125 28064 9137 28067
rect 5592 28036 9137 28064
rect 5592 28024 5598 28036
rect 9125 28033 9137 28036
rect 9171 28033 9183 28067
rect 9125 28027 9183 28033
rect 10505 28067 10563 28073
rect 10505 28033 10517 28067
rect 10551 28033 10563 28067
rect 11146 28064 11152 28076
rect 11107 28036 11152 28064
rect 10505 28027 10563 28033
rect 10520 27996 10548 28027
rect 11146 28024 11152 28036
rect 11204 28024 11210 28076
rect 11793 28067 11851 28073
rect 11793 28033 11805 28067
rect 11839 28033 11851 28067
rect 11793 28027 11851 28033
rect 11606 27996 11612 28008
rect 10520 27968 11612 27996
rect 11606 27956 11612 27968
rect 11664 27996 11670 28008
rect 11808 27996 11836 28027
rect 11974 28024 11980 28076
rect 12032 28064 12038 28076
rect 12621 28067 12679 28073
rect 12621 28064 12633 28067
rect 12032 28036 12633 28064
rect 12032 28024 12038 28036
rect 12621 28033 12633 28036
rect 12667 28033 12679 28067
rect 12621 28027 12679 28033
rect 12986 28024 12992 28076
rect 13044 28064 13050 28076
rect 13449 28067 13507 28073
rect 13449 28064 13461 28067
rect 13044 28036 13461 28064
rect 13044 28024 13050 28036
rect 13449 28033 13461 28036
rect 13495 28033 13507 28067
rect 13449 28027 13507 28033
rect 11664 27968 11836 27996
rect 11664 27956 11670 27968
rect 10965 27931 11023 27937
rect 10965 27897 10977 27931
rect 11011 27928 11023 27931
rect 12066 27928 12072 27940
rect 11011 27900 12072 27928
rect 11011 27897 11023 27900
rect 10965 27891 11023 27897
rect 12066 27888 12072 27900
rect 12124 27888 12130 27940
rect 9214 27860 9220 27872
rect 9175 27832 9220 27860
rect 9214 27820 9220 27832
rect 9272 27820 9278 27872
rect 11882 27860 11888 27872
rect 11843 27832 11888 27860
rect 11882 27820 11888 27832
rect 11940 27820 11946 27872
rect 12710 27860 12716 27872
rect 12671 27832 12716 27860
rect 12710 27820 12716 27832
rect 12768 27820 12774 27872
rect 13262 27860 13268 27872
rect 13223 27832 13268 27860
rect 13262 27820 13268 27832
rect 13320 27820 13326 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 9214 27616 9220 27668
rect 9272 27656 9278 27668
rect 21818 27656 21824 27668
rect 9272 27628 21824 27656
rect 9272 27616 9278 27628
rect 21818 27616 21824 27628
rect 21876 27616 21882 27668
rect 10413 27591 10471 27597
rect 10413 27557 10425 27591
rect 10459 27588 10471 27591
rect 11146 27588 11152 27600
rect 10459 27560 11152 27588
rect 10459 27557 10471 27560
rect 10413 27551 10471 27557
rect 11146 27548 11152 27560
rect 11204 27548 11210 27600
rect 13446 27588 13452 27600
rect 13407 27560 13452 27588
rect 13446 27548 13452 27560
rect 13504 27548 13510 27600
rect 17678 27548 17684 27600
rect 17736 27588 17742 27600
rect 25498 27588 25504 27600
rect 17736 27560 25504 27588
rect 17736 27548 17742 27560
rect 25498 27548 25504 27560
rect 25556 27548 25562 27600
rect 11882 27520 11888 27532
rect 11843 27492 11888 27520
rect 11882 27480 11888 27492
rect 11940 27480 11946 27532
rect 12526 27520 12532 27532
rect 11992 27492 12532 27520
rect 1578 27452 1584 27464
rect 1539 27424 1584 27452
rect 1578 27412 1584 27424
rect 1636 27412 1642 27464
rect 1857 27455 1915 27461
rect 1857 27421 1869 27455
rect 1903 27452 1915 27455
rect 5534 27452 5540 27464
rect 1903 27424 5540 27452
rect 1903 27421 1915 27424
rect 1857 27415 1915 27421
rect 5534 27412 5540 27424
rect 5592 27412 5598 27464
rect 10597 27455 10655 27461
rect 10597 27421 10609 27455
rect 10643 27421 10655 27455
rect 10597 27415 10655 27421
rect 11057 27455 11115 27461
rect 11057 27421 11069 27455
rect 11103 27421 11115 27455
rect 11057 27415 11115 27421
rect 11149 27455 11207 27461
rect 11149 27421 11161 27455
rect 11195 27452 11207 27455
rect 11701 27455 11759 27461
rect 11701 27452 11713 27455
rect 11195 27424 11713 27452
rect 11195 27421 11207 27424
rect 11149 27415 11207 27421
rect 11701 27421 11713 27424
rect 11747 27452 11759 27455
rect 11992 27452 12020 27492
rect 12526 27480 12532 27492
rect 12584 27480 12590 27532
rect 12710 27480 12716 27532
rect 12768 27520 12774 27532
rect 12989 27523 13047 27529
rect 12989 27520 13001 27523
rect 12768 27492 13001 27520
rect 12768 27480 12774 27492
rect 12989 27489 13001 27492
rect 13035 27489 13047 27523
rect 38194 27520 38200 27532
rect 12989 27483 13047 27489
rect 22066 27492 38200 27520
rect 11747 27424 12020 27452
rect 12345 27455 12403 27461
rect 11747 27421 11759 27424
rect 11701 27415 11759 27421
rect 12345 27421 12357 27455
rect 12391 27452 12403 27455
rect 12434 27452 12440 27464
rect 12391 27424 12440 27452
rect 12391 27421 12403 27424
rect 12345 27415 12403 27421
rect 10612 27316 10640 27415
rect 10962 27344 10968 27396
rect 11020 27384 11026 27396
rect 11072 27384 11100 27415
rect 12434 27412 12440 27424
rect 12492 27452 12498 27464
rect 12805 27455 12863 27461
rect 12805 27452 12817 27455
rect 12492 27424 12817 27452
rect 12492 27412 12498 27424
rect 12805 27421 12817 27424
rect 12851 27421 12863 27455
rect 12805 27415 12863 27421
rect 22066 27384 22094 27492
rect 38194 27480 38200 27492
rect 38252 27480 38258 27532
rect 38286 27452 38292 27464
rect 38247 27424 38292 27452
rect 38286 27412 38292 27424
rect 38344 27412 38350 27464
rect 11020 27356 22094 27384
rect 11020 27344 11026 27356
rect 11146 27316 11152 27328
rect 10612 27288 11152 27316
rect 11146 27276 11152 27288
rect 11204 27316 11210 27328
rect 11974 27316 11980 27328
rect 11204 27288 11980 27316
rect 11204 27276 11210 27288
rect 11974 27276 11980 27288
rect 12032 27276 12038 27328
rect 14734 27316 14740 27328
rect 14695 27288 14740 27316
rect 14734 27276 14740 27288
rect 14792 27276 14798 27328
rect 34606 27276 34612 27328
rect 34664 27316 34670 27328
rect 38105 27319 38163 27325
rect 38105 27316 38117 27319
rect 34664 27288 38117 27316
rect 34664 27276 34670 27288
rect 38105 27285 38117 27288
rect 38151 27285 38163 27319
rect 38105 27279 38163 27285
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 12434 27072 12440 27124
rect 12492 27112 12498 27124
rect 12492 27084 12537 27112
rect 12492 27072 12498 27084
rect 13446 27072 13452 27124
rect 13504 27112 13510 27124
rect 13541 27115 13599 27121
rect 13541 27112 13553 27115
rect 13504 27084 13553 27112
rect 13504 27072 13510 27084
rect 13541 27081 13553 27084
rect 13587 27081 13599 27115
rect 13541 27075 13599 27081
rect 22465 27115 22523 27121
rect 22465 27081 22477 27115
rect 22511 27081 22523 27115
rect 22465 27075 22523 27081
rect 10962 27044 10968 27056
rect 10923 27016 10968 27044
rect 10962 27004 10968 27016
rect 11020 27004 11026 27056
rect 12250 27044 12256 27056
rect 11440 27016 12256 27044
rect 10042 26936 10048 26988
rect 10100 26976 10106 26988
rect 10413 26979 10471 26985
rect 10413 26976 10425 26979
rect 10100 26948 10425 26976
rect 10100 26936 10106 26948
rect 10413 26945 10425 26948
rect 10459 26945 10471 26979
rect 10413 26939 10471 26945
rect 9398 26868 9404 26920
rect 9456 26908 9462 26920
rect 11440 26908 11468 27016
rect 12250 27004 12256 27016
rect 12308 27004 12314 27056
rect 22480 27044 22508 27075
rect 22480 27016 23336 27044
rect 11514 26936 11520 26988
rect 11572 26976 11578 26988
rect 11977 26979 12035 26985
rect 11977 26976 11989 26979
rect 11572 26948 11989 26976
rect 11572 26936 11578 26948
rect 11977 26945 11989 26948
rect 12023 26945 12035 26979
rect 11977 26939 12035 26945
rect 12066 26936 12072 26988
rect 12124 26976 12130 26988
rect 13081 26979 13139 26985
rect 13081 26976 13093 26979
rect 12124 26948 13093 26976
rect 12124 26936 12130 26948
rect 13081 26945 13093 26948
rect 13127 26945 13139 26979
rect 13081 26939 13139 26945
rect 13998 26936 14004 26988
rect 14056 26976 14062 26988
rect 14737 26979 14795 26985
rect 14737 26976 14749 26979
rect 14056 26948 14749 26976
rect 14056 26936 14062 26948
rect 14737 26945 14749 26948
rect 14783 26945 14795 26979
rect 15378 26976 15384 26988
rect 15339 26948 15384 26976
rect 14737 26939 14795 26945
rect 15378 26936 15384 26948
rect 15436 26936 15442 26988
rect 21910 26936 21916 26988
rect 21968 26976 21974 26988
rect 23308 26985 23336 27016
rect 22649 26979 22707 26985
rect 22649 26976 22661 26979
rect 21968 26948 22661 26976
rect 21968 26936 21974 26948
rect 22649 26945 22661 26948
rect 22695 26945 22707 26979
rect 22649 26939 22707 26945
rect 23293 26979 23351 26985
rect 23293 26945 23305 26979
rect 23339 26945 23351 26979
rect 23293 26939 23351 26945
rect 11790 26908 11796 26920
rect 9456 26880 11468 26908
rect 11751 26880 11796 26908
rect 9456 26868 9462 26880
rect 11790 26868 11796 26880
rect 11848 26868 11854 26920
rect 12894 26908 12900 26920
rect 12855 26880 12900 26908
rect 12894 26868 12900 26880
rect 12952 26868 12958 26920
rect 10229 26843 10287 26849
rect 10229 26809 10241 26843
rect 10275 26840 10287 26843
rect 12802 26840 12808 26852
rect 10275 26812 12808 26840
rect 10275 26809 10287 26812
rect 10229 26803 10287 26809
rect 12802 26800 12808 26812
rect 12860 26800 12866 26852
rect 11054 26772 11060 26784
rect 11015 26744 11060 26772
rect 11054 26732 11060 26744
rect 11112 26732 11118 26784
rect 14550 26772 14556 26784
rect 14511 26744 14556 26772
rect 14550 26732 14556 26744
rect 14608 26732 14614 26784
rect 15194 26772 15200 26784
rect 15155 26744 15200 26772
rect 15194 26732 15200 26744
rect 15252 26732 15258 26784
rect 23109 26775 23167 26781
rect 23109 26741 23121 26775
rect 23155 26772 23167 26775
rect 23290 26772 23296 26784
rect 23155 26744 23296 26772
rect 23155 26741 23167 26744
rect 23109 26735 23167 26741
rect 23290 26732 23296 26744
rect 23348 26732 23354 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 9398 26568 9404 26580
rect 9359 26540 9404 26568
rect 9398 26528 9404 26540
rect 9456 26528 9462 26580
rect 10042 26568 10048 26580
rect 10003 26540 10048 26568
rect 10042 26528 10048 26540
rect 10100 26528 10106 26580
rect 10686 26528 10692 26580
rect 10744 26568 10750 26580
rect 12618 26568 12624 26580
rect 10744 26540 12624 26568
rect 10744 26528 10750 26540
rect 12618 26528 12624 26540
rect 12676 26568 12682 26580
rect 13449 26571 13507 26577
rect 13449 26568 13461 26571
rect 12676 26540 13461 26568
rect 12676 26528 12682 26540
rect 13449 26537 13461 26540
rect 13495 26537 13507 26571
rect 13449 26531 13507 26537
rect 14645 26571 14703 26577
rect 14645 26537 14657 26571
rect 14691 26568 14703 26571
rect 15378 26568 15384 26580
rect 14691 26540 15384 26568
rect 14691 26537 14703 26540
rect 14645 26531 14703 26537
rect 15378 26528 15384 26540
rect 15436 26528 15442 26580
rect 20346 26528 20352 26580
rect 20404 26568 20410 26580
rect 21269 26571 21327 26577
rect 21269 26568 21281 26571
rect 20404 26540 21281 26568
rect 20404 26528 20410 26540
rect 21269 26537 21281 26540
rect 21315 26537 21327 26571
rect 33778 26568 33784 26580
rect 21269 26531 21327 26537
rect 22066 26540 33784 26568
rect 1857 26503 1915 26509
rect 1857 26469 1869 26503
rect 1903 26500 1915 26503
rect 22066 26500 22094 26540
rect 33778 26528 33784 26540
rect 33836 26528 33842 26580
rect 1903 26472 22094 26500
rect 1903 26469 1915 26472
rect 1857 26463 1915 26469
rect 34514 26460 34520 26512
rect 34572 26500 34578 26512
rect 38105 26503 38163 26509
rect 38105 26500 38117 26503
rect 34572 26472 38117 26500
rect 34572 26460 34578 26472
rect 38105 26469 38117 26472
rect 38151 26469 38163 26503
rect 38105 26463 38163 26469
rect 6730 26392 6736 26444
rect 6788 26432 6794 26444
rect 11977 26435 12035 26441
rect 11977 26432 11989 26435
rect 6788 26404 11989 26432
rect 6788 26392 6794 26404
rect 11977 26401 11989 26404
rect 12023 26401 12035 26435
rect 11977 26395 12035 26401
rect 12802 26392 12808 26444
rect 12860 26432 12866 26444
rect 13265 26435 13323 26441
rect 13265 26432 13277 26435
rect 12860 26404 13277 26432
rect 12860 26392 12866 26404
rect 13265 26401 13277 26404
rect 13311 26401 13323 26435
rect 15102 26432 15108 26444
rect 13265 26395 13323 26401
rect 14844 26404 15108 26432
rect 2498 26324 2504 26376
rect 2556 26364 2562 26376
rect 9309 26367 9367 26373
rect 9309 26364 9321 26367
rect 2556 26336 9321 26364
rect 2556 26324 2562 26336
rect 9309 26333 9321 26336
rect 9355 26333 9367 26367
rect 9309 26327 9367 26333
rect 10229 26367 10287 26373
rect 10229 26333 10241 26367
rect 10275 26364 10287 26367
rect 10502 26364 10508 26376
rect 10275 26336 10508 26364
rect 10275 26333 10287 26336
rect 10229 26327 10287 26333
rect 10502 26324 10508 26336
rect 10560 26324 10566 26376
rect 10686 26364 10692 26376
rect 10647 26336 10692 26364
rect 10686 26324 10692 26336
rect 10744 26324 10750 26376
rect 11517 26367 11575 26373
rect 11517 26333 11529 26367
rect 11563 26364 11575 26367
rect 11606 26364 11612 26376
rect 11563 26336 11612 26364
rect 11563 26333 11575 26336
rect 11517 26327 11575 26333
rect 11606 26324 11612 26336
rect 11664 26324 11670 26376
rect 12066 26324 12072 26376
rect 12124 26364 12130 26376
rect 12161 26367 12219 26373
rect 12161 26364 12173 26367
rect 12124 26336 12173 26364
rect 12124 26324 12130 26336
rect 12161 26333 12173 26336
rect 12207 26333 12219 26367
rect 12161 26327 12219 26333
rect 13081 26367 13139 26373
rect 13081 26333 13093 26367
rect 13127 26333 13139 26367
rect 13081 26327 13139 26333
rect 1670 26296 1676 26308
rect 1631 26268 1676 26296
rect 1670 26256 1676 26268
rect 1728 26256 1734 26308
rect 8202 26256 8208 26308
rect 8260 26296 8266 26308
rect 10781 26299 10839 26305
rect 10781 26296 10793 26299
rect 8260 26268 10793 26296
rect 8260 26256 8266 26268
rect 10781 26265 10793 26268
rect 10827 26265 10839 26299
rect 12986 26296 12992 26308
rect 10781 26259 10839 26265
rect 11348 26268 12992 26296
rect 11348 26237 11376 26268
rect 12986 26256 12992 26268
rect 13044 26256 13050 26308
rect 13096 26296 13124 26327
rect 14182 26324 14188 26376
rect 14240 26364 14246 26376
rect 14844 26373 14872 26404
rect 15102 26392 15108 26404
rect 15160 26432 15166 26444
rect 15473 26435 15531 26441
rect 15160 26404 15424 26432
rect 15160 26392 15166 26404
rect 14829 26367 14887 26373
rect 14829 26364 14841 26367
rect 14240 26336 14841 26364
rect 14240 26324 14246 26336
rect 14829 26333 14841 26336
rect 14875 26333 14887 26367
rect 14829 26327 14887 26333
rect 15289 26367 15347 26373
rect 15289 26333 15301 26367
rect 15335 26333 15347 26367
rect 15396 26364 15424 26404
rect 15473 26401 15485 26435
rect 15519 26432 15531 26435
rect 16485 26435 16543 26441
rect 16485 26432 16497 26435
rect 15519 26404 16497 26432
rect 15519 26401 15531 26404
rect 15473 26395 15531 26401
rect 16485 26401 16497 26404
rect 16531 26401 16543 26435
rect 16485 26395 16543 26401
rect 16393 26367 16451 26373
rect 16393 26364 16405 26367
rect 15396 26336 16405 26364
rect 15289 26327 15347 26333
rect 16393 26333 16405 26336
rect 16439 26333 16451 26367
rect 20806 26364 20812 26376
rect 20767 26336 20812 26364
rect 16393 26327 16451 26333
rect 15304 26296 15332 26327
rect 20806 26324 20812 26336
rect 20864 26324 20870 26376
rect 21453 26367 21511 26373
rect 21453 26333 21465 26367
rect 21499 26333 21511 26367
rect 21453 26327 21511 26333
rect 17954 26296 17960 26308
rect 13096 26268 15240 26296
rect 15304 26268 17960 26296
rect 11333 26231 11391 26237
rect 11333 26197 11345 26231
rect 11379 26197 11391 26231
rect 11333 26191 11391 26197
rect 12621 26231 12679 26237
rect 12621 26197 12633 26231
rect 12667 26228 12679 26231
rect 12894 26228 12900 26240
rect 12667 26200 12900 26228
rect 12667 26197 12679 26200
rect 12621 26191 12679 26197
rect 12894 26188 12900 26200
rect 12952 26228 12958 26240
rect 13446 26228 13452 26240
rect 12952 26200 13452 26228
rect 12952 26188 12958 26200
rect 13446 26188 13452 26200
rect 13504 26188 13510 26240
rect 15212 26228 15240 26268
rect 17954 26256 17960 26268
rect 18012 26296 18018 26308
rect 18230 26296 18236 26308
rect 18012 26268 18236 26296
rect 18012 26256 18018 26268
rect 18230 26256 18236 26268
rect 18288 26256 18294 26308
rect 21468 26296 21496 26327
rect 21910 26324 21916 26376
rect 21968 26364 21974 26376
rect 22649 26367 22707 26373
rect 22649 26364 22661 26367
rect 21968 26336 22661 26364
rect 21968 26324 21974 26336
rect 22649 26333 22661 26336
rect 22695 26333 22707 26367
rect 38286 26364 38292 26376
rect 38247 26336 38292 26364
rect 22649 26327 22707 26333
rect 38286 26324 38292 26336
rect 38344 26324 38350 26376
rect 20640 26268 21496 26296
rect 15286 26228 15292 26240
rect 15212 26200 15292 26228
rect 15286 26188 15292 26200
rect 15344 26228 15350 26240
rect 20640 26237 20668 26268
rect 15933 26231 15991 26237
rect 15933 26228 15945 26231
rect 15344 26200 15945 26228
rect 15344 26188 15350 26200
rect 15933 26197 15945 26200
rect 15979 26197 15991 26231
rect 15933 26191 15991 26197
rect 20625 26231 20683 26237
rect 20625 26197 20637 26231
rect 20671 26197 20683 26231
rect 22462 26228 22468 26240
rect 22423 26200 22468 26228
rect 20625 26191 20683 26197
rect 22462 26188 22468 26200
rect 22520 26188 22526 26240
rect 23106 26228 23112 26240
rect 23067 26200 23112 26228
rect 23106 26188 23112 26200
rect 23164 26188 23170 26240
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 13998 26024 14004 26036
rect 2746 25996 12434 26024
rect 13959 25996 14004 26024
rect 1762 25916 1768 25968
rect 1820 25956 1826 25968
rect 2746 25956 2774 25996
rect 1820 25928 2774 25956
rect 8389 25959 8447 25965
rect 1820 25916 1826 25928
rect 8389 25925 8401 25959
rect 8435 25956 8447 25959
rect 8478 25956 8484 25968
rect 8435 25928 8484 25956
rect 8435 25925 8447 25928
rect 8389 25919 8447 25925
rect 8478 25916 8484 25928
rect 8536 25916 8542 25968
rect 10778 25916 10784 25968
rect 10836 25956 10842 25968
rect 12069 25959 12127 25965
rect 12069 25956 12081 25959
rect 10836 25928 12081 25956
rect 10836 25916 10842 25928
rect 12069 25925 12081 25928
rect 12115 25925 12127 25959
rect 12406 25956 12434 25996
rect 13998 25984 14004 25996
rect 14056 25984 14062 26036
rect 15286 26024 15292 26036
rect 15247 25996 15292 26024
rect 15286 25984 15292 25996
rect 15344 25984 15350 26036
rect 20257 26027 20315 26033
rect 20257 26024 20269 26027
rect 16040 25996 20269 26024
rect 16040 25956 16068 25996
rect 20257 25993 20269 25996
rect 20303 25993 20315 26027
rect 20257 25987 20315 25993
rect 18414 25956 18420 25968
rect 12406 25928 16068 25956
rect 17236 25928 18420 25956
rect 12069 25919 12127 25925
rect 8297 25891 8355 25897
rect 8297 25857 8309 25891
rect 8343 25888 8355 25891
rect 9950 25888 9956 25900
rect 8343 25860 9956 25888
rect 8343 25857 8355 25860
rect 8297 25851 8355 25857
rect 9950 25848 9956 25860
rect 10008 25848 10014 25900
rect 10502 25888 10508 25900
rect 10463 25860 10508 25888
rect 10502 25848 10508 25860
rect 10560 25848 10566 25900
rect 13170 25848 13176 25900
rect 13228 25888 13234 25900
rect 14182 25888 14188 25900
rect 13228 25860 14188 25888
rect 13228 25848 13234 25860
rect 14182 25848 14188 25860
rect 14240 25848 14246 25900
rect 14645 25891 14703 25897
rect 14645 25857 14657 25891
rect 14691 25888 14703 25891
rect 14734 25888 14740 25900
rect 14691 25860 14740 25888
rect 14691 25857 14703 25860
rect 14645 25851 14703 25857
rect 14734 25848 14740 25860
rect 14792 25848 14798 25900
rect 14829 25891 14887 25897
rect 14829 25857 14841 25891
rect 14875 25888 14887 25891
rect 15194 25888 15200 25900
rect 14875 25860 15200 25888
rect 14875 25857 14887 25860
rect 14829 25851 14887 25857
rect 15194 25848 15200 25860
rect 15252 25848 15258 25900
rect 15746 25848 15752 25900
rect 15804 25888 15810 25900
rect 17236 25888 17264 25928
rect 18414 25916 18420 25928
rect 18472 25916 18478 25968
rect 18509 25959 18567 25965
rect 18509 25925 18521 25959
rect 18555 25956 18567 25959
rect 19518 25956 19524 25968
rect 18555 25928 19524 25956
rect 18555 25925 18567 25928
rect 18509 25919 18567 25925
rect 19518 25916 19524 25928
rect 19576 25916 19582 25968
rect 20165 25959 20223 25965
rect 20165 25925 20177 25959
rect 20211 25956 20223 25959
rect 24210 25956 24216 25968
rect 20211 25928 24216 25956
rect 20211 25925 20223 25928
rect 20165 25919 20223 25925
rect 24210 25916 24216 25928
rect 24268 25916 24274 25968
rect 15804 25860 17264 25888
rect 15804 25848 15810 25860
rect 19334 25848 19340 25900
rect 19392 25888 19398 25900
rect 20809 25891 20867 25897
rect 20809 25888 20821 25891
rect 19392 25860 20821 25888
rect 19392 25848 19398 25860
rect 20809 25857 20821 25860
rect 20855 25857 20867 25891
rect 20809 25851 20867 25857
rect 21818 25848 21824 25900
rect 21876 25888 21882 25900
rect 22005 25891 22063 25897
rect 22005 25888 22017 25891
rect 21876 25860 22017 25888
rect 21876 25848 21882 25860
rect 22005 25857 22017 25860
rect 22051 25857 22063 25891
rect 23106 25888 23112 25900
rect 23067 25860 23112 25888
rect 22005 25851 22063 25857
rect 23106 25848 23112 25860
rect 23164 25848 23170 25900
rect 23290 25888 23296 25900
rect 23251 25860 23296 25888
rect 23290 25848 23296 25860
rect 23348 25848 23354 25900
rect 30377 25891 30435 25897
rect 30377 25857 30389 25891
rect 30423 25888 30435 25891
rect 38102 25888 38108 25900
rect 30423 25860 38108 25888
rect 30423 25857 30435 25860
rect 30377 25851 30435 25857
rect 38102 25848 38108 25860
rect 38160 25848 38166 25900
rect 11790 25780 11796 25832
rect 11848 25820 11854 25832
rect 11977 25823 12035 25829
rect 11977 25820 11989 25823
rect 11848 25792 11989 25820
rect 11848 25780 11854 25792
rect 11977 25789 11989 25792
rect 12023 25789 12035 25823
rect 11977 25783 12035 25789
rect 12989 25823 13047 25829
rect 12989 25789 13001 25823
rect 13035 25820 13047 25823
rect 17954 25820 17960 25832
rect 13035 25792 17960 25820
rect 13035 25789 13047 25792
rect 12989 25783 13047 25789
rect 17954 25780 17960 25792
rect 18012 25780 18018 25832
rect 19242 25820 19248 25832
rect 19203 25792 19248 25820
rect 19242 25780 19248 25792
rect 19300 25780 19306 25832
rect 22186 25820 22192 25832
rect 22147 25792 22192 25820
rect 22186 25780 22192 25792
rect 22244 25780 22250 25832
rect 15194 25712 15200 25764
rect 15252 25752 15258 25764
rect 22922 25752 22928 25764
rect 15252 25724 22928 25752
rect 15252 25712 15258 25724
rect 22922 25712 22928 25724
rect 22980 25712 22986 25764
rect 10597 25687 10655 25693
rect 10597 25653 10609 25687
rect 10643 25684 10655 25687
rect 12158 25684 12164 25696
rect 10643 25656 12164 25684
rect 10643 25653 10655 25656
rect 10597 25647 10655 25653
rect 12158 25644 12164 25656
rect 12216 25644 12222 25696
rect 20901 25687 20959 25693
rect 20901 25653 20913 25687
rect 20947 25684 20959 25687
rect 21266 25684 21272 25696
rect 20947 25656 21272 25684
rect 20947 25653 20959 25656
rect 20901 25647 20959 25653
rect 21266 25644 21272 25656
rect 21324 25644 21330 25696
rect 22649 25687 22707 25693
rect 22649 25653 22661 25687
rect 22695 25684 22707 25687
rect 23753 25687 23811 25693
rect 23753 25684 23765 25687
rect 22695 25656 23765 25684
rect 22695 25653 22707 25656
rect 22649 25647 22707 25653
rect 23753 25653 23765 25656
rect 23799 25684 23811 25687
rect 24394 25684 24400 25696
rect 23799 25656 24400 25684
rect 23799 25653 23811 25656
rect 23753 25647 23811 25653
rect 24394 25644 24400 25656
rect 24452 25644 24458 25696
rect 24762 25644 24768 25696
rect 24820 25684 24826 25696
rect 30469 25687 30527 25693
rect 30469 25684 30481 25687
rect 24820 25656 30481 25684
rect 24820 25644 24826 25656
rect 30469 25653 30481 25656
rect 30515 25653 30527 25687
rect 30469 25647 30527 25653
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 10778 25480 10784 25492
rect 10739 25452 10784 25480
rect 10778 25440 10784 25452
rect 10836 25440 10842 25492
rect 12618 25480 12624 25492
rect 12579 25452 12624 25480
rect 12618 25440 12624 25452
rect 12676 25440 12682 25492
rect 13446 25480 13452 25492
rect 13407 25452 13452 25480
rect 13446 25440 13452 25452
rect 13504 25440 13510 25492
rect 16390 25480 16396 25492
rect 15028 25452 16396 25480
rect 6365 25415 6423 25421
rect 6365 25381 6377 25415
rect 6411 25412 6423 25415
rect 11790 25412 11796 25424
rect 6411 25384 11796 25412
rect 6411 25381 6423 25384
rect 6365 25375 6423 25381
rect 11790 25372 11796 25384
rect 11848 25372 11854 25424
rect 14642 25412 14648 25424
rect 12406 25384 14648 25412
rect 11977 25347 12035 25353
rect 11977 25313 11989 25347
rect 12023 25344 12035 25347
rect 12406 25344 12434 25384
rect 14642 25372 14648 25384
rect 14700 25372 14706 25424
rect 13262 25344 13268 25356
rect 12023 25316 12434 25344
rect 13223 25316 13268 25344
rect 12023 25313 12035 25316
rect 11977 25307 12035 25313
rect 13262 25304 13268 25316
rect 13320 25304 13326 25356
rect 1946 25236 1952 25288
rect 2004 25276 2010 25288
rect 2130 25276 2136 25288
rect 2004 25248 2136 25276
rect 2004 25236 2010 25248
rect 2130 25236 2136 25248
rect 2188 25276 2194 25288
rect 6273 25279 6331 25285
rect 6273 25276 6285 25279
rect 2188 25248 6285 25276
rect 2188 25236 2194 25248
rect 6273 25245 6285 25248
rect 6319 25245 6331 25279
rect 10686 25276 10692 25288
rect 10647 25248 10692 25276
rect 6273 25239 6331 25245
rect 10686 25236 10692 25248
rect 10744 25236 10750 25288
rect 12158 25276 12164 25288
rect 12119 25248 12164 25276
rect 12158 25236 12164 25248
rect 12216 25236 12222 25288
rect 13081 25279 13139 25285
rect 13081 25276 13093 25279
rect 12406 25248 13093 25276
rect 11333 25211 11391 25217
rect 11333 25177 11345 25211
rect 11379 25208 11391 25211
rect 12406 25208 12434 25248
rect 13081 25245 13093 25248
rect 13127 25245 13139 25279
rect 13081 25239 13139 25245
rect 14277 25279 14335 25285
rect 14277 25245 14289 25279
rect 14323 25276 14335 25279
rect 15028 25276 15056 25452
rect 16390 25440 16396 25452
rect 16448 25440 16454 25492
rect 19518 25480 19524 25492
rect 19479 25452 19524 25480
rect 19518 25440 19524 25452
rect 19576 25440 19582 25492
rect 24670 25480 24676 25492
rect 24631 25452 24676 25480
rect 24670 25440 24676 25452
rect 24728 25440 24734 25492
rect 15102 25372 15108 25424
rect 15160 25372 15166 25424
rect 17954 25372 17960 25424
rect 18012 25412 18018 25424
rect 18012 25384 21496 25412
rect 18012 25372 18018 25384
rect 15120 25344 15148 25372
rect 21468 25356 21496 25384
rect 21174 25344 21180 25356
rect 15120 25316 15700 25344
rect 21135 25316 21180 25344
rect 14323 25248 15056 25276
rect 15105 25279 15163 25285
rect 14323 25245 14335 25248
rect 14277 25239 14335 25245
rect 15105 25245 15117 25279
rect 15151 25276 15163 25279
rect 15194 25276 15200 25288
rect 15151 25248 15200 25276
rect 15151 25245 15163 25248
rect 15105 25239 15163 25245
rect 15194 25236 15200 25248
rect 15252 25236 15258 25288
rect 15672 25278 15700 25316
rect 21174 25304 21180 25316
rect 21232 25304 21238 25356
rect 21450 25344 21456 25356
rect 21363 25316 21456 25344
rect 21450 25304 21456 25316
rect 21508 25304 21514 25356
rect 15749 25279 15807 25285
rect 15749 25278 15761 25279
rect 15672 25250 15761 25278
rect 15749 25245 15761 25250
rect 15795 25245 15807 25279
rect 15749 25239 15807 25245
rect 16390 25236 16396 25288
rect 16448 25276 16454 25288
rect 16669 25279 16727 25285
rect 16669 25276 16681 25279
rect 16448 25248 16681 25276
rect 16448 25236 16454 25248
rect 16669 25245 16681 25248
rect 16715 25245 16727 25279
rect 16669 25239 16727 25245
rect 19334 25236 19340 25288
rect 19392 25276 19398 25288
rect 19429 25279 19487 25285
rect 19429 25276 19441 25279
rect 19392 25248 19441 25276
rect 19392 25236 19398 25248
rect 19429 25245 19441 25248
rect 19475 25245 19487 25279
rect 19429 25239 19487 25245
rect 22462 25236 22468 25288
rect 22520 25276 22526 25288
rect 23109 25279 23167 25285
rect 23109 25276 23121 25279
rect 22520 25248 23121 25276
rect 22520 25236 22526 25248
rect 23109 25245 23121 25248
rect 23155 25245 23167 25279
rect 23109 25239 23167 25245
rect 24581 25279 24639 25285
rect 24581 25245 24593 25279
rect 24627 25276 24639 25279
rect 27430 25276 27436 25288
rect 24627 25248 27436 25276
rect 24627 25245 24639 25248
rect 24581 25239 24639 25245
rect 27430 25236 27436 25248
rect 27488 25236 27494 25288
rect 31113 25279 31171 25285
rect 31113 25245 31125 25279
rect 31159 25276 31171 25279
rect 34514 25276 34520 25288
rect 31159 25248 34520 25276
rect 31159 25245 31171 25248
rect 31113 25239 31171 25245
rect 34514 25236 34520 25248
rect 34572 25236 34578 25288
rect 38010 25276 38016 25288
rect 37971 25248 38016 25276
rect 38010 25236 38016 25248
rect 38068 25236 38074 25288
rect 11379 25180 12434 25208
rect 11379 25177 11391 25180
rect 11333 25171 11391 25177
rect 14734 25168 14740 25220
rect 14792 25208 14798 25220
rect 15841 25211 15899 25217
rect 15841 25208 15853 25211
rect 14792 25180 15853 25208
rect 14792 25168 14798 25180
rect 15841 25177 15853 25180
rect 15887 25177 15899 25211
rect 15841 25171 15899 25177
rect 21266 25168 21272 25220
rect 21324 25208 21330 25220
rect 21324 25180 21369 25208
rect 21324 25168 21330 25180
rect 14366 25140 14372 25152
rect 14327 25112 14372 25140
rect 14366 25100 14372 25112
rect 14424 25100 14430 25152
rect 15194 25140 15200 25152
rect 15155 25112 15200 25140
rect 15194 25100 15200 25112
rect 15252 25100 15258 25152
rect 16761 25143 16819 25149
rect 16761 25109 16773 25143
rect 16807 25140 16819 25143
rect 17218 25140 17224 25152
rect 16807 25112 17224 25140
rect 16807 25109 16819 25112
rect 16761 25103 16819 25109
rect 17218 25100 17224 25112
rect 17276 25100 17282 25152
rect 22925 25143 22983 25149
rect 22925 25109 22937 25143
rect 22971 25140 22983 25143
rect 24762 25140 24768 25152
rect 22971 25112 24768 25140
rect 22971 25109 22983 25112
rect 22925 25103 22983 25109
rect 24762 25100 24768 25112
rect 24820 25100 24826 25152
rect 31202 25140 31208 25152
rect 31163 25112 31208 25140
rect 31202 25100 31208 25112
rect 31260 25100 31266 25152
rect 38194 25140 38200 25152
rect 38155 25112 38200 25140
rect 38194 25100 38200 25112
rect 38252 25100 38258 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 19242 24936 19248 24948
rect 14660 24908 19248 24936
rect 13173 24871 13231 24877
rect 13173 24837 13185 24871
rect 13219 24868 13231 24871
rect 14366 24868 14372 24880
rect 13219 24840 14372 24868
rect 13219 24837 13231 24840
rect 13173 24831 13231 24837
rect 14366 24828 14372 24840
rect 14424 24828 14430 24880
rect 14660 24868 14688 24908
rect 19242 24896 19248 24908
rect 19300 24896 19306 24948
rect 22097 24939 22155 24945
rect 22097 24905 22109 24939
rect 22143 24936 22155 24939
rect 22186 24936 22192 24948
rect 22143 24908 22192 24936
rect 22143 24905 22155 24908
rect 22097 24899 22155 24905
rect 22186 24896 22192 24908
rect 22244 24896 22250 24948
rect 24213 24939 24271 24945
rect 24213 24905 24225 24939
rect 24259 24905 24271 24939
rect 24213 24899 24271 24905
rect 14476 24840 14688 24868
rect 14737 24871 14795 24877
rect 1581 24803 1639 24809
rect 1581 24769 1593 24803
rect 1627 24800 1639 24803
rect 4062 24800 4068 24812
rect 1627 24772 4068 24800
rect 1627 24769 1639 24772
rect 1581 24763 1639 24769
rect 4062 24760 4068 24772
rect 4120 24760 4126 24812
rect 8662 24760 8668 24812
rect 8720 24800 8726 24812
rect 10597 24803 10655 24809
rect 10597 24800 10609 24803
rect 8720 24772 10609 24800
rect 8720 24760 8726 24772
rect 10597 24769 10609 24772
rect 10643 24800 10655 24803
rect 10686 24800 10692 24812
rect 10643 24772 10692 24800
rect 10643 24769 10655 24772
rect 10597 24763 10655 24769
rect 10686 24760 10692 24772
rect 10744 24760 10750 24812
rect 11606 24760 11612 24812
rect 11664 24800 11670 24812
rect 11701 24803 11759 24809
rect 11701 24800 11713 24803
rect 11664 24772 11713 24800
rect 11664 24760 11670 24772
rect 11701 24769 11713 24772
rect 11747 24769 11759 24803
rect 11701 24763 11759 24769
rect 11793 24803 11851 24809
rect 11793 24769 11805 24803
rect 11839 24800 11851 24803
rect 12066 24800 12072 24812
rect 11839 24772 12072 24800
rect 11839 24769 11851 24772
rect 11793 24763 11851 24769
rect 11716 24732 11744 24763
rect 12066 24760 12072 24772
rect 12124 24760 12130 24812
rect 12345 24803 12403 24809
rect 12345 24769 12357 24803
rect 12391 24800 12403 24803
rect 12894 24800 12900 24812
rect 12391 24772 12900 24800
rect 12391 24769 12403 24772
rect 12345 24763 12403 24769
rect 12894 24760 12900 24772
rect 12952 24760 12958 24812
rect 12710 24732 12716 24744
rect 11716 24704 12716 24732
rect 12710 24692 12716 24704
rect 12768 24692 12774 24744
rect 13078 24732 13084 24744
rect 13039 24704 13084 24732
rect 13078 24692 13084 24704
rect 13136 24692 13142 24744
rect 13354 24692 13360 24744
rect 13412 24732 13418 24744
rect 14093 24735 14151 24741
rect 14093 24732 14105 24735
rect 13412 24704 14105 24732
rect 13412 24692 13418 24704
rect 14093 24701 14105 24704
rect 14139 24732 14151 24735
rect 14476 24732 14504 24840
rect 14737 24837 14749 24871
rect 14783 24868 14795 24871
rect 18049 24871 18107 24877
rect 18049 24868 18061 24871
rect 14783 24840 15516 24868
rect 14783 24837 14795 24840
rect 14737 24831 14795 24837
rect 15488 24800 15516 24840
rect 17788 24840 18061 24868
rect 16117 24803 16175 24809
rect 15488 24772 15792 24800
rect 14139 24704 14504 24732
rect 14645 24735 14703 24741
rect 14139 24701 14151 24704
rect 14093 24695 14151 24701
rect 14645 24701 14657 24735
rect 14691 24732 14703 24735
rect 15194 24732 15200 24744
rect 14691 24704 15200 24732
rect 14691 24701 14703 24704
rect 14645 24695 14703 24701
rect 15194 24692 15200 24704
rect 15252 24692 15258 24744
rect 15289 24735 15347 24741
rect 15289 24701 15301 24735
rect 15335 24701 15347 24735
rect 15764 24732 15792 24772
rect 16117 24769 16129 24803
rect 16163 24800 16175 24803
rect 16298 24800 16304 24812
rect 16163 24772 16304 24800
rect 16163 24769 16175 24772
rect 16117 24763 16175 24769
rect 16298 24760 16304 24772
rect 16356 24800 16362 24812
rect 17221 24803 17279 24809
rect 17221 24800 17233 24803
rect 16356 24772 17233 24800
rect 16356 24760 16362 24772
rect 17221 24769 17233 24772
rect 17267 24769 17279 24803
rect 17221 24763 17279 24769
rect 17313 24803 17371 24809
rect 17313 24769 17325 24803
rect 17359 24800 17371 24803
rect 17788 24800 17816 24840
rect 18049 24837 18061 24840
rect 18095 24837 18107 24871
rect 22922 24868 22928 24880
rect 22883 24840 22928 24868
rect 18049 24831 18107 24837
rect 22922 24828 22928 24840
rect 22980 24828 22986 24880
rect 24228 24868 24256 24899
rect 24228 24840 24532 24868
rect 17359 24772 17816 24800
rect 19613 24803 19671 24809
rect 17359 24769 17371 24772
rect 17313 24763 17371 24769
rect 19613 24769 19625 24803
rect 19659 24800 19671 24803
rect 19978 24800 19984 24812
rect 19659 24772 19984 24800
rect 19659 24769 19671 24772
rect 19613 24763 19671 24769
rect 19978 24760 19984 24772
rect 20036 24760 20042 24812
rect 21910 24760 21916 24812
rect 21968 24800 21974 24812
rect 22005 24803 22063 24809
rect 22005 24800 22017 24803
rect 21968 24772 22017 24800
rect 21968 24760 21974 24772
rect 22005 24769 22017 24772
rect 22051 24769 22063 24803
rect 22005 24763 22063 24769
rect 24302 24760 24308 24812
rect 24360 24800 24366 24812
rect 24397 24803 24455 24809
rect 24397 24800 24409 24803
rect 24360 24772 24409 24800
rect 24360 24760 24366 24772
rect 24397 24769 24409 24772
rect 24443 24769 24455 24803
rect 24504 24800 24532 24840
rect 25041 24803 25099 24809
rect 25041 24800 25053 24803
rect 24504 24772 25053 24800
rect 24397 24763 24455 24769
rect 25041 24769 25053 24772
rect 25087 24769 25099 24803
rect 25774 24800 25780 24812
rect 25735 24772 25780 24800
rect 25041 24763 25099 24769
rect 25774 24760 25780 24772
rect 25832 24760 25838 24812
rect 25869 24803 25927 24809
rect 25869 24769 25881 24803
rect 25915 24800 25927 24803
rect 26878 24800 26884 24812
rect 25915 24772 26884 24800
rect 25915 24769 25927 24772
rect 25869 24763 25927 24769
rect 26878 24760 26884 24772
rect 26936 24760 26942 24812
rect 30653 24803 30711 24809
rect 30653 24769 30665 24803
rect 30699 24800 30711 24803
rect 37642 24800 37648 24812
rect 30699 24772 37648 24800
rect 30699 24769 30711 24772
rect 30653 24763 30711 24769
rect 37642 24760 37648 24772
rect 37700 24760 37706 24812
rect 16209 24735 16267 24741
rect 16209 24732 16221 24735
rect 15764 24704 16221 24732
rect 15289 24695 15347 24701
rect 16209 24701 16221 24704
rect 16255 24701 16267 24735
rect 16209 24695 16267 24701
rect 17957 24723 18015 24729
rect 15102 24624 15108 24676
rect 15160 24664 15166 24676
rect 15304 24664 15332 24695
rect 17957 24689 17969 24723
rect 18003 24689 18015 24723
rect 18046 24692 18052 24744
rect 18104 24732 18110 24744
rect 18233 24735 18291 24741
rect 18233 24732 18245 24735
rect 18104 24704 18245 24732
rect 18104 24692 18110 24704
rect 18233 24701 18245 24704
rect 18279 24701 18291 24735
rect 18233 24695 18291 24701
rect 20714 24692 20720 24744
rect 20772 24732 20778 24744
rect 22833 24735 22891 24741
rect 22833 24732 22845 24735
rect 20772 24704 22845 24732
rect 20772 24692 20778 24704
rect 22833 24701 22845 24704
rect 22879 24701 22891 24735
rect 31202 24732 31208 24744
rect 22833 24695 22891 24701
rect 22940 24704 31208 24732
rect 17957 24683 18015 24689
rect 15160 24636 15332 24664
rect 15160 24624 15166 24636
rect 1762 24596 1768 24608
rect 1723 24568 1768 24596
rect 1762 24556 1768 24568
rect 1820 24556 1826 24608
rect 10318 24556 10324 24608
rect 10376 24596 10382 24608
rect 10689 24599 10747 24605
rect 10689 24596 10701 24599
rect 10376 24568 10701 24596
rect 10376 24556 10382 24568
rect 10689 24565 10701 24568
rect 10735 24565 10747 24599
rect 10689 24559 10747 24565
rect 12437 24599 12495 24605
rect 12437 24565 12449 24599
rect 12483 24596 12495 24599
rect 12618 24596 12624 24608
rect 12483 24568 12624 24596
rect 12483 24565 12495 24568
rect 12437 24559 12495 24565
rect 12618 24556 12624 24568
rect 12676 24556 12682 24608
rect 17972 24596 18000 24683
rect 22940 24664 22968 24704
rect 31202 24692 31208 24704
rect 31260 24692 31266 24744
rect 19352 24636 22968 24664
rect 23385 24667 23443 24673
rect 19352 24596 19380 24636
rect 23385 24633 23397 24667
rect 23431 24664 23443 24667
rect 27154 24664 27160 24676
rect 23431 24636 27160 24664
rect 23431 24633 23443 24636
rect 23385 24627 23443 24633
rect 27154 24624 27160 24636
rect 27212 24664 27218 24676
rect 27522 24664 27528 24676
rect 27212 24636 27528 24664
rect 27212 24624 27218 24636
rect 27522 24624 27528 24636
rect 27580 24624 27586 24676
rect 17972 24568 19380 24596
rect 19429 24599 19487 24605
rect 19429 24565 19441 24599
rect 19475 24596 19487 24599
rect 22830 24596 22836 24608
rect 19475 24568 22836 24596
rect 19475 24565 19487 24568
rect 19429 24559 19487 24565
rect 22830 24556 22836 24568
rect 22888 24556 22894 24608
rect 22922 24556 22928 24608
rect 22980 24596 22986 24608
rect 24857 24599 24915 24605
rect 24857 24596 24869 24599
rect 22980 24568 24869 24596
rect 22980 24556 22986 24568
rect 24857 24565 24869 24568
rect 24903 24565 24915 24599
rect 24857 24559 24915 24565
rect 30650 24556 30656 24608
rect 30708 24596 30714 24608
rect 30745 24599 30803 24605
rect 30745 24596 30757 24599
rect 30708 24568 30757 24596
rect 30708 24556 30714 24568
rect 30745 24565 30757 24568
rect 30791 24565 30803 24599
rect 30745 24559 30803 24565
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 14642 24352 14648 24404
rect 14700 24392 14706 24404
rect 14737 24395 14795 24401
rect 14737 24392 14749 24395
rect 14700 24364 14749 24392
rect 14700 24352 14706 24364
rect 14737 24361 14749 24364
rect 14783 24361 14795 24395
rect 14737 24355 14795 24361
rect 23106 24352 23112 24404
rect 23164 24392 23170 24404
rect 25774 24392 25780 24404
rect 23164 24364 25780 24392
rect 23164 24352 23170 24364
rect 25774 24352 25780 24364
rect 25832 24352 25838 24404
rect 11882 24284 11888 24336
rect 11940 24324 11946 24336
rect 16850 24324 16856 24336
rect 11940 24296 16856 24324
rect 11940 24284 11946 24296
rect 16850 24284 16856 24296
rect 16908 24284 16914 24336
rect 17678 24324 17684 24336
rect 17639 24296 17684 24324
rect 17678 24284 17684 24296
rect 17736 24284 17742 24336
rect 23290 24284 23296 24336
rect 23348 24324 23354 24336
rect 23348 24296 24624 24324
rect 23348 24284 23354 24296
rect 24596 24268 24624 24296
rect 24854 24284 24860 24336
rect 24912 24324 24918 24336
rect 24949 24327 25007 24333
rect 24949 24324 24961 24327
rect 24912 24296 24961 24324
rect 24912 24284 24918 24296
rect 24949 24293 24961 24296
rect 24995 24293 25007 24327
rect 24949 24287 25007 24293
rect 12526 24256 12532 24268
rect 12487 24228 12532 24256
rect 12526 24216 12532 24228
rect 12584 24216 12590 24268
rect 12894 24216 12900 24268
rect 12952 24256 12958 24268
rect 13262 24256 13268 24268
rect 12952 24228 13268 24256
rect 12952 24216 12958 24228
rect 13262 24216 13268 24228
rect 13320 24256 13326 24268
rect 14550 24256 14556 24268
rect 13320 24228 13860 24256
rect 14511 24228 14556 24256
rect 13320 24216 13326 24228
rect 1578 24188 1584 24200
rect 1539 24160 1584 24188
rect 1578 24148 1584 24160
rect 1636 24148 1642 24200
rect 1854 24188 1860 24200
rect 1815 24160 1860 24188
rect 1854 24148 1860 24160
rect 1912 24148 1918 24200
rect 12618 24080 12624 24132
rect 12676 24120 12682 24132
rect 13173 24123 13231 24129
rect 12676 24092 12721 24120
rect 12676 24080 12682 24092
rect 13173 24089 13185 24123
rect 13219 24120 13231 24123
rect 13722 24120 13728 24132
rect 13219 24092 13728 24120
rect 13219 24089 13231 24092
rect 13173 24083 13231 24089
rect 13722 24080 13728 24092
rect 13780 24080 13786 24132
rect 13832 24120 13860 24228
rect 14550 24216 14556 24228
rect 14608 24216 14614 24268
rect 22094 24216 22100 24268
rect 22152 24256 22158 24268
rect 22741 24259 22799 24265
rect 22741 24256 22753 24259
rect 22152 24228 22753 24256
rect 22152 24216 22158 24228
rect 22741 24225 22753 24228
rect 22787 24256 22799 24259
rect 24578 24256 24584 24268
rect 22787 24228 23888 24256
rect 24491 24228 24584 24256
rect 22787 24225 22799 24228
rect 22741 24219 22799 24225
rect 14369 24191 14427 24197
rect 14369 24157 14381 24191
rect 14415 24188 14427 24191
rect 15194 24188 15200 24200
rect 14415 24160 15200 24188
rect 14415 24157 14427 24160
rect 14369 24151 14427 24157
rect 15194 24148 15200 24160
rect 15252 24148 15258 24200
rect 15286 24148 15292 24200
rect 15344 24188 15350 24200
rect 15565 24191 15623 24197
rect 15565 24188 15577 24191
rect 15344 24160 15577 24188
rect 15344 24148 15350 24160
rect 15565 24157 15577 24160
rect 15611 24157 15623 24191
rect 16761 24191 16819 24197
rect 16761 24188 16773 24191
rect 15565 24151 15623 24157
rect 15672 24160 16773 24188
rect 15672 24120 15700 24160
rect 16761 24157 16773 24160
rect 16807 24157 16819 24191
rect 16761 24151 16819 24157
rect 16853 24191 16911 24197
rect 16853 24157 16865 24191
rect 16899 24188 16911 24191
rect 16899 24160 18276 24188
rect 16899 24157 16911 24160
rect 16853 24151 16911 24157
rect 13832 24092 15700 24120
rect 15838 24080 15844 24132
rect 15896 24120 15902 24132
rect 17497 24123 17555 24129
rect 17497 24120 17509 24123
rect 15896 24092 17509 24120
rect 15896 24080 15902 24092
rect 17497 24089 17509 24092
rect 17543 24089 17555 24123
rect 18248 24120 18276 24160
rect 18322 24148 18328 24200
rect 18380 24188 18386 24200
rect 18380 24160 18425 24188
rect 18380 24148 18386 24160
rect 22833 24123 22891 24129
rect 18248 24092 22692 24120
rect 17497 24083 17555 24089
rect 15654 24052 15660 24064
rect 15615 24024 15660 24052
rect 15654 24012 15660 24024
rect 15712 24012 15718 24064
rect 18417 24055 18475 24061
rect 18417 24021 18429 24055
rect 18463 24052 18475 24055
rect 18782 24052 18788 24064
rect 18463 24024 18788 24052
rect 18463 24021 18475 24024
rect 18417 24015 18475 24021
rect 18782 24012 18788 24024
rect 18840 24012 18846 24064
rect 20070 24052 20076 24064
rect 20031 24024 20076 24052
rect 20070 24012 20076 24024
rect 20128 24012 20134 24064
rect 22664 24052 22692 24092
rect 22833 24089 22845 24123
rect 22879 24089 22891 24123
rect 23753 24123 23811 24129
rect 23753 24120 23765 24123
rect 22833 24083 22891 24089
rect 23492 24092 23765 24120
rect 22848 24052 22876 24083
rect 23492 24064 23520 24092
rect 23753 24089 23765 24092
rect 23799 24089 23811 24123
rect 23860 24120 23888 24228
rect 24578 24216 24584 24228
rect 24636 24216 24642 24268
rect 24762 24256 24768 24268
rect 24723 24228 24768 24256
rect 24762 24216 24768 24228
rect 24820 24216 24826 24268
rect 37734 24256 37740 24268
rect 35866 24228 37740 24256
rect 29733 24191 29791 24197
rect 29733 24157 29745 24191
rect 29779 24188 29791 24191
rect 35866 24188 35894 24228
rect 37734 24216 37740 24228
rect 37792 24216 37798 24268
rect 37458 24188 37464 24200
rect 29779 24160 35894 24188
rect 37419 24160 37464 24188
rect 29779 24157 29791 24160
rect 29733 24151 29791 24157
rect 37458 24148 37464 24160
rect 37516 24148 37522 24200
rect 30466 24120 30472 24132
rect 23860 24092 30472 24120
rect 23753 24083 23811 24089
rect 30466 24080 30472 24092
rect 30524 24080 30530 24132
rect 22664 24024 22876 24052
rect 23474 24012 23480 24064
rect 23532 24012 23538 24064
rect 24302 24012 24308 24064
rect 24360 24052 24366 24064
rect 24762 24052 24768 24064
rect 24360 24024 24768 24052
rect 24360 24012 24366 24024
rect 24762 24012 24768 24024
rect 24820 24012 24826 24064
rect 27982 24012 27988 24064
rect 28040 24052 28046 24064
rect 29825 24055 29883 24061
rect 29825 24052 29837 24055
rect 28040 24024 29837 24052
rect 28040 24012 28046 24024
rect 29825 24021 29837 24024
rect 29871 24021 29883 24055
rect 29825 24015 29883 24021
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 1854 23808 1860 23860
rect 1912 23848 1918 23860
rect 15838 23848 15844 23860
rect 1912 23820 15844 23848
rect 1912 23808 1918 23820
rect 15838 23808 15844 23820
rect 15896 23808 15902 23860
rect 19245 23851 19303 23857
rect 19245 23817 19257 23851
rect 19291 23848 19303 23851
rect 20714 23848 20720 23860
rect 19291 23820 20720 23848
rect 19291 23817 19303 23820
rect 19245 23811 19303 23817
rect 20714 23808 20720 23820
rect 20772 23808 20778 23860
rect 22830 23808 22836 23860
rect 22888 23848 22894 23860
rect 30466 23848 30472 23860
rect 22888 23820 26234 23848
rect 30427 23820 30472 23848
rect 22888 23808 22894 23820
rect 12986 23780 12992 23792
rect 12947 23752 12992 23780
rect 12986 23740 12992 23752
rect 13044 23740 13050 23792
rect 15381 23783 15439 23789
rect 15381 23749 15393 23783
rect 15427 23780 15439 23783
rect 16945 23783 17003 23789
rect 16945 23780 16957 23783
rect 15427 23752 16957 23780
rect 15427 23749 15439 23752
rect 15381 23743 15439 23749
rect 16945 23749 16957 23752
rect 16991 23749 17003 23783
rect 21634 23780 21640 23792
rect 16945 23743 17003 23749
rect 17788 23752 21640 23780
rect 2130 23712 2136 23724
rect 2091 23684 2136 23712
rect 2130 23672 2136 23684
rect 2188 23672 2194 23724
rect 4709 23715 4767 23721
rect 4709 23681 4721 23715
rect 4755 23712 4767 23715
rect 7006 23712 7012 23724
rect 4755 23684 7012 23712
rect 4755 23681 4767 23684
rect 4709 23675 4767 23681
rect 7006 23672 7012 23684
rect 7064 23672 7070 23724
rect 10042 23672 10048 23724
rect 10100 23712 10106 23724
rect 10137 23715 10195 23721
rect 10137 23712 10149 23715
rect 10100 23684 10149 23712
rect 10100 23672 10106 23684
rect 10137 23681 10149 23684
rect 10183 23681 10195 23715
rect 10137 23675 10195 23681
rect 10410 23672 10416 23724
rect 10468 23712 10474 23724
rect 11885 23715 11943 23721
rect 11885 23712 11897 23715
rect 10468 23684 11897 23712
rect 10468 23672 10474 23684
rect 11885 23681 11897 23684
rect 11931 23712 11943 23715
rect 14553 23715 14611 23721
rect 11931 23684 12434 23712
rect 11931 23681 11943 23684
rect 11885 23675 11943 23681
rect 4062 23536 4068 23588
rect 4120 23576 4126 23588
rect 4525 23579 4583 23585
rect 4525 23576 4537 23579
rect 4120 23548 4537 23576
rect 4120 23536 4126 23548
rect 4525 23545 4537 23548
rect 4571 23545 4583 23579
rect 12406 23576 12434 23684
rect 14553 23681 14565 23715
rect 14599 23712 14611 23715
rect 14918 23712 14924 23724
rect 14599 23684 14924 23712
rect 14599 23681 14611 23684
rect 14553 23675 14611 23681
rect 12897 23647 12955 23653
rect 12897 23613 12909 23647
rect 12943 23644 12955 23647
rect 13078 23644 13084 23656
rect 12943 23616 13084 23644
rect 12943 23613 12955 23616
rect 12897 23607 12955 23613
rect 13078 23604 13084 23616
rect 13136 23604 13142 23656
rect 14568 23644 14596 23675
rect 14918 23672 14924 23684
rect 14976 23672 14982 23724
rect 16850 23712 16856 23724
rect 16811 23684 16856 23712
rect 16850 23672 16856 23684
rect 16908 23672 16914 23724
rect 17788 23721 17816 23752
rect 21634 23740 21640 23752
rect 21692 23780 21698 23792
rect 21910 23780 21916 23792
rect 21692 23752 21916 23780
rect 21692 23740 21698 23752
rect 21910 23740 21916 23752
rect 21968 23740 21974 23792
rect 22186 23780 22192 23792
rect 22147 23752 22192 23780
rect 22186 23740 22192 23752
rect 22244 23740 22250 23792
rect 23382 23780 23388 23792
rect 23343 23752 23388 23780
rect 23382 23740 23388 23752
rect 23440 23740 23446 23792
rect 26206 23780 26234 23820
rect 30466 23808 30472 23820
rect 30524 23808 30530 23860
rect 38010 23780 38016 23792
rect 26206 23752 38016 23780
rect 38010 23740 38016 23752
rect 38068 23740 38074 23792
rect 17773 23715 17831 23721
rect 17773 23681 17785 23715
rect 17819 23681 17831 23715
rect 18598 23712 18604 23724
rect 18559 23684 18604 23712
rect 17773 23675 17831 23681
rect 18598 23672 18604 23684
rect 18656 23672 18662 23724
rect 18782 23712 18788 23724
rect 18743 23684 18788 23712
rect 18782 23672 18788 23684
rect 18840 23672 18846 23724
rect 20070 23712 20076 23724
rect 20031 23684 20076 23712
rect 20070 23672 20076 23684
rect 20128 23672 20134 23724
rect 20257 23715 20315 23721
rect 20257 23681 20269 23715
rect 20303 23712 20315 23715
rect 20346 23712 20352 23724
rect 20303 23684 20352 23712
rect 20303 23681 20315 23684
rect 20257 23675 20315 23681
rect 20346 23672 20352 23684
rect 20404 23672 20410 23724
rect 24578 23672 24584 23724
rect 24636 23712 24642 23724
rect 27982 23712 27988 23724
rect 24636 23684 27988 23712
rect 24636 23672 24642 23684
rect 27982 23672 27988 23684
rect 28040 23672 28046 23724
rect 29733 23715 29791 23721
rect 29733 23681 29745 23715
rect 29779 23681 29791 23715
rect 29733 23675 29791 23681
rect 30377 23715 30435 23721
rect 30377 23681 30389 23715
rect 30423 23712 30435 23715
rect 34606 23712 34612 23724
rect 30423 23684 34612 23712
rect 30423 23681 30435 23684
rect 30377 23675 30435 23681
rect 15286 23644 15292 23656
rect 13372 23616 14596 23644
rect 15247 23616 15292 23644
rect 13372 23576 13400 23616
rect 15286 23604 15292 23616
rect 15344 23604 15350 23656
rect 15565 23647 15623 23653
rect 15565 23613 15577 23647
rect 15611 23613 15623 23647
rect 22094 23644 22100 23656
rect 22055 23616 22100 23644
rect 15565 23607 15623 23613
rect 12406 23548 13400 23576
rect 4525 23539 4583 23545
rect 13446 23536 13452 23588
rect 13504 23576 13510 23588
rect 13504 23548 13549 23576
rect 13504 23536 13510 23548
rect 14182 23536 14188 23588
rect 14240 23576 14246 23588
rect 15102 23576 15108 23588
rect 14240 23548 15108 23576
rect 14240 23536 14246 23548
rect 15102 23536 15108 23548
rect 15160 23576 15166 23588
rect 15580 23576 15608 23607
rect 22094 23604 22100 23616
rect 22152 23604 22158 23656
rect 22370 23644 22376 23656
rect 22331 23616 22376 23644
rect 22370 23604 22376 23616
rect 22428 23604 22434 23656
rect 23293 23647 23351 23653
rect 23293 23613 23305 23647
rect 23339 23613 23351 23647
rect 23293 23607 23351 23613
rect 15160 23548 15608 23576
rect 23308 23576 23336 23607
rect 23474 23604 23480 23656
rect 23532 23644 23538 23656
rect 23569 23647 23627 23653
rect 23569 23644 23581 23647
rect 23532 23616 23581 23644
rect 23532 23604 23538 23616
rect 23569 23613 23581 23616
rect 23615 23613 23627 23647
rect 29748 23644 29776 23675
rect 34606 23672 34612 23684
rect 34664 23672 34670 23724
rect 37918 23644 37924 23656
rect 29748 23616 37924 23644
rect 23569 23607 23627 23613
rect 37918 23604 37924 23616
rect 37976 23604 37982 23656
rect 24670 23576 24676 23588
rect 23308 23548 24676 23576
rect 15160 23536 15166 23548
rect 24670 23536 24676 23548
rect 24728 23536 24734 23588
rect 27154 23576 27160 23588
rect 24780 23548 27160 23576
rect 1946 23508 1952 23520
rect 1907 23480 1952 23508
rect 1946 23468 1952 23480
rect 2004 23468 2010 23520
rect 9858 23468 9864 23520
rect 9916 23508 9922 23520
rect 10229 23511 10287 23517
rect 10229 23508 10241 23511
rect 9916 23480 10241 23508
rect 9916 23468 9922 23480
rect 10229 23477 10241 23480
rect 10275 23477 10287 23511
rect 10229 23471 10287 23477
rect 11514 23468 11520 23520
rect 11572 23508 11578 23520
rect 11977 23511 12035 23517
rect 11977 23508 11989 23511
rect 11572 23480 11989 23508
rect 11572 23468 11578 23480
rect 11977 23477 11989 23480
rect 12023 23477 12035 23511
rect 11977 23471 12035 23477
rect 14645 23511 14703 23517
rect 14645 23477 14657 23511
rect 14691 23508 14703 23511
rect 14826 23508 14832 23520
rect 14691 23480 14832 23508
rect 14691 23477 14703 23480
rect 14645 23471 14703 23477
rect 14826 23468 14832 23480
rect 14884 23468 14890 23520
rect 15286 23468 15292 23520
rect 15344 23508 15350 23520
rect 15562 23508 15568 23520
rect 15344 23480 15568 23508
rect 15344 23468 15350 23480
rect 15562 23468 15568 23480
rect 15620 23468 15626 23520
rect 17034 23468 17040 23520
rect 17092 23508 17098 23520
rect 17865 23511 17923 23517
rect 17865 23508 17877 23511
rect 17092 23480 17877 23508
rect 17092 23468 17098 23480
rect 17865 23477 17877 23480
rect 17911 23477 17923 23511
rect 17865 23471 17923 23477
rect 18322 23468 18328 23520
rect 18380 23508 18386 23520
rect 20806 23508 20812 23520
rect 18380 23480 20812 23508
rect 18380 23468 18386 23480
rect 20806 23468 20812 23480
rect 20864 23508 20870 23520
rect 24780 23508 24808 23548
rect 27154 23536 27160 23548
rect 27212 23536 27218 23588
rect 20864 23480 24808 23508
rect 20864 23468 20870 23480
rect 25130 23468 25136 23520
rect 25188 23508 25194 23520
rect 29825 23511 29883 23517
rect 29825 23508 29837 23511
rect 25188 23480 29837 23508
rect 25188 23468 25194 23480
rect 29825 23477 29837 23480
rect 29871 23477 29883 23511
rect 29825 23471 29883 23477
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 17957 23307 18015 23313
rect 17957 23273 17969 23307
rect 18003 23304 18015 23307
rect 23382 23304 23388 23316
rect 18003 23276 23388 23304
rect 18003 23273 18015 23276
rect 17957 23267 18015 23273
rect 23382 23264 23388 23276
rect 23440 23264 23446 23316
rect 29546 23304 29552 23316
rect 23492 23276 29552 23304
rect 23492 23236 23520 23276
rect 29546 23264 29552 23276
rect 29604 23264 29610 23316
rect 20180 23208 23520 23236
rect 10226 23168 10232 23180
rect 10187 23140 10232 23168
rect 10226 23128 10232 23140
rect 10284 23128 10290 23180
rect 11241 23171 11299 23177
rect 11241 23137 11253 23171
rect 11287 23168 11299 23171
rect 13354 23168 13360 23180
rect 11287 23140 13360 23168
rect 11287 23137 11299 23140
rect 11241 23131 11299 23137
rect 13354 23128 13360 23140
rect 13412 23128 13418 23180
rect 13446 23128 13452 23180
rect 13504 23168 13510 23180
rect 15013 23171 15071 23177
rect 15013 23168 15025 23171
rect 13504 23140 15025 23168
rect 13504 23128 13510 23140
rect 15013 23137 15025 23140
rect 15059 23137 15071 23171
rect 15013 23131 15071 23137
rect 16945 23171 17003 23177
rect 16945 23137 16957 23171
rect 16991 23168 17003 23171
rect 17034 23168 17040 23180
rect 16991 23140 17040 23168
rect 16991 23137 17003 23140
rect 16945 23131 17003 23137
rect 17034 23128 17040 23140
rect 17092 23128 17098 23180
rect 18966 23128 18972 23180
rect 19024 23168 19030 23180
rect 20180 23177 20208 23208
rect 24670 23196 24676 23248
rect 24728 23196 24734 23248
rect 20165 23171 20223 23177
rect 20165 23168 20177 23171
rect 19024 23140 20177 23168
rect 19024 23128 19030 23140
rect 20165 23137 20177 23140
rect 20211 23137 20223 23171
rect 20165 23131 20223 23137
rect 21085 23171 21143 23177
rect 21085 23137 21097 23171
rect 21131 23168 21143 23171
rect 23290 23168 23296 23180
rect 21131 23140 23296 23168
rect 21131 23137 21143 23140
rect 21085 23131 21143 23137
rect 23290 23128 23296 23140
rect 23348 23128 23354 23180
rect 24688 23168 24716 23196
rect 24765 23171 24823 23177
rect 24765 23168 24777 23171
rect 24688 23140 24777 23168
rect 24765 23137 24777 23140
rect 24811 23137 24823 23171
rect 24765 23131 24823 23137
rect 11882 23060 11888 23112
rect 11940 23100 11946 23112
rect 12253 23103 12311 23109
rect 12253 23100 12265 23103
rect 11940 23072 12265 23100
rect 11940 23060 11946 23072
rect 12253 23069 12265 23072
rect 12299 23069 12311 23103
rect 13372 23100 13400 23128
rect 13906 23100 13912 23112
rect 13372 23072 13912 23100
rect 12253 23063 12311 23069
rect 13906 23060 13912 23072
rect 13964 23060 13970 23112
rect 15838 23100 15844 23112
rect 15799 23072 15844 23100
rect 15838 23060 15844 23072
rect 15896 23060 15902 23112
rect 16482 23060 16488 23112
rect 16540 23100 16546 23112
rect 16761 23103 16819 23109
rect 16761 23100 16773 23103
rect 16540 23072 16773 23100
rect 16540 23060 16546 23072
rect 16761 23069 16773 23072
rect 16807 23069 16819 23103
rect 16761 23063 16819 23069
rect 17865 23103 17923 23109
rect 17865 23069 17877 23103
rect 17911 23069 17923 23103
rect 17865 23063 17923 23069
rect 10318 22992 10324 23044
rect 10376 23032 10382 23044
rect 14737 23035 14795 23041
rect 10376 23004 10421 23032
rect 10376 22992 10382 23004
rect 14737 23001 14749 23035
rect 14783 23001 14795 23035
rect 14737 22995 14795 23001
rect 9493 22967 9551 22973
rect 9493 22933 9505 22967
rect 9539 22964 9551 22967
rect 9766 22964 9772 22976
rect 9539 22936 9772 22964
rect 9539 22933 9551 22936
rect 9493 22927 9551 22933
rect 9766 22924 9772 22936
rect 9824 22924 9830 22976
rect 12342 22964 12348 22976
rect 12303 22936 12348 22964
rect 12342 22924 12348 22936
rect 12400 22924 12406 22976
rect 14752 22964 14780 22995
rect 14826 22992 14832 23044
rect 14884 23032 14890 23044
rect 15746 23032 15752 23044
rect 14884 23004 14929 23032
rect 15580 23004 15752 23032
rect 14884 22992 14890 23004
rect 15580 22964 15608 23004
rect 15746 22992 15752 23004
rect 15804 22992 15810 23044
rect 16022 22992 16028 23044
rect 16080 23032 16086 23044
rect 17880 23032 17908 23063
rect 16080 23004 17908 23032
rect 19889 23035 19947 23041
rect 16080 22992 16086 23004
rect 19889 23001 19901 23035
rect 19935 23001 19947 23035
rect 19889 22995 19947 23001
rect 19981 23035 20039 23041
rect 19981 23001 19993 23035
rect 20027 23032 20039 23035
rect 20027 23004 20484 23032
rect 20027 23001 20039 23004
rect 19981 22995 20039 23001
rect 14752 22936 15608 22964
rect 15654 22924 15660 22976
rect 15712 22964 15718 22976
rect 15933 22967 15991 22973
rect 15933 22964 15945 22967
rect 15712 22936 15945 22964
rect 15712 22924 15718 22936
rect 15933 22933 15945 22936
rect 15979 22933 15991 22967
rect 15933 22927 15991 22933
rect 17405 22967 17463 22973
rect 17405 22933 17417 22967
rect 17451 22964 17463 22967
rect 19426 22964 19432 22976
rect 17451 22936 19432 22964
rect 17451 22933 17463 22936
rect 17405 22927 17463 22933
rect 19426 22924 19432 22936
rect 19484 22924 19490 22976
rect 19904 22964 19932 22995
rect 20346 22964 20352 22976
rect 19904 22936 20352 22964
rect 20346 22924 20352 22936
rect 20404 22924 20410 22976
rect 20456 22964 20484 23004
rect 21174 22992 21180 23044
rect 21232 23032 21238 23044
rect 21232 23004 21277 23032
rect 21232 22992 21238 23004
rect 21358 22992 21364 23044
rect 21416 23032 21422 23044
rect 22097 23035 22155 23041
rect 22097 23032 22109 23035
rect 21416 23004 22109 23032
rect 21416 22992 21422 23004
rect 22097 23001 22109 23004
rect 22143 23001 22155 23035
rect 22097 22995 22155 23001
rect 24857 23035 24915 23041
rect 24857 23001 24869 23035
rect 24903 23032 24915 23035
rect 25038 23032 25044 23044
rect 24903 23004 25044 23032
rect 24903 23001 24915 23004
rect 24857 22995 24915 23001
rect 25038 22992 25044 23004
rect 25096 22992 25102 23044
rect 25409 23035 25467 23041
rect 25409 23001 25421 23035
rect 25455 23001 25467 23035
rect 25409 22995 25467 23001
rect 21910 22964 21916 22976
rect 20456 22936 21916 22964
rect 21910 22924 21916 22936
rect 21968 22924 21974 22976
rect 22370 22924 22376 22976
rect 22428 22964 22434 22976
rect 25424 22964 25452 22995
rect 22428 22936 25452 22964
rect 22428 22924 22434 22936
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 2038 22720 2044 22772
rect 2096 22760 2102 22772
rect 9033 22763 9091 22769
rect 9033 22760 9045 22763
rect 2096 22732 9045 22760
rect 2096 22720 2102 22732
rect 9033 22729 9045 22732
rect 9079 22729 9091 22763
rect 11885 22763 11943 22769
rect 9033 22723 9091 22729
rect 9600 22732 10088 22760
rect 7285 22695 7343 22701
rect 7285 22692 7297 22695
rect 7024 22664 7297 22692
rect 1762 22624 1768 22636
rect 1723 22596 1768 22624
rect 1762 22584 1768 22596
rect 1820 22584 1826 22636
rect 7024 22488 7052 22664
rect 7285 22661 7297 22664
rect 7331 22661 7343 22695
rect 7285 22655 7343 22661
rect 7837 22695 7895 22701
rect 7837 22661 7849 22695
rect 7883 22692 7895 22695
rect 9600 22692 9628 22732
rect 9766 22692 9772 22704
rect 7883 22664 9628 22692
rect 9727 22664 9772 22692
rect 7883 22661 7895 22664
rect 7837 22655 7895 22661
rect 9766 22652 9772 22664
rect 9824 22652 9830 22704
rect 9858 22652 9864 22704
rect 9916 22692 9922 22704
rect 10060 22692 10088 22732
rect 11885 22729 11897 22763
rect 11931 22760 11943 22763
rect 12986 22760 12992 22772
rect 11931 22732 12992 22760
rect 11931 22729 11943 22732
rect 11885 22723 11943 22729
rect 12986 22720 12992 22732
rect 13044 22720 13050 22772
rect 14642 22720 14648 22772
rect 14700 22760 14706 22772
rect 15197 22763 15255 22769
rect 15197 22760 15209 22763
rect 14700 22732 15209 22760
rect 14700 22720 14706 22732
rect 15197 22729 15209 22732
rect 15243 22729 15255 22763
rect 20346 22760 20352 22772
rect 20307 22732 20352 22760
rect 15197 22723 15255 22729
rect 20346 22720 20352 22732
rect 20404 22720 20410 22772
rect 22097 22763 22155 22769
rect 22097 22729 22109 22763
rect 22143 22760 22155 22763
rect 22186 22760 22192 22772
rect 22143 22732 22192 22760
rect 22143 22729 22155 22732
rect 22097 22723 22155 22729
rect 22186 22720 22192 22732
rect 22244 22720 22250 22772
rect 25038 22760 25044 22772
rect 24999 22732 25044 22760
rect 25038 22720 25044 22732
rect 25096 22720 25102 22772
rect 30745 22763 30803 22769
rect 30745 22729 30757 22763
rect 30791 22760 30803 22763
rect 32398 22760 32404 22772
rect 30791 22732 32404 22760
rect 30791 22729 30803 22732
rect 30745 22723 30803 22729
rect 32398 22720 32404 22732
rect 32456 22720 32462 22772
rect 12434 22692 12440 22704
rect 9916 22664 9961 22692
rect 10060 22664 12440 22692
rect 9916 22652 9922 22664
rect 12434 22652 12440 22664
rect 12492 22692 12498 22704
rect 13354 22692 13360 22704
rect 12492 22664 13360 22692
rect 12492 22652 12498 22664
rect 13354 22652 13360 22664
rect 13412 22652 13418 22704
rect 13449 22695 13507 22701
rect 13449 22661 13461 22695
rect 13495 22692 13507 22695
rect 14366 22692 14372 22704
rect 13495 22664 14372 22692
rect 13495 22661 13507 22664
rect 13449 22655 13507 22661
rect 14366 22652 14372 22664
rect 14424 22652 14430 22704
rect 17218 22692 17224 22704
rect 17179 22664 17224 22692
rect 17218 22652 17224 22664
rect 17276 22652 17282 22704
rect 19426 22652 19432 22704
rect 19484 22692 19490 22704
rect 24854 22692 24860 22704
rect 19484 22664 24860 22692
rect 19484 22652 19490 22664
rect 24854 22652 24860 22664
rect 24912 22652 24918 22704
rect 27246 22692 27252 22704
rect 27207 22664 27252 22692
rect 27246 22652 27252 22664
rect 27304 22652 27310 22704
rect 27338 22652 27344 22704
rect 27396 22692 27402 22704
rect 27396 22664 27441 22692
rect 27396 22652 27402 22664
rect 9217 22627 9275 22633
rect 9217 22593 9229 22627
rect 9263 22593 9275 22627
rect 10870 22624 10876 22636
rect 10831 22596 10876 22624
rect 9217 22587 9275 22593
rect 7193 22559 7251 22565
rect 7193 22525 7205 22559
rect 7239 22556 7251 22559
rect 7558 22556 7564 22568
rect 7239 22528 7564 22556
rect 7239 22525 7251 22528
rect 7193 22519 7251 22525
rect 7558 22516 7564 22528
rect 7616 22516 7622 22568
rect 8570 22488 8576 22500
rect 7024 22460 8576 22488
rect 8570 22448 8576 22460
rect 8628 22448 8634 22500
rect 9232 22488 9260 22587
rect 10870 22584 10876 22596
rect 10928 22624 10934 22636
rect 11793 22627 11851 22633
rect 11793 22624 11805 22627
rect 10928 22596 11805 22624
rect 10928 22584 10934 22596
rect 11793 22593 11805 22596
rect 11839 22593 11851 22627
rect 14734 22624 14740 22636
rect 14695 22596 14740 22624
rect 11793 22587 11851 22593
rect 14734 22584 14740 22596
rect 14792 22584 14798 22636
rect 14918 22584 14924 22636
rect 14976 22624 14982 22636
rect 16117 22627 16175 22633
rect 16117 22624 16129 22627
rect 14976 22596 16129 22624
rect 14976 22584 14982 22596
rect 16117 22593 16129 22596
rect 16163 22593 16175 22627
rect 18598 22624 18604 22636
rect 18559 22596 18604 22624
rect 16117 22587 16175 22593
rect 18598 22584 18604 22596
rect 18656 22624 18662 22636
rect 22005 22627 22063 22633
rect 22005 22624 22017 22627
rect 18656 22596 22017 22624
rect 18656 22584 18662 22596
rect 22005 22593 22017 22596
rect 22051 22593 22063 22627
rect 22005 22587 22063 22593
rect 24949 22627 25007 22633
rect 24949 22593 24961 22627
rect 24995 22624 25007 22627
rect 25038 22624 25044 22636
rect 24995 22596 25044 22624
rect 24995 22593 25007 22596
rect 24949 22587 25007 22593
rect 25038 22584 25044 22596
rect 25096 22584 25102 22636
rect 26145 22627 26203 22633
rect 26145 22593 26157 22627
rect 26191 22593 26203 22627
rect 26145 22587 26203 22593
rect 30469 22627 30527 22633
rect 30469 22593 30481 22627
rect 30515 22624 30527 22627
rect 30926 22624 30932 22636
rect 30515 22596 30932 22624
rect 30515 22593 30527 22596
rect 30469 22587 30527 22593
rect 10413 22559 10471 22565
rect 10413 22525 10425 22559
rect 10459 22556 10471 22559
rect 11606 22556 11612 22568
rect 10459 22528 11612 22556
rect 10459 22525 10471 22528
rect 10413 22519 10471 22525
rect 11606 22516 11612 22528
rect 11664 22516 11670 22568
rect 13357 22559 13415 22565
rect 13357 22525 13369 22559
rect 13403 22525 13415 22559
rect 13357 22519 13415 22525
rect 11698 22488 11704 22500
rect 9232 22460 11704 22488
rect 11698 22448 11704 22460
rect 11756 22448 11762 22500
rect 13372 22488 13400 22519
rect 13722 22516 13728 22568
rect 13780 22556 13786 22568
rect 13817 22559 13875 22565
rect 13817 22556 13829 22559
rect 13780 22528 13829 22556
rect 13780 22516 13786 22528
rect 13817 22525 13829 22528
rect 13863 22525 13875 22559
rect 14550 22556 14556 22568
rect 14511 22528 14556 22556
rect 13817 22519 13875 22525
rect 14550 22516 14556 22528
rect 14608 22516 14614 22568
rect 16206 22516 16212 22568
rect 16264 22556 16270 22568
rect 17129 22559 17187 22565
rect 17129 22556 17141 22559
rect 16264 22528 17141 22556
rect 16264 22516 16270 22528
rect 17129 22525 17141 22528
rect 17175 22525 17187 22559
rect 17954 22556 17960 22568
rect 17915 22528 17960 22556
rect 17129 22519 17187 22525
rect 17954 22516 17960 22528
rect 18012 22516 18018 22568
rect 19242 22516 19248 22568
rect 19300 22556 19306 22568
rect 21358 22556 21364 22568
rect 19300 22528 21364 22556
rect 19300 22516 19306 22528
rect 21358 22516 21364 22528
rect 21416 22516 21422 22568
rect 24762 22516 24768 22568
rect 24820 22556 24826 22568
rect 26160 22556 26188 22587
rect 30926 22584 30932 22596
rect 30984 22584 30990 22636
rect 38010 22624 38016 22636
rect 37971 22596 38016 22624
rect 38010 22584 38016 22596
rect 38068 22584 38074 22636
rect 24820 22528 26188 22556
rect 24820 22516 24826 22528
rect 26878 22516 26884 22568
rect 26936 22556 26942 22568
rect 27525 22559 27583 22565
rect 27525 22556 27537 22559
rect 26936 22528 27537 22556
rect 26936 22516 26942 22528
rect 27525 22525 27537 22528
rect 27571 22525 27583 22559
rect 27525 22519 27583 22525
rect 16114 22488 16120 22500
rect 13372 22460 16120 22488
rect 16114 22448 16120 22460
rect 16172 22488 16178 22500
rect 16482 22488 16488 22500
rect 16172 22460 16488 22488
rect 16172 22448 16178 22460
rect 16482 22448 16488 22460
rect 16540 22448 16546 22500
rect 38194 22488 38200 22500
rect 38155 22460 38200 22488
rect 38194 22448 38200 22460
rect 38252 22448 38258 22500
rect 1581 22423 1639 22429
rect 1581 22389 1593 22423
rect 1627 22420 1639 22423
rect 8294 22420 8300 22432
rect 1627 22392 8300 22420
rect 1627 22389 1639 22392
rect 1581 22383 1639 22389
rect 8294 22380 8300 22392
rect 8352 22380 8358 22432
rect 10134 22380 10140 22432
rect 10192 22420 10198 22432
rect 10965 22423 11023 22429
rect 10965 22420 10977 22423
rect 10192 22392 10977 22420
rect 10192 22380 10198 22392
rect 10965 22389 10977 22392
rect 11011 22389 11023 22423
rect 10965 22383 11023 22389
rect 16209 22423 16267 22429
rect 16209 22389 16221 22423
rect 16255 22420 16267 22423
rect 16574 22420 16580 22432
rect 16255 22392 16580 22420
rect 16255 22389 16267 22392
rect 16209 22383 16267 22389
rect 16574 22380 16580 22392
rect 16632 22380 16638 22432
rect 17954 22380 17960 22432
rect 18012 22420 18018 22432
rect 18693 22423 18751 22429
rect 18693 22420 18705 22423
rect 18012 22392 18705 22420
rect 18012 22380 18018 22392
rect 18693 22389 18705 22392
rect 18739 22389 18751 22423
rect 18693 22383 18751 22389
rect 26237 22423 26295 22429
rect 26237 22389 26249 22423
rect 26283 22420 26295 22423
rect 27062 22420 27068 22432
rect 26283 22392 27068 22420
rect 26283 22389 26295 22392
rect 26237 22383 26295 22389
rect 27062 22380 27068 22392
rect 27120 22380 27126 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 8846 22176 8852 22228
rect 8904 22216 8910 22228
rect 10042 22216 10048 22228
rect 8904 22188 10048 22216
rect 8904 22176 8910 22188
rect 10042 22176 10048 22188
rect 10100 22216 10106 22228
rect 10870 22216 10876 22228
rect 10100 22188 10876 22216
rect 10100 22176 10106 22188
rect 10870 22176 10876 22188
rect 10928 22176 10934 22228
rect 19702 22216 19708 22228
rect 17696 22188 19708 22216
rect 8202 22108 8208 22160
rect 8260 22148 8266 22160
rect 13722 22148 13728 22160
rect 8260 22120 13728 22148
rect 8260 22108 8266 22120
rect 13722 22108 13728 22120
rect 13780 22108 13786 22160
rect 16022 22148 16028 22160
rect 14568 22120 16028 22148
rect 7006 22080 7012 22092
rect 6967 22052 7012 22080
rect 7006 22040 7012 22052
rect 7064 22040 7070 22092
rect 11606 22040 11612 22092
rect 11664 22080 11670 22092
rect 11701 22083 11759 22089
rect 11701 22080 11713 22083
rect 11664 22052 11713 22080
rect 11664 22040 11670 22052
rect 11701 22049 11713 22052
rect 11747 22049 11759 22083
rect 14366 22080 14372 22092
rect 14327 22052 14372 22080
rect 11701 22043 11759 22049
rect 14366 22040 14372 22052
rect 14424 22040 14430 22092
rect 6917 22015 6975 22021
rect 6917 21981 6929 22015
rect 6963 22012 6975 22015
rect 7098 22012 7104 22024
rect 6963 21984 7104 22012
rect 6963 21981 6975 21984
rect 6917 21975 6975 21981
rect 7098 21972 7104 21984
rect 7156 21972 7162 22024
rect 8021 22015 8079 22021
rect 8021 21981 8033 22015
rect 8067 21981 8079 22015
rect 8021 21975 8079 21981
rect 8036 21944 8064 21975
rect 8294 21972 8300 22024
rect 8352 22012 8358 22024
rect 9125 22015 9183 22021
rect 9125 22012 9137 22015
rect 8352 21984 9137 22012
rect 8352 21972 8358 21984
rect 9125 21981 9137 21984
rect 9171 21981 9183 22015
rect 9125 21975 9183 21981
rect 13998 21972 14004 22024
rect 14056 22012 14062 22024
rect 14277 22015 14335 22021
rect 14277 22012 14289 22015
rect 14056 21984 14289 22012
rect 14056 21972 14062 21984
rect 14277 21981 14289 21984
rect 14323 22012 14335 22015
rect 14568 22012 14596 22120
rect 16022 22108 16028 22120
rect 16080 22108 16086 22160
rect 17218 22108 17224 22160
rect 17276 22148 17282 22160
rect 17696 22148 17724 22188
rect 19702 22176 19708 22188
rect 19760 22176 19766 22228
rect 26329 22219 26387 22225
rect 26329 22185 26341 22219
rect 26375 22216 26387 22219
rect 27338 22216 27344 22228
rect 26375 22188 27344 22216
rect 26375 22185 26387 22188
rect 26329 22179 26387 22185
rect 27338 22176 27344 22188
rect 27396 22176 27402 22228
rect 17276 22120 17724 22148
rect 17276 22108 17282 22120
rect 17604 22089 17632 22120
rect 17862 22108 17868 22160
rect 17920 22148 17926 22160
rect 25038 22148 25044 22160
rect 17920 22120 25044 22148
rect 17920 22108 17926 22120
rect 17589 22083 17647 22089
rect 14323 21984 14596 22012
rect 14660 22052 16528 22080
rect 14323 21981 14335 21984
rect 14277 21975 14335 21981
rect 9030 21944 9036 21956
rect 8036 21916 9036 21944
rect 9030 21904 9036 21916
rect 9088 21904 9094 21956
rect 9217 21947 9275 21953
rect 9217 21913 9229 21947
rect 9263 21944 9275 21947
rect 10045 21947 10103 21953
rect 10045 21944 10057 21947
rect 9263 21916 10057 21944
rect 9263 21913 9275 21916
rect 9217 21907 9275 21913
rect 10045 21913 10057 21916
rect 10091 21913 10103 21947
rect 10045 21907 10103 21913
rect 10134 21904 10140 21956
rect 10192 21944 10198 21956
rect 10689 21947 10747 21953
rect 10192 21916 10237 21944
rect 10192 21904 10198 21916
rect 10689 21913 10701 21947
rect 10735 21913 10747 21947
rect 10689 21907 10747 21913
rect 7466 21836 7472 21888
rect 7524 21876 7530 21888
rect 8113 21879 8171 21885
rect 8113 21876 8125 21879
rect 7524 21848 8125 21876
rect 7524 21836 7530 21848
rect 8113 21845 8125 21848
rect 8159 21845 8171 21879
rect 10704 21876 10732 21907
rect 10870 21904 10876 21956
rect 10928 21944 10934 21956
rect 11425 21947 11483 21953
rect 11425 21944 11437 21947
rect 10928 21916 11437 21944
rect 10928 21904 10934 21916
rect 11425 21913 11437 21916
rect 11471 21913 11483 21947
rect 11425 21907 11483 21913
rect 11514 21904 11520 21956
rect 11572 21944 11578 21956
rect 11572 21916 11617 21944
rect 11572 21904 11578 21916
rect 12526 21904 12532 21956
rect 12584 21944 12590 21956
rect 14660 21944 14688 22052
rect 16500 22024 16528 22052
rect 17589 22049 17601 22083
rect 17635 22049 17647 22083
rect 17954 22080 17960 22092
rect 17915 22052 17960 22080
rect 17589 22043 17647 22049
rect 17954 22040 17960 22052
rect 18012 22040 18018 22092
rect 19628 22080 19656 22120
rect 25038 22108 25044 22120
rect 25096 22148 25102 22160
rect 25406 22148 25412 22160
rect 25096 22120 25412 22148
rect 25096 22108 25102 22120
rect 25406 22108 25412 22120
rect 25464 22108 25470 22160
rect 27522 22148 27528 22160
rect 27483 22120 27528 22148
rect 27522 22108 27528 22120
rect 27580 22108 27586 22160
rect 19536 22052 19656 22080
rect 15378 22012 15384 22024
rect 15339 21984 15384 22012
rect 15378 21972 15384 21984
rect 15436 21972 15442 22024
rect 15838 22012 15844 22024
rect 15799 21984 15844 22012
rect 15838 21972 15844 21984
rect 15896 21972 15902 22024
rect 16114 22012 16120 22024
rect 15948 21984 16120 22012
rect 15194 21944 15200 21956
rect 12584 21916 14688 21944
rect 15155 21916 15200 21944
rect 12584 21904 12590 21916
rect 15194 21904 15200 21916
rect 15252 21904 15258 21956
rect 15948 21953 15976 21984
rect 16114 21972 16120 21984
rect 16172 21972 16178 22024
rect 16482 21972 16488 22024
rect 16540 21972 16546 22024
rect 16850 22012 16856 22024
rect 16811 21984 16856 22012
rect 16850 21972 16856 21984
rect 16908 21972 16914 22024
rect 19536 22021 19564 22052
rect 20254 22040 20260 22092
rect 20312 22080 20318 22092
rect 28258 22080 28264 22092
rect 20312 22052 28264 22080
rect 20312 22040 20318 22052
rect 28258 22040 28264 22052
rect 28316 22040 28322 22092
rect 19521 22015 19579 22021
rect 19521 21981 19533 22015
rect 19567 21981 19579 22015
rect 19521 21975 19579 21981
rect 20898 21972 20904 22024
rect 20956 22012 20962 22024
rect 24581 22015 24639 22021
rect 24581 22012 24593 22015
rect 20956 21984 24593 22012
rect 20956 21972 20962 21984
rect 24581 21981 24593 21984
rect 24627 22012 24639 22015
rect 26237 22015 26295 22021
rect 26237 22012 26249 22015
rect 24627 21984 26249 22012
rect 24627 21981 24639 21984
rect 24581 21975 24639 21981
rect 26237 21981 26249 21984
rect 26283 21981 26295 22015
rect 26237 21975 26295 21981
rect 34790 21972 34796 22024
rect 34848 22012 34854 22024
rect 34885 22015 34943 22021
rect 34885 22012 34897 22015
rect 34848 21984 34897 22012
rect 34848 21972 34854 21984
rect 34885 21981 34897 21984
rect 34931 21981 34943 22015
rect 34885 21975 34943 21981
rect 34977 22015 35035 22021
rect 34977 21981 34989 22015
rect 35023 22012 35035 22015
rect 37553 22015 37611 22021
rect 37553 22012 37565 22015
rect 35023 21984 37565 22012
rect 35023 21981 35035 21984
rect 34977 21975 35035 21981
rect 37553 21981 37565 21984
rect 37599 21981 37611 22015
rect 37553 21975 37611 21981
rect 38013 22015 38071 22021
rect 38013 21981 38025 22015
rect 38059 21981 38071 22015
rect 38013 21975 38071 21981
rect 15933 21947 15991 21953
rect 15304 21916 15792 21944
rect 12986 21876 12992 21888
rect 10704 21848 12992 21876
rect 8113 21839 8171 21845
rect 12986 21836 12992 21848
rect 13044 21836 13050 21888
rect 13170 21836 13176 21888
rect 13228 21876 13234 21888
rect 15304 21876 15332 21916
rect 13228 21848 15332 21876
rect 15764 21876 15792 21916
rect 15933 21913 15945 21947
rect 15979 21913 15991 21947
rect 17681 21947 17739 21953
rect 15933 21907 15991 21913
rect 16040 21916 17632 21944
rect 16040 21876 16068 21916
rect 15764 21848 16068 21876
rect 13228 21836 13234 21848
rect 16114 21836 16120 21888
rect 16172 21876 16178 21888
rect 16945 21879 17003 21885
rect 16945 21876 16957 21879
rect 16172 21848 16957 21876
rect 16172 21836 16178 21848
rect 16945 21845 16957 21848
rect 16991 21845 17003 21879
rect 17604 21876 17632 21916
rect 17681 21913 17693 21947
rect 17727 21944 17739 21947
rect 17770 21944 17776 21956
rect 17727 21916 17776 21944
rect 17727 21913 17739 21916
rect 17681 21907 17739 21913
rect 17770 21904 17776 21916
rect 17828 21904 17834 21956
rect 22370 21944 22376 21956
rect 17880 21916 22376 21944
rect 17880 21876 17908 21916
rect 22370 21904 22376 21916
rect 22428 21944 22434 21956
rect 22830 21944 22836 21956
rect 22428 21916 22836 21944
rect 22428 21904 22434 21916
rect 22830 21904 22836 21916
rect 22888 21904 22894 21956
rect 26970 21944 26976 21956
rect 26931 21916 26976 21944
rect 26970 21904 26976 21916
rect 27028 21904 27034 21956
rect 27062 21904 27068 21956
rect 27120 21944 27126 21956
rect 38028 21944 38056 21975
rect 27120 21916 27165 21944
rect 37384 21916 38056 21944
rect 27120 21904 27126 21916
rect 17604 21848 17908 21876
rect 16945 21839 17003 21845
rect 19426 21836 19432 21888
rect 19484 21876 19490 21888
rect 19613 21879 19671 21885
rect 19613 21876 19625 21879
rect 19484 21848 19625 21876
rect 19484 21836 19490 21848
rect 19613 21845 19625 21848
rect 19659 21845 19671 21879
rect 19613 21839 19671 21845
rect 19702 21836 19708 21888
rect 19760 21876 19766 21888
rect 23474 21876 23480 21888
rect 19760 21848 23480 21876
rect 19760 21836 19766 21848
rect 23474 21836 23480 21848
rect 23532 21836 23538 21888
rect 23566 21836 23572 21888
rect 23624 21876 23630 21888
rect 37384 21885 37412 21916
rect 24673 21879 24731 21885
rect 24673 21876 24685 21879
rect 23624 21848 24685 21876
rect 23624 21836 23630 21848
rect 24673 21845 24685 21848
rect 24719 21845 24731 21879
rect 24673 21839 24731 21845
rect 37369 21879 37427 21885
rect 37369 21845 37381 21879
rect 37415 21845 37427 21879
rect 38194 21876 38200 21888
rect 38155 21848 38200 21876
rect 37369 21839 37427 21845
rect 38194 21836 38200 21848
rect 38252 21836 38258 21888
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 8570 21672 8576 21684
rect 8531 21644 8576 21672
rect 8570 21632 8576 21644
rect 8628 21632 8634 21684
rect 8754 21632 8760 21684
rect 8812 21672 8818 21684
rect 15194 21672 15200 21684
rect 8812 21644 15200 21672
rect 8812 21632 8818 21644
rect 5445 21607 5503 21613
rect 5445 21573 5457 21607
rect 5491 21604 5503 21607
rect 6730 21604 6736 21616
rect 5491 21576 6736 21604
rect 5491 21573 5503 21576
rect 5445 21567 5503 21573
rect 6730 21564 6736 21576
rect 6788 21564 6794 21616
rect 7374 21604 7380 21616
rect 7335 21576 7380 21604
rect 7374 21564 7380 21576
rect 7432 21564 7438 21616
rect 7466 21564 7472 21616
rect 7524 21604 7530 21616
rect 10686 21604 10692 21616
rect 7524 21576 7569 21604
rect 8496 21576 10692 21604
rect 7524 21564 7530 21576
rect 1670 21536 1676 21548
rect 1631 21508 1676 21536
rect 1670 21496 1676 21508
rect 1728 21496 1734 21548
rect 5997 21539 6055 21545
rect 5997 21505 6009 21539
rect 6043 21536 6055 21539
rect 7098 21536 7104 21548
rect 6043 21508 7104 21536
rect 6043 21505 6055 21508
rect 5997 21499 6055 21505
rect 7098 21496 7104 21508
rect 7156 21496 7162 21548
rect 8496 21545 8524 21576
rect 10686 21564 10692 21576
rect 10744 21564 10750 21616
rect 12802 21604 12808 21616
rect 12763 21576 12808 21604
rect 12802 21564 12808 21576
rect 12860 21564 12866 21616
rect 8481 21539 8539 21545
rect 8481 21505 8493 21539
rect 8527 21505 8539 21539
rect 8481 21499 8539 21505
rect 9125 21539 9183 21545
rect 9125 21505 9137 21539
rect 9171 21536 9183 21539
rect 11606 21536 11612 21548
rect 9171 21508 11612 21536
rect 9171 21505 9183 21508
rect 9125 21499 9183 21505
rect 11606 21496 11612 21508
rect 11664 21496 11670 21548
rect 14108 21545 14136 21644
rect 15194 21632 15200 21644
rect 15252 21632 15258 21684
rect 16022 21672 16028 21684
rect 15856 21644 16028 21672
rect 14185 21607 14243 21613
rect 14185 21573 14197 21607
rect 14231 21604 14243 21607
rect 14550 21604 14556 21616
rect 14231 21576 14556 21604
rect 14231 21573 14243 21576
rect 14185 21567 14243 21573
rect 14550 21564 14556 21576
rect 14608 21564 14614 21616
rect 15381 21607 15439 21613
rect 15381 21573 15393 21607
rect 15427 21604 15439 21607
rect 15856 21604 15884 21644
rect 16022 21632 16028 21644
rect 16080 21632 16086 21684
rect 18064 21644 19104 21672
rect 15427 21576 15884 21604
rect 15427 21573 15439 21576
rect 15381 21567 15439 21573
rect 15930 21564 15936 21616
rect 15988 21604 15994 21616
rect 16945 21607 17003 21613
rect 16945 21604 16957 21607
rect 15988 21576 16957 21604
rect 15988 21564 15994 21576
rect 16945 21573 16957 21576
rect 16991 21573 17003 21607
rect 16945 21567 17003 21573
rect 17494 21564 17500 21616
rect 17552 21604 17558 21616
rect 17862 21604 17868 21616
rect 17552 21576 17868 21604
rect 17552 21564 17558 21576
rect 17862 21564 17868 21576
rect 17920 21564 17926 21616
rect 14093 21539 14151 21545
rect 14093 21505 14105 21539
rect 14139 21505 14151 21539
rect 17589 21539 17647 21545
rect 17589 21536 17601 21539
rect 14093 21499 14151 21505
rect 16132 21508 17601 21536
rect 5353 21471 5411 21477
rect 5353 21437 5365 21471
rect 5399 21468 5411 21471
rect 5626 21468 5632 21480
rect 5399 21440 5632 21468
rect 5399 21437 5411 21440
rect 5353 21431 5411 21437
rect 5626 21428 5632 21440
rect 5684 21428 5690 21480
rect 5828 21440 9352 21468
rect 1857 21403 1915 21409
rect 1857 21369 1869 21403
rect 1903 21400 1915 21403
rect 5828 21400 5856 21440
rect 1903 21372 5856 21400
rect 1903 21369 1915 21372
rect 1857 21363 1915 21369
rect 6914 21360 6920 21412
rect 6972 21400 6978 21412
rect 7929 21403 7987 21409
rect 7929 21400 7941 21403
rect 6972 21372 7941 21400
rect 6972 21360 6978 21372
rect 7929 21369 7941 21372
rect 7975 21400 7987 21403
rect 8202 21400 8208 21412
rect 7975 21372 8208 21400
rect 7975 21369 7987 21372
rect 7929 21363 7987 21369
rect 8202 21360 8208 21372
rect 8260 21360 8266 21412
rect 8386 21292 8392 21344
rect 8444 21332 8450 21344
rect 9217 21335 9275 21341
rect 9217 21332 9229 21335
rect 8444 21304 9229 21332
rect 8444 21292 8450 21304
rect 9217 21301 9229 21304
rect 9263 21301 9275 21335
rect 9324 21332 9352 21440
rect 9950 21428 9956 21480
rect 10008 21468 10014 21480
rect 12713 21471 12771 21477
rect 10008 21440 12664 21468
rect 10008 21428 10014 21440
rect 9398 21360 9404 21412
rect 9456 21400 9462 21412
rect 12526 21400 12532 21412
rect 9456 21372 12532 21400
rect 9456 21360 9462 21372
rect 12526 21360 12532 21372
rect 12584 21360 12590 21412
rect 12636 21400 12664 21440
rect 12713 21437 12725 21471
rect 12759 21468 12771 21471
rect 13170 21468 13176 21480
rect 12759 21440 13176 21468
rect 12759 21437 12771 21440
rect 12713 21431 12771 21437
rect 13170 21428 13176 21440
rect 13228 21428 13234 21480
rect 13357 21471 13415 21477
rect 13357 21437 13369 21471
rect 13403 21468 13415 21471
rect 13446 21468 13452 21480
rect 13403 21440 13452 21468
rect 13403 21437 13415 21440
rect 13357 21431 13415 21437
rect 13372 21400 13400 21431
rect 13446 21428 13452 21440
rect 13504 21428 13510 21480
rect 15289 21471 15347 21477
rect 15289 21437 15301 21471
rect 15335 21468 15347 21471
rect 15562 21468 15568 21480
rect 15335 21440 15568 21468
rect 15335 21437 15347 21440
rect 15289 21431 15347 21437
rect 15562 21428 15568 21440
rect 15620 21428 15626 21480
rect 16132 21468 16160 21508
rect 17589 21505 17601 21508
rect 17635 21505 17647 21539
rect 17589 21499 17647 21505
rect 15672 21440 16160 21468
rect 16301 21471 16359 21477
rect 12636 21372 13400 21400
rect 13722 21360 13728 21412
rect 13780 21400 13786 21412
rect 15672 21400 15700 21440
rect 16301 21437 16313 21471
rect 16347 21468 16359 21471
rect 16482 21468 16488 21480
rect 16347 21440 16488 21468
rect 16347 21437 16359 21440
rect 16301 21431 16359 21437
rect 16482 21428 16488 21440
rect 16540 21468 16546 21480
rect 18064 21468 18092 21644
rect 18414 21604 18420 21616
rect 18375 21576 18420 21604
rect 18414 21564 18420 21576
rect 18472 21564 18478 21616
rect 18966 21604 18972 21616
rect 18927 21576 18972 21604
rect 18966 21564 18972 21576
rect 19024 21564 19030 21616
rect 19076 21604 19104 21644
rect 19426 21632 19432 21684
rect 19484 21672 19490 21684
rect 22373 21675 22431 21681
rect 19484 21644 19656 21672
rect 19484 21632 19490 21644
rect 19518 21604 19524 21616
rect 19076 21576 19524 21604
rect 19518 21564 19524 21576
rect 19576 21564 19582 21616
rect 19628 21613 19656 21644
rect 22373 21641 22385 21675
rect 22419 21672 22431 21675
rect 28258 21672 28264 21684
rect 22419 21644 24808 21672
rect 28219 21644 28264 21672
rect 22419 21641 22431 21644
rect 22373 21635 22431 21641
rect 19613 21607 19671 21613
rect 19613 21573 19625 21607
rect 19659 21573 19671 21607
rect 23566 21604 23572 21616
rect 23527 21576 23572 21604
rect 19613 21567 19671 21573
rect 23566 21564 23572 21576
rect 23624 21564 23630 21616
rect 20625 21539 20683 21545
rect 20625 21505 20637 21539
rect 20671 21536 20683 21539
rect 20898 21536 20904 21548
rect 20671 21508 20904 21536
rect 20671 21505 20683 21508
rect 20625 21499 20683 21505
rect 20898 21496 20904 21508
rect 20956 21496 20962 21548
rect 21082 21496 21088 21548
rect 21140 21536 21146 21548
rect 24780 21545 24808 21644
rect 28258 21632 28264 21644
rect 28316 21632 28322 21684
rect 37366 21604 37372 21616
rect 26896 21576 37372 21604
rect 22557 21539 22615 21545
rect 22557 21536 22569 21539
rect 21140 21508 22569 21536
rect 21140 21496 21146 21508
rect 22557 21505 22569 21508
rect 22603 21505 22615 21539
rect 22557 21499 22615 21505
rect 24765 21539 24823 21545
rect 24765 21505 24777 21539
rect 24811 21505 24823 21539
rect 24765 21499 24823 21505
rect 18322 21468 18328 21480
rect 16540 21440 18092 21468
rect 18235 21440 18328 21468
rect 16540 21428 16546 21440
rect 18322 21428 18328 21440
rect 18380 21468 18386 21480
rect 18506 21468 18512 21480
rect 18380 21440 18512 21468
rect 18380 21428 18386 21440
rect 18506 21428 18512 21440
rect 18564 21428 18570 21480
rect 19521 21471 19579 21477
rect 19521 21437 19533 21471
rect 19567 21468 19579 21471
rect 19610 21468 19616 21480
rect 19567 21440 19616 21468
rect 19567 21437 19579 21440
rect 19521 21431 19579 21437
rect 19610 21428 19616 21440
rect 19668 21428 19674 21480
rect 19996 21440 22094 21468
rect 13780 21372 15700 21400
rect 13780 21360 13786 21372
rect 15746 21360 15752 21412
rect 15804 21400 15810 21412
rect 19996 21400 20024 21440
rect 15804 21372 20024 21400
rect 20073 21403 20131 21409
rect 15804 21360 15810 21372
rect 20073 21369 20085 21403
rect 20119 21400 20131 21403
rect 20990 21400 20996 21412
rect 20119 21372 20996 21400
rect 20119 21369 20131 21372
rect 20073 21363 20131 21369
rect 14366 21332 14372 21344
rect 9324 21304 14372 21332
rect 9217 21295 9275 21301
rect 14366 21292 14372 21304
rect 14424 21292 14430 21344
rect 17037 21335 17095 21341
rect 17037 21301 17049 21335
rect 17083 21332 17095 21335
rect 17402 21332 17408 21344
rect 17083 21304 17408 21332
rect 17083 21301 17095 21304
rect 17037 21295 17095 21301
rect 17402 21292 17408 21304
rect 17460 21292 17466 21344
rect 17678 21332 17684 21344
rect 17639 21304 17684 21332
rect 17678 21292 17684 21304
rect 17736 21292 17742 21344
rect 17954 21292 17960 21344
rect 18012 21332 18018 21344
rect 20088 21332 20116 21363
rect 20990 21360 20996 21372
rect 21048 21360 21054 21412
rect 22066 21400 22094 21440
rect 23290 21428 23296 21480
rect 23348 21468 23354 21480
rect 23477 21471 23535 21477
rect 23477 21468 23489 21471
rect 23348 21440 23489 21468
rect 23348 21428 23354 21440
rect 23477 21437 23489 21440
rect 23523 21437 23535 21471
rect 26896 21468 26924 21576
rect 37366 21564 37372 21576
rect 37424 21564 37430 21616
rect 28169 21539 28227 21545
rect 28169 21505 28181 21539
rect 28215 21536 28227 21539
rect 37734 21536 37740 21548
rect 28215 21508 37740 21536
rect 28215 21505 28227 21508
rect 28169 21499 28227 21505
rect 37734 21496 37740 21508
rect 37792 21496 37798 21548
rect 23477 21431 23535 21437
rect 23584 21440 26924 21468
rect 23584 21400 23612 21440
rect 22066 21372 23612 21400
rect 24029 21403 24087 21409
rect 24029 21369 24041 21403
rect 24075 21369 24087 21403
rect 24029 21363 24087 21369
rect 18012 21304 20116 21332
rect 18012 21292 18018 21304
rect 20438 21292 20444 21344
rect 20496 21332 20502 21344
rect 20717 21335 20775 21341
rect 20717 21332 20729 21335
rect 20496 21304 20729 21332
rect 20496 21292 20502 21304
rect 20717 21301 20729 21304
rect 20763 21301 20775 21335
rect 20717 21295 20775 21301
rect 22830 21292 22836 21344
rect 22888 21332 22894 21344
rect 24044 21332 24072 21363
rect 22888 21304 24072 21332
rect 24581 21335 24639 21341
rect 22888 21292 22894 21304
rect 24581 21301 24593 21335
rect 24627 21332 24639 21335
rect 24762 21332 24768 21344
rect 24627 21304 24768 21332
rect 24627 21301 24639 21304
rect 24581 21295 24639 21301
rect 24762 21292 24768 21304
rect 24820 21292 24826 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 2222 21088 2228 21140
rect 2280 21128 2286 21140
rect 15930 21128 15936 21140
rect 2280 21100 15936 21128
rect 2280 21088 2286 21100
rect 15930 21088 15936 21100
rect 15988 21088 15994 21140
rect 18046 21128 18052 21140
rect 16040 21100 18052 21128
rect 9030 21020 9036 21072
rect 9088 21060 9094 21072
rect 13538 21060 13544 21072
rect 9088 21032 13544 21060
rect 9088 21020 9094 21032
rect 13538 21020 13544 21032
rect 13596 21020 13602 21072
rect 15378 21020 15384 21072
rect 15436 21020 15442 21072
rect 4798 20992 4804 21004
rect 4759 20964 4804 20992
rect 4798 20952 4804 20964
rect 4856 20952 4862 21004
rect 5626 20992 5632 21004
rect 5587 20964 5632 20992
rect 5626 20952 5632 20964
rect 5684 20952 5690 21004
rect 9950 20952 9956 21004
rect 10008 20992 10014 21004
rect 10413 20995 10471 21001
rect 10413 20992 10425 20995
rect 10008 20964 10425 20992
rect 10008 20952 10014 20964
rect 10413 20961 10425 20964
rect 10459 20961 10471 20995
rect 10413 20955 10471 20961
rect 11330 20952 11336 21004
rect 11388 20992 11394 21004
rect 12250 20992 12256 21004
rect 11388 20964 12256 20992
rect 11388 20952 11394 20964
rect 12250 20952 12256 20964
rect 12308 20952 12314 21004
rect 13262 20992 13268 21004
rect 13175 20964 13268 20992
rect 13262 20952 13268 20964
rect 13320 20992 13326 21004
rect 15396 20992 15424 21020
rect 16040 20992 16068 21100
rect 18046 21088 18052 21100
rect 18104 21088 18110 21140
rect 22738 21128 22744 21140
rect 18340 21100 22744 21128
rect 18138 21060 18144 21072
rect 16776 21032 18144 21060
rect 13320 20964 16068 20992
rect 16577 20995 16635 21001
rect 13320 20952 13326 20964
rect 16577 20961 16589 20995
rect 16623 20992 16635 20995
rect 16776 20992 16804 21032
rect 18138 21020 18144 21032
rect 18196 21020 18202 21072
rect 16942 20992 16948 21004
rect 16623 20964 16804 20992
rect 16903 20964 16948 20992
rect 16623 20961 16635 20964
rect 16577 20955 16635 20961
rect 16942 20952 16948 20964
rect 17000 20992 17006 21004
rect 18340 20992 18368 21100
rect 22738 21088 22744 21100
rect 22796 21088 22802 21140
rect 28534 21128 28540 21140
rect 22848 21100 28540 21128
rect 18598 21020 18604 21072
rect 18656 21060 18662 21072
rect 22848 21060 22876 21100
rect 28534 21088 28540 21100
rect 28592 21088 28598 21140
rect 37829 21131 37887 21137
rect 37829 21097 37841 21131
rect 37875 21128 37887 21131
rect 38010 21128 38016 21140
rect 37875 21100 38016 21128
rect 37875 21097 37887 21100
rect 37829 21091 37887 21097
rect 38010 21088 38016 21100
rect 38068 21088 38074 21140
rect 18656 21032 22876 21060
rect 18656 21020 18662 21032
rect 22922 21020 22928 21072
rect 22980 21060 22986 21072
rect 23566 21060 23572 21072
rect 22980 21032 23572 21060
rect 22980 21020 22986 21032
rect 23566 21020 23572 21032
rect 23624 21020 23630 21072
rect 23750 21060 23756 21072
rect 23711 21032 23756 21060
rect 23750 21020 23756 21032
rect 23808 21020 23814 21072
rect 17000 20964 18368 20992
rect 18877 20995 18935 21001
rect 17000 20952 17006 20964
rect 18877 20961 18889 20995
rect 18923 20992 18935 20995
rect 18966 20992 18972 21004
rect 18923 20964 18972 20992
rect 18923 20961 18935 20964
rect 18877 20955 18935 20961
rect 18966 20952 18972 20964
rect 19024 20952 19030 21004
rect 19610 20992 19616 21004
rect 19571 20964 19616 20992
rect 19610 20952 19616 20964
rect 19668 20952 19674 21004
rect 20349 20995 20407 21001
rect 20349 20961 20361 20995
rect 20395 20992 20407 20995
rect 21266 20992 21272 21004
rect 20395 20964 21272 20992
rect 20395 20961 20407 20964
rect 20349 20955 20407 20961
rect 21266 20952 21272 20964
rect 21324 20952 21330 21004
rect 23201 20995 23259 21001
rect 23201 20961 23213 20995
rect 23247 20992 23259 20995
rect 25774 20992 25780 21004
rect 23247 20964 25780 20992
rect 23247 20961 23259 20964
rect 23201 20955 23259 20961
rect 25774 20952 25780 20964
rect 25832 20952 25838 21004
rect 1578 20924 1584 20936
rect 1539 20896 1584 20924
rect 1578 20884 1584 20896
rect 1636 20884 1642 20936
rect 1854 20924 1860 20936
rect 1815 20896 1860 20924
rect 1854 20884 1860 20896
rect 1912 20884 1918 20936
rect 6273 20927 6331 20933
rect 6273 20893 6285 20927
rect 6319 20924 6331 20927
rect 7466 20924 7472 20936
rect 6319 20896 7472 20924
rect 6319 20893 6331 20896
rect 6273 20887 6331 20893
rect 7466 20884 7472 20896
rect 7524 20884 7530 20936
rect 8389 20927 8447 20933
rect 8389 20893 8401 20927
rect 8435 20924 8447 20927
rect 9125 20927 9183 20933
rect 9125 20924 9137 20927
rect 8435 20896 9137 20924
rect 8435 20893 8447 20896
rect 8389 20887 8447 20893
rect 9125 20893 9137 20896
rect 9171 20924 9183 20927
rect 9306 20924 9312 20936
rect 9171 20896 9312 20924
rect 9171 20893 9183 20896
rect 9125 20887 9183 20893
rect 9306 20884 9312 20896
rect 9364 20884 9370 20936
rect 13722 20924 13728 20936
rect 13188 20896 13728 20924
rect 4522 20856 4528 20868
rect 4483 20828 4528 20856
rect 4522 20816 4528 20828
rect 4580 20816 4586 20868
rect 4617 20859 4675 20865
rect 4617 20825 4629 20859
rect 4663 20825 4675 20859
rect 4617 20819 4675 20825
rect 4632 20788 4660 20819
rect 7742 20816 7748 20868
rect 7800 20856 7806 20868
rect 8662 20856 8668 20868
rect 7800 20828 8668 20856
rect 7800 20816 7806 20828
rect 8662 20816 8668 20828
rect 8720 20816 8726 20868
rect 10134 20856 10140 20868
rect 10095 20828 10140 20856
rect 10134 20816 10140 20828
rect 10192 20816 10198 20868
rect 10229 20859 10287 20865
rect 10229 20825 10241 20859
rect 10275 20825 10287 20859
rect 12342 20856 12348 20868
rect 12303 20828 12348 20856
rect 10229 20819 10287 20825
rect 6365 20791 6423 20797
rect 6365 20788 6377 20791
rect 4632 20760 6377 20788
rect 6365 20757 6377 20760
rect 6411 20757 6423 20791
rect 8478 20788 8484 20800
rect 8439 20760 8484 20788
rect 6365 20751 6423 20757
rect 8478 20748 8484 20760
rect 8536 20748 8542 20800
rect 9214 20788 9220 20800
rect 9175 20760 9220 20788
rect 9214 20748 9220 20760
rect 9272 20748 9278 20800
rect 9950 20748 9956 20800
rect 10008 20788 10014 20800
rect 10237 20788 10265 20819
rect 12342 20816 12348 20828
rect 12400 20816 12406 20868
rect 12618 20856 12624 20868
rect 12544 20828 12624 20856
rect 10008 20760 10265 20788
rect 10008 20748 10014 20760
rect 10686 20748 10692 20800
rect 10744 20788 10750 20800
rect 12544 20788 12572 20828
rect 12618 20816 12624 20828
rect 12676 20856 12682 20868
rect 13188 20856 13216 20896
rect 13722 20884 13728 20896
rect 13780 20884 13786 20936
rect 19518 20884 19524 20936
rect 19576 20924 19582 20936
rect 20070 20924 20076 20936
rect 19576 20896 20076 20924
rect 19576 20884 19582 20896
rect 20070 20884 20076 20896
rect 20128 20884 20134 20936
rect 20990 20884 20996 20936
rect 21048 20924 21054 20936
rect 22462 20924 22468 20936
rect 21048 20896 21093 20924
rect 22375 20896 22468 20924
rect 21048 20884 21054 20896
rect 22462 20884 22468 20896
rect 22520 20884 22526 20936
rect 22554 20884 22560 20936
rect 22612 20924 22618 20936
rect 25222 20924 25228 20936
rect 22612 20896 22657 20924
rect 25183 20896 25228 20924
rect 22612 20884 22618 20896
rect 25222 20884 25228 20896
rect 25280 20884 25286 20936
rect 38013 20927 38071 20933
rect 38013 20893 38025 20927
rect 38059 20924 38071 20927
rect 38378 20924 38384 20936
rect 38059 20896 38384 20924
rect 38059 20893 38071 20896
rect 38013 20887 38071 20893
rect 38378 20884 38384 20896
rect 38436 20884 38442 20936
rect 14642 20856 14648 20868
rect 12676 20828 13216 20856
rect 14603 20828 14648 20856
rect 12676 20816 12682 20828
rect 14642 20816 14648 20828
rect 14700 20816 14706 20868
rect 14734 20816 14740 20868
rect 14792 20856 14798 20868
rect 15657 20859 15715 20865
rect 14792 20828 14837 20856
rect 14792 20816 14798 20828
rect 15657 20825 15669 20859
rect 15703 20856 15715 20859
rect 15930 20856 15936 20868
rect 15703 20828 15936 20856
rect 15703 20825 15715 20828
rect 15657 20819 15715 20825
rect 15930 20816 15936 20828
rect 15988 20816 15994 20868
rect 16669 20859 16727 20865
rect 16669 20825 16681 20859
rect 16715 20825 16727 20859
rect 16669 20819 16727 20825
rect 10744 20760 12572 20788
rect 10744 20748 10750 20760
rect 16574 20748 16580 20800
rect 16632 20788 16638 20800
rect 16684 20788 16712 20819
rect 17770 20816 17776 20868
rect 17828 20856 17834 20868
rect 18233 20859 18291 20865
rect 18233 20856 18245 20859
rect 17828 20828 18245 20856
rect 17828 20816 17834 20828
rect 18233 20825 18245 20828
rect 18279 20825 18291 20859
rect 18233 20819 18291 20825
rect 18322 20816 18328 20868
rect 18380 20856 18386 20868
rect 18380 20828 18425 20856
rect 18380 20816 18386 20828
rect 20438 20816 20444 20868
rect 20496 20856 20502 20868
rect 22480 20856 22508 20884
rect 22922 20856 22928 20868
rect 20496 20828 20541 20856
rect 22480 20828 22928 20856
rect 20496 20816 20502 20828
rect 22922 20816 22928 20828
rect 22980 20816 22986 20868
rect 23293 20859 23351 20865
rect 23293 20856 23305 20859
rect 23032 20828 23305 20856
rect 16632 20760 16712 20788
rect 16632 20748 16638 20760
rect 17678 20748 17684 20800
rect 17736 20788 17742 20800
rect 23032 20788 23060 20828
rect 23293 20825 23305 20828
rect 23339 20825 23351 20859
rect 23293 20819 23351 20825
rect 25038 20788 25044 20800
rect 17736 20760 23060 20788
rect 24999 20760 25044 20788
rect 17736 20748 17742 20760
rect 25038 20748 25044 20760
rect 25096 20748 25102 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 6730 20544 6736 20596
rect 6788 20584 6794 20596
rect 7745 20587 7803 20593
rect 7745 20584 7757 20587
rect 6788 20556 7757 20584
rect 6788 20544 6794 20556
rect 7745 20553 7757 20556
rect 7791 20553 7803 20587
rect 7745 20547 7803 20553
rect 7926 20544 7932 20596
rect 7984 20584 7990 20596
rect 8846 20584 8852 20596
rect 7984 20556 8852 20584
rect 7984 20544 7990 20556
rect 8846 20544 8852 20556
rect 8904 20544 8910 20596
rect 10226 20544 10232 20596
rect 10284 20544 10290 20596
rect 12250 20544 12256 20596
rect 12308 20584 12314 20596
rect 14090 20584 14096 20596
rect 12308 20556 14096 20584
rect 12308 20544 12314 20556
rect 14090 20544 14096 20556
rect 14148 20544 14154 20596
rect 14369 20587 14427 20593
rect 14369 20553 14381 20587
rect 14415 20584 14427 20587
rect 14734 20584 14740 20596
rect 14415 20556 14740 20584
rect 14415 20553 14427 20556
rect 14369 20547 14427 20553
rect 14734 20544 14740 20556
rect 14792 20544 14798 20596
rect 16850 20584 16856 20596
rect 15212 20556 16856 20584
rect 1854 20476 1860 20528
rect 1912 20516 1918 20528
rect 1912 20488 2774 20516
rect 1912 20476 1918 20488
rect 2746 20244 2774 20488
rect 8110 20476 8116 20528
rect 8168 20516 8174 20528
rect 8389 20519 8447 20525
rect 8389 20516 8401 20519
rect 8168 20488 8401 20516
rect 8168 20476 8174 20488
rect 8389 20485 8401 20488
rect 8435 20485 8447 20519
rect 8389 20479 8447 20485
rect 8481 20519 8539 20525
rect 8481 20485 8493 20519
rect 8527 20516 8539 20519
rect 9214 20516 9220 20528
rect 8527 20488 9220 20516
rect 8527 20485 8539 20488
rect 8481 20479 8539 20485
rect 9214 20476 9220 20488
rect 9272 20476 9278 20528
rect 10244 20516 10272 20544
rect 10321 20519 10379 20525
rect 10321 20516 10333 20519
rect 10244 20488 10333 20516
rect 10321 20485 10333 20488
rect 10367 20485 10379 20519
rect 10321 20479 10379 20485
rect 10413 20519 10471 20525
rect 10413 20485 10425 20519
rect 10459 20516 10471 20519
rect 10778 20516 10784 20528
rect 10459 20488 10784 20516
rect 10459 20485 10471 20488
rect 10413 20479 10471 20485
rect 10778 20476 10784 20488
rect 10836 20476 10842 20528
rect 10962 20476 10968 20528
rect 11020 20516 11026 20528
rect 11885 20519 11943 20525
rect 11885 20516 11897 20519
rect 11020 20488 11897 20516
rect 11020 20476 11026 20488
rect 11885 20485 11897 20488
rect 11931 20485 11943 20519
rect 13262 20516 13268 20528
rect 13223 20488 13268 20516
rect 11885 20479 11943 20485
rect 13262 20476 13268 20488
rect 13320 20476 13326 20528
rect 15212 20516 15240 20556
rect 16850 20544 16856 20556
rect 16908 20544 16914 20596
rect 19242 20584 19248 20596
rect 17052 20556 19248 20584
rect 14292 20488 15240 20516
rect 14292 20460 14320 20488
rect 15286 20476 15292 20528
rect 15344 20516 15350 20528
rect 15381 20519 15439 20525
rect 15381 20516 15393 20519
rect 15344 20488 15393 20516
rect 15344 20476 15350 20488
rect 15381 20485 15393 20488
rect 15427 20485 15439 20519
rect 15381 20479 15439 20485
rect 15930 20476 15936 20528
rect 15988 20516 15994 20528
rect 16574 20516 16580 20528
rect 15988 20488 16580 20516
rect 15988 20476 15994 20488
rect 16574 20476 16580 20488
rect 16632 20476 16638 20528
rect 7650 20448 7656 20460
rect 7611 20420 7656 20448
rect 7650 20408 7656 20420
rect 7708 20408 7714 20460
rect 14274 20448 14280 20460
rect 14235 20420 14280 20448
rect 14274 20408 14280 20420
rect 14332 20408 14338 20460
rect 9214 20380 9220 20392
rect 9175 20352 9220 20380
rect 9214 20340 9220 20352
rect 9272 20380 9278 20392
rect 9582 20380 9588 20392
rect 9272 20352 9588 20380
rect 9272 20340 9278 20352
rect 9582 20340 9588 20352
rect 9640 20340 9646 20392
rect 10965 20383 11023 20389
rect 10965 20349 10977 20383
rect 11011 20380 11023 20383
rect 11514 20380 11520 20392
rect 11011 20352 11520 20380
rect 11011 20349 11023 20352
rect 10965 20343 11023 20349
rect 11514 20340 11520 20352
rect 11572 20340 11578 20392
rect 11790 20380 11796 20392
rect 11751 20352 11796 20380
rect 11790 20340 11796 20352
rect 11848 20340 11854 20392
rect 12069 20383 12127 20389
rect 12069 20349 12081 20383
rect 12115 20349 12127 20383
rect 13170 20380 13176 20392
rect 13131 20352 13176 20380
rect 12069 20343 12127 20349
rect 7098 20272 7104 20324
rect 7156 20312 7162 20324
rect 12084 20312 12112 20343
rect 13170 20340 13176 20352
rect 13228 20340 13234 20392
rect 13446 20380 13452 20392
rect 13407 20352 13452 20380
rect 13446 20340 13452 20352
rect 13504 20340 13510 20392
rect 13814 20340 13820 20392
rect 13872 20380 13878 20392
rect 15289 20383 15347 20389
rect 13872 20352 15148 20380
rect 13872 20340 13878 20352
rect 7156 20284 12112 20312
rect 15120 20312 15148 20352
rect 15289 20349 15301 20383
rect 15335 20380 15347 20383
rect 15470 20380 15476 20392
rect 15335 20352 15476 20380
rect 15335 20349 15347 20352
rect 15289 20343 15347 20349
rect 15470 20340 15476 20352
rect 15528 20340 15534 20392
rect 16301 20383 16359 20389
rect 16301 20349 16313 20383
rect 16347 20380 16359 20383
rect 17052 20380 17080 20556
rect 19242 20544 19248 20556
rect 19300 20544 19306 20596
rect 25130 20584 25136 20596
rect 19352 20556 25136 20584
rect 19352 20528 19380 20556
rect 25130 20544 25136 20556
rect 25188 20544 25194 20596
rect 26421 20587 26479 20593
rect 26421 20553 26433 20587
rect 26467 20584 26479 20587
rect 26970 20584 26976 20596
rect 26467 20556 26976 20584
rect 26467 20553 26479 20556
rect 26421 20547 26479 20553
rect 26970 20544 26976 20556
rect 27028 20544 27034 20596
rect 17310 20516 17316 20528
rect 17271 20488 17316 20516
rect 17310 20476 17316 20488
rect 17368 20476 17374 20528
rect 18138 20476 18144 20528
rect 18196 20516 18202 20528
rect 18417 20519 18475 20525
rect 18417 20516 18429 20519
rect 18196 20488 18429 20516
rect 18196 20476 18202 20488
rect 18417 20485 18429 20488
rect 18463 20485 18475 20519
rect 19334 20516 19340 20528
rect 19247 20488 19340 20516
rect 18417 20479 18475 20485
rect 19334 20476 19340 20488
rect 19392 20476 19398 20528
rect 19429 20519 19487 20525
rect 19429 20485 19441 20519
rect 19475 20516 19487 20519
rect 19886 20516 19892 20528
rect 19475 20488 19892 20516
rect 19475 20485 19487 20488
rect 19429 20479 19487 20485
rect 19886 20476 19892 20488
rect 19944 20476 19950 20528
rect 21358 20476 21364 20528
rect 21416 20516 21422 20528
rect 22189 20519 22247 20525
rect 22189 20516 22201 20519
rect 21416 20488 22201 20516
rect 21416 20476 21422 20488
rect 22189 20485 22201 20488
rect 22235 20485 22247 20519
rect 22189 20479 22247 20485
rect 23014 20476 23020 20528
rect 23072 20516 23078 20528
rect 23385 20519 23443 20525
rect 23385 20516 23397 20519
rect 23072 20488 23397 20516
rect 23072 20476 23078 20488
rect 23385 20485 23397 20488
rect 23431 20485 23443 20519
rect 23385 20479 23443 20485
rect 18325 20451 18383 20457
rect 18325 20417 18337 20451
rect 18371 20417 18383 20451
rect 24394 20448 24400 20460
rect 24355 20420 24400 20448
rect 18325 20411 18383 20417
rect 16347 20352 17080 20380
rect 17221 20383 17279 20389
rect 16347 20349 16359 20352
rect 16301 20343 16359 20349
rect 17221 20349 17233 20383
rect 17267 20380 17279 20383
rect 17586 20380 17592 20392
rect 17267 20352 17592 20380
rect 17267 20349 17279 20352
rect 17221 20343 17279 20349
rect 16316 20312 16344 20343
rect 17586 20340 17592 20352
rect 17644 20340 17650 20392
rect 18340 20380 18368 20411
rect 24394 20408 24400 20420
rect 24452 20408 24458 20460
rect 24581 20451 24639 20457
rect 24581 20417 24593 20451
rect 24627 20448 24639 20451
rect 25038 20448 25044 20460
rect 24627 20420 25044 20448
rect 24627 20417 24639 20420
rect 24581 20411 24639 20417
rect 25038 20408 25044 20420
rect 25096 20408 25102 20460
rect 25774 20448 25780 20460
rect 25735 20420 25780 20448
rect 25774 20408 25780 20420
rect 25832 20408 25838 20460
rect 27154 20448 27160 20460
rect 27115 20420 27160 20448
rect 27154 20408 27160 20420
rect 27212 20408 27218 20460
rect 38286 20448 38292 20460
rect 38247 20420 38292 20448
rect 38286 20408 38292 20420
rect 38344 20408 38350 20460
rect 19978 20380 19984 20392
rect 17696 20352 19984 20380
rect 17696 20312 17724 20352
rect 19978 20340 19984 20352
rect 20036 20340 20042 20392
rect 20162 20380 20168 20392
rect 20123 20352 20168 20380
rect 20162 20340 20168 20352
rect 20220 20340 20226 20392
rect 20990 20340 20996 20392
rect 21048 20380 21054 20392
rect 21634 20380 21640 20392
rect 21048 20352 21640 20380
rect 21048 20340 21054 20352
rect 21634 20340 21640 20352
rect 21692 20340 21698 20392
rect 22097 20383 22155 20389
rect 22097 20349 22109 20383
rect 22143 20349 22155 20383
rect 22097 20343 22155 20349
rect 15120 20284 16344 20312
rect 17052 20284 17724 20312
rect 7156 20272 7162 20284
rect 17052 20244 17080 20284
rect 17770 20272 17776 20324
rect 17828 20312 17834 20324
rect 17828 20284 17873 20312
rect 17828 20272 17834 20284
rect 18138 20272 18144 20324
rect 18196 20312 18202 20324
rect 22112 20312 22140 20343
rect 22554 20340 22560 20392
rect 22612 20380 22618 20392
rect 23290 20380 23296 20392
rect 22612 20352 23296 20380
rect 22612 20340 22618 20352
rect 23290 20340 23296 20352
rect 23348 20340 23354 20392
rect 25961 20383 26019 20389
rect 25961 20349 25973 20383
rect 26007 20380 26019 20383
rect 27249 20383 27307 20389
rect 27249 20380 27261 20383
rect 26007 20352 27261 20380
rect 26007 20349 26019 20352
rect 25961 20343 26019 20349
rect 27249 20349 27261 20352
rect 27295 20349 27307 20383
rect 27249 20343 27307 20349
rect 18196 20284 22140 20312
rect 22649 20315 22707 20321
rect 18196 20272 18202 20284
rect 22649 20281 22661 20315
rect 22695 20312 22707 20315
rect 23845 20315 23903 20321
rect 23845 20312 23857 20315
rect 22695 20284 23857 20312
rect 22695 20281 22707 20284
rect 22649 20275 22707 20281
rect 23845 20281 23857 20284
rect 23891 20312 23903 20315
rect 26786 20312 26792 20324
rect 23891 20284 26792 20312
rect 23891 20281 23903 20284
rect 23845 20275 23903 20281
rect 26786 20272 26792 20284
rect 26844 20272 26850 20324
rect 2746 20216 17080 20244
rect 17126 20204 17132 20256
rect 17184 20244 17190 20256
rect 21542 20244 21548 20256
rect 17184 20216 21548 20244
rect 17184 20204 17190 20216
rect 21542 20204 21548 20216
rect 21600 20204 21606 20256
rect 25041 20247 25099 20253
rect 25041 20213 25053 20247
rect 25087 20244 25099 20247
rect 25130 20244 25136 20256
rect 25087 20216 25136 20244
rect 25087 20213 25099 20216
rect 25041 20207 25099 20213
rect 25130 20204 25136 20216
rect 25188 20204 25194 20256
rect 34698 20204 34704 20256
rect 34756 20244 34762 20256
rect 38105 20247 38163 20253
rect 38105 20244 38117 20247
rect 34756 20216 38117 20244
rect 34756 20204 34762 20216
rect 38105 20213 38117 20216
rect 38151 20213 38163 20247
rect 38105 20207 38163 20213
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 9217 20043 9275 20049
rect 9217 20009 9229 20043
rect 9263 20040 9275 20043
rect 9950 20040 9956 20052
rect 9263 20012 9956 20040
rect 9263 20009 9275 20012
rect 9217 20003 9275 20009
rect 9950 20000 9956 20012
rect 10008 20000 10014 20052
rect 10778 20040 10784 20052
rect 10739 20012 10784 20040
rect 10778 20000 10784 20012
rect 10836 20000 10842 20052
rect 11790 20000 11796 20052
rect 11848 20040 11854 20052
rect 17218 20040 17224 20052
rect 11848 20012 17224 20040
rect 11848 20000 11854 20012
rect 17218 20000 17224 20012
rect 17276 20000 17282 20052
rect 22278 20040 22284 20052
rect 19306 20012 22284 20040
rect 6917 19975 6975 19981
rect 6917 19941 6929 19975
rect 6963 19972 6975 19975
rect 7098 19972 7104 19984
rect 6963 19944 7104 19972
rect 6963 19941 6975 19944
rect 6917 19935 6975 19941
rect 7098 19932 7104 19944
rect 7156 19932 7162 19984
rect 7650 19932 7656 19984
rect 7708 19972 7714 19984
rect 11330 19972 11336 19984
rect 7708 19944 11336 19972
rect 7708 19932 7714 19944
rect 11330 19932 11336 19944
rect 11388 19932 11394 19984
rect 19306 19972 19334 20012
rect 22278 20000 22284 20012
rect 22336 20040 22342 20052
rect 23382 20040 23388 20052
rect 22336 20012 23388 20040
rect 22336 20000 22342 20012
rect 23382 20000 23388 20012
rect 23440 20000 23446 20052
rect 25222 20000 25228 20052
rect 25280 20040 25286 20052
rect 25685 20043 25743 20049
rect 25685 20040 25697 20043
rect 25280 20012 25697 20040
rect 25280 20000 25286 20012
rect 25685 20009 25697 20012
rect 25731 20009 25743 20043
rect 25685 20003 25743 20009
rect 22738 19972 22744 19984
rect 13740 19944 19334 19972
rect 19812 19944 22744 19972
rect 5261 19907 5319 19913
rect 5261 19873 5273 19907
rect 5307 19904 5319 19907
rect 6365 19907 6423 19913
rect 6365 19904 6377 19907
rect 5307 19876 6377 19904
rect 5307 19873 5319 19876
rect 5261 19867 5319 19873
rect 6365 19873 6377 19876
rect 6411 19904 6423 19907
rect 6411 19876 13584 19904
rect 6411 19873 6423 19876
rect 6365 19867 6423 19873
rect 8938 19796 8944 19848
rect 8996 19836 9002 19848
rect 9125 19839 9183 19845
rect 9125 19836 9137 19839
rect 8996 19808 9137 19836
rect 8996 19796 9002 19808
rect 9125 19805 9137 19808
rect 9171 19805 9183 19839
rect 9766 19836 9772 19848
rect 9727 19808 9772 19836
rect 9125 19799 9183 19805
rect 9766 19796 9772 19808
rect 9824 19796 9830 19848
rect 10686 19836 10692 19848
rect 10647 19808 10692 19836
rect 10686 19796 10692 19808
rect 10744 19796 10750 19848
rect 11517 19839 11575 19845
rect 11517 19805 11529 19839
rect 11563 19836 11575 19839
rect 11606 19836 11612 19848
rect 11563 19808 11612 19836
rect 11563 19805 11575 19808
rect 11517 19799 11575 19805
rect 11606 19796 11612 19808
rect 11664 19796 11670 19848
rect 13556 19836 13584 19876
rect 13740 19836 13768 19944
rect 14090 19864 14096 19916
rect 14148 19904 14154 19916
rect 14369 19907 14427 19913
rect 14369 19904 14381 19907
rect 14148 19876 14381 19904
rect 14148 19864 14154 19876
rect 14369 19873 14381 19876
rect 14415 19873 14427 19907
rect 14369 19867 14427 19873
rect 17589 19907 17647 19913
rect 17589 19873 17601 19907
rect 17635 19904 17647 19907
rect 19334 19904 19340 19916
rect 17635 19876 19340 19904
rect 17635 19873 17647 19876
rect 17589 19867 17647 19873
rect 19334 19864 19340 19876
rect 19392 19864 19398 19916
rect 13556 19808 13768 19836
rect 16209 19839 16267 19845
rect 16209 19805 16221 19839
rect 16255 19805 16267 19839
rect 16209 19799 16267 19805
rect 17037 19839 17095 19845
rect 17037 19805 17049 19839
rect 17083 19836 17095 19839
rect 17402 19836 17408 19848
rect 17083 19808 17408 19836
rect 17083 19805 17095 19808
rect 17037 19799 17095 19805
rect 3970 19728 3976 19780
rect 4028 19768 4034 19780
rect 4249 19771 4307 19777
rect 4249 19768 4261 19771
rect 4028 19740 4261 19768
rect 4028 19728 4034 19740
rect 4249 19737 4261 19740
rect 4295 19737 4307 19771
rect 4249 19731 4307 19737
rect 4341 19771 4399 19777
rect 4341 19737 4353 19771
rect 4387 19768 4399 19771
rect 5074 19768 5080 19780
rect 4387 19740 5080 19768
rect 4387 19737 4399 19740
rect 4341 19731 4399 19737
rect 5074 19728 5080 19740
rect 5132 19728 5138 19780
rect 6457 19771 6515 19777
rect 6457 19737 6469 19771
rect 6503 19737 6515 19771
rect 6457 19731 6515 19737
rect 6472 19700 6500 19731
rect 6730 19728 6736 19780
rect 6788 19768 6794 19780
rect 7561 19771 7619 19777
rect 7561 19768 7573 19771
rect 6788 19740 7573 19768
rect 6788 19728 6794 19740
rect 7561 19737 7573 19740
rect 7607 19737 7619 19771
rect 7561 19731 7619 19737
rect 7653 19771 7711 19777
rect 7653 19737 7665 19771
rect 7699 19768 7711 19771
rect 8478 19768 8484 19780
rect 7699 19740 8484 19768
rect 7699 19737 7711 19740
rect 7653 19731 7711 19737
rect 8478 19728 8484 19740
rect 8536 19728 8542 19780
rect 8570 19728 8576 19780
rect 8628 19768 8634 19780
rect 8628 19740 8673 19768
rect 8628 19728 8634 19740
rect 10134 19728 10140 19780
rect 10192 19768 10198 19780
rect 11054 19768 11060 19780
rect 10192 19740 11060 19768
rect 10192 19728 10198 19740
rect 11054 19728 11060 19740
rect 11112 19728 11118 19780
rect 12250 19728 12256 19780
rect 12308 19768 12314 19780
rect 12437 19771 12495 19777
rect 12437 19768 12449 19771
rect 12308 19740 12449 19768
rect 12308 19728 12314 19740
rect 12437 19737 12449 19740
rect 12483 19737 12495 19771
rect 12437 19731 12495 19737
rect 12526 19728 12532 19780
rect 12584 19768 12590 19780
rect 13446 19768 13452 19780
rect 12584 19740 12629 19768
rect 13407 19740 13452 19768
rect 12584 19728 12590 19740
rect 13446 19728 13452 19740
rect 13504 19728 13510 19780
rect 14458 19728 14464 19780
rect 14516 19768 14522 19780
rect 15381 19771 15439 19777
rect 14516 19740 14561 19768
rect 14516 19728 14522 19740
rect 15381 19737 15393 19771
rect 15427 19768 15439 19771
rect 16114 19768 16120 19780
rect 15427 19740 16120 19768
rect 15427 19737 15439 19740
rect 15381 19731 15439 19737
rect 16114 19728 16120 19740
rect 16172 19728 16178 19780
rect 8202 19700 8208 19712
rect 6472 19672 8208 19700
rect 8202 19660 8208 19672
rect 8260 19660 8266 19712
rect 9861 19703 9919 19709
rect 9861 19669 9873 19703
rect 9907 19700 9919 19703
rect 10042 19700 10048 19712
rect 9907 19672 10048 19700
rect 9907 19669 9919 19672
rect 9861 19663 9919 19669
rect 10042 19660 10048 19672
rect 10100 19660 10106 19712
rect 10226 19660 10232 19712
rect 10284 19700 10290 19712
rect 10962 19700 10968 19712
rect 10284 19672 10968 19700
rect 10284 19660 10290 19672
rect 10962 19660 10968 19672
rect 11020 19660 11026 19712
rect 11609 19703 11667 19709
rect 11609 19669 11621 19703
rect 11655 19700 11667 19703
rect 12894 19700 12900 19712
rect 11655 19672 12900 19700
rect 11655 19669 11667 19672
rect 11609 19663 11667 19669
rect 12894 19660 12900 19672
rect 12952 19660 12958 19712
rect 13538 19660 13544 19712
rect 13596 19700 13602 19712
rect 16224 19700 16252 19799
rect 17402 19796 17408 19808
rect 17460 19796 17466 19848
rect 19812 19845 19840 19944
rect 22738 19932 22744 19944
rect 22796 19932 22802 19984
rect 24504 19944 25084 19972
rect 19886 19864 19892 19916
rect 19944 19904 19950 19916
rect 21266 19904 21272 19916
rect 19944 19876 19989 19904
rect 21227 19876 21272 19904
rect 19944 19864 19950 19876
rect 21266 19864 21272 19876
rect 21324 19904 21330 19916
rect 22094 19904 22100 19916
rect 21324 19876 22100 19904
rect 21324 19864 21330 19876
rect 22094 19864 22100 19876
rect 22152 19864 22158 19916
rect 22278 19904 22284 19916
rect 22239 19876 22284 19904
rect 22278 19864 22284 19876
rect 22336 19864 22342 19916
rect 24504 19848 24532 19944
rect 24581 19907 24639 19913
rect 24581 19873 24593 19907
rect 24627 19904 24639 19907
rect 24946 19904 24952 19916
rect 24627 19876 24952 19904
rect 24627 19873 24639 19876
rect 24581 19867 24639 19873
rect 24946 19864 24952 19876
rect 25004 19864 25010 19916
rect 19797 19839 19855 19845
rect 19797 19805 19809 19839
rect 19843 19805 19855 19839
rect 24486 19836 24492 19848
rect 19797 19799 19855 19805
rect 22204 19808 24492 19836
rect 16301 19771 16359 19777
rect 16301 19737 16313 19771
rect 16347 19768 16359 19771
rect 16347 19740 17540 19768
rect 16347 19737 16359 19740
rect 16301 19731 16359 19737
rect 13596 19672 16252 19700
rect 16853 19703 16911 19709
rect 13596 19660 13602 19672
rect 16853 19669 16865 19703
rect 16899 19700 16911 19703
rect 17034 19700 17040 19712
rect 16899 19672 17040 19700
rect 16899 19669 16911 19672
rect 16853 19663 16911 19669
rect 17034 19660 17040 19672
rect 17092 19660 17098 19712
rect 17512 19700 17540 19740
rect 17678 19728 17684 19780
rect 17736 19768 17742 19780
rect 18598 19768 18604 19780
rect 17736 19740 17781 19768
rect 18559 19740 18604 19768
rect 17736 19728 17742 19740
rect 18598 19728 18604 19740
rect 18656 19728 18662 19780
rect 19334 19728 19340 19780
rect 19392 19768 19398 19780
rect 20162 19768 20168 19780
rect 19392 19740 20168 19768
rect 19392 19728 19398 19740
rect 20162 19728 20168 19740
rect 20220 19728 20226 19780
rect 21361 19771 21419 19777
rect 21361 19737 21373 19771
rect 21407 19737 21419 19771
rect 21361 19731 21419 19737
rect 21376 19700 21404 19731
rect 21634 19728 21640 19780
rect 21692 19768 21698 19780
rect 22204 19768 22232 19808
rect 24486 19796 24492 19808
rect 24544 19796 24550 19848
rect 24670 19796 24676 19848
rect 24728 19836 24734 19848
rect 24765 19839 24823 19845
rect 24765 19836 24777 19839
rect 24728 19808 24777 19836
rect 24728 19796 24734 19808
rect 24765 19805 24777 19808
rect 24811 19805 24823 19839
rect 25056 19836 25084 19944
rect 25130 19932 25136 19984
rect 25188 19972 25194 19984
rect 27614 19972 27620 19984
rect 25188 19944 27620 19972
rect 25188 19932 25194 19944
rect 27614 19932 27620 19944
rect 27672 19932 27678 19984
rect 25406 19864 25412 19916
rect 25464 19904 25470 19916
rect 25464 19876 27016 19904
rect 25464 19864 25470 19876
rect 25869 19839 25927 19845
rect 25869 19836 25881 19839
rect 25056 19808 25881 19836
rect 24765 19799 24823 19805
rect 25869 19805 25881 19808
rect 25915 19805 25927 19839
rect 25869 19799 25927 19805
rect 26329 19839 26387 19845
rect 26329 19805 26341 19839
rect 26375 19836 26387 19839
rect 26694 19836 26700 19848
rect 26375 19808 26700 19836
rect 26375 19805 26387 19808
rect 26329 19799 26387 19805
rect 26694 19796 26700 19808
rect 26752 19796 26758 19848
rect 26988 19845 27016 19876
rect 26973 19839 27031 19845
rect 26973 19805 26985 19839
rect 27019 19805 27031 19839
rect 26973 19799 27031 19805
rect 28626 19796 28632 19848
rect 28684 19836 28690 19848
rect 29917 19839 29975 19845
rect 29917 19836 29929 19839
rect 28684 19808 29929 19836
rect 28684 19796 28690 19808
rect 29917 19805 29929 19808
rect 29963 19805 29975 19839
rect 29917 19799 29975 19805
rect 21692 19740 22232 19768
rect 23385 19771 23443 19777
rect 21692 19728 21698 19740
rect 23385 19737 23397 19771
rect 23431 19768 23443 19771
rect 25498 19768 25504 19780
rect 23431 19740 25504 19768
rect 23431 19737 23443 19740
rect 23385 19731 23443 19737
rect 25498 19728 25504 19740
rect 25556 19768 25562 19780
rect 37826 19768 37832 19780
rect 25556 19740 37832 19768
rect 25556 19728 25562 19740
rect 37826 19728 37832 19740
rect 37884 19728 37890 19780
rect 17512 19672 21404 19700
rect 21542 19660 21548 19712
rect 21600 19700 21606 19712
rect 23477 19703 23535 19709
rect 23477 19700 23489 19703
rect 21600 19672 23489 19700
rect 21600 19660 21606 19672
rect 23477 19669 23489 19672
rect 23523 19669 23535 19703
rect 23477 19663 23535 19669
rect 25314 19660 25320 19712
rect 25372 19700 25378 19712
rect 26421 19703 26479 19709
rect 26421 19700 26433 19703
rect 25372 19672 26433 19700
rect 25372 19660 25378 19672
rect 26421 19669 26433 19672
rect 26467 19669 26479 19703
rect 26421 19663 26479 19669
rect 26510 19660 26516 19712
rect 26568 19700 26574 19712
rect 27065 19703 27123 19709
rect 27065 19700 27077 19703
rect 26568 19672 27077 19700
rect 26568 19660 26574 19672
rect 27065 19669 27077 19672
rect 27111 19669 27123 19703
rect 27065 19663 27123 19669
rect 29733 19703 29791 19709
rect 29733 19669 29745 19703
rect 29779 19700 29791 19703
rect 29914 19700 29920 19712
rect 29779 19672 29920 19700
rect 29779 19669 29791 19672
rect 29733 19663 29791 19669
rect 29914 19660 29920 19672
rect 29972 19660 29978 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 1486 19456 1492 19508
rect 1544 19496 1550 19508
rect 1765 19499 1823 19505
rect 1765 19496 1777 19499
rect 1544 19468 1777 19496
rect 1544 19456 1550 19468
rect 1765 19465 1777 19468
rect 1811 19465 1823 19499
rect 5074 19496 5080 19508
rect 5035 19468 5080 19496
rect 1765 19459 1823 19465
rect 5074 19456 5080 19468
rect 5132 19456 5138 19508
rect 6730 19456 6736 19508
rect 6788 19496 6794 19508
rect 6788 19468 7972 19496
rect 6788 19456 6794 19468
rect 6825 19431 6883 19437
rect 6825 19397 6837 19431
rect 6871 19428 6883 19431
rect 7834 19428 7840 19440
rect 6871 19400 7840 19428
rect 6871 19397 6883 19400
rect 6825 19391 6883 19397
rect 7834 19388 7840 19400
rect 7892 19388 7898 19440
rect 1854 19320 1860 19372
rect 1912 19360 1918 19372
rect 1949 19363 2007 19369
rect 1949 19360 1961 19363
rect 1912 19332 1961 19360
rect 1912 19320 1918 19332
rect 1949 19329 1961 19332
rect 1995 19329 2007 19363
rect 1949 19323 2007 19329
rect 4985 19363 5043 19369
rect 4985 19329 4997 19363
rect 5031 19360 5043 19363
rect 5031 19332 5580 19360
rect 5031 19329 5043 19332
rect 4985 19323 5043 19329
rect 5552 19292 5580 19332
rect 5626 19320 5632 19372
rect 5684 19360 5690 19372
rect 7944 19360 7972 19468
rect 8110 19456 8116 19508
rect 8168 19496 8174 19508
rect 10413 19499 10471 19505
rect 8168 19468 10364 19496
rect 8168 19456 8174 19468
rect 8386 19428 8392 19440
rect 8347 19400 8392 19428
rect 8386 19388 8392 19400
rect 8444 19388 8450 19440
rect 8570 19388 8576 19440
rect 8628 19428 8634 19440
rect 9309 19431 9367 19437
rect 9309 19428 9321 19431
rect 8628 19400 9321 19428
rect 8628 19388 8634 19400
rect 9309 19397 9321 19400
rect 9355 19428 9367 19431
rect 9398 19428 9404 19440
rect 9355 19400 9404 19428
rect 9355 19397 9367 19400
rect 9309 19391 9367 19397
rect 9398 19388 9404 19400
rect 9456 19388 9462 19440
rect 10336 19369 10364 19468
rect 10413 19465 10425 19499
rect 10459 19496 10471 19499
rect 13262 19496 13268 19508
rect 10459 19468 13268 19496
rect 10459 19465 10471 19468
rect 10413 19459 10471 19465
rect 13262 19456 13268 19468
rect 13320 19456 13326 19508
rect 14553 19499 14611 19505
rect 14553 19465 14565 19499
rect 14599 19496 14611 19499
rect 15102 19496 15108 19508
rect 14599 19468 15108 19496
rect 14599 19465 14611 19468
rect 14553 19459 14611 19465
rect 15102 19456 15108 19468
rect 15160 19456 15166 19508
rect 15286 19496 15292 19508
rect 15247 19468 15292 19496
rect 15286 19456 15292 19468
rect 15344 19456 15350 19508
rect 16025 19499 16083 19505
rect 16025 19465 16037 19499
rect 16071 19496 16083 19499
rect 16206 19496 16212 19508
rect 16071 19468 16212 19496
rect 16071 19465 16083 19468
rect 16025 19459 16083 19465
rect 16206 19456 16212 19468
rect 16264 19456 16270 19508
rect 17402 19456 17408 19508
rect 17460 19496 17466 19508
rect 17865 19499 17923 19505
rect 17865 19496 17877 19499
rect 17460 19468 17877 19496
rect 17460 19456 17466 19468
rect 17865 19465 17877 19468
rect 17911 19465 17923 19499
rect 19426 19496 19432 19508
rect 17865 19459 17923 19465
rect 17972 19468 19432 19496
rect 11057 19431 11115 19437
rect 11057 19397 11069 19431
rect 11103 19428 11115 19431
rect 12526 19428 12532 19440
rect 11103 19400 12532 19428
rect 11103 19397 11115 19400
rect 11057 19391 11115 19397
rect 12526 19388 12532 19400
rect 12584 19388 12590 19440
rect 13078 19428 13084 19440
rect 13039 19400 13084 19428
rect 13078 19388 13084 19400
rect 13136 19388 13142 19440
rect 13446 19388 13452 19440
rect 13504 19428 13510 19440
rect 14001 19431 14059 19437
rect 14001 19428 14013 19431
rect 13504 19400 14013 19428
rect 13504 19388 13510 19400
rect 14001 19397 14013 19400
rect 14047 19428 14059 19431
rect 14366 19428 14372 19440
rect 14047 19400 14372 19428
rect 14047 19397 14059 19400
rect 14001 19391 14059 19397
rect 14366 19388 14372 19400
rect 14424 19388 14430 19440
rect 16114 19388 16120 19440
rect 16172 19428 16178 19440
rect 17972 19428 18000 19468
rect 19426 19456 19432 19468
rect 19484 19456 19490 19508
rect 20257 19499 20315 19505
rect 20257 19465 20269 19499
rect 20303 19496 20315 19499
rect 23014 19496 23020 19508
rect 20303 19468 22692 19496
rect 22975 19468 23020 19496
rect 20303 19465 20315 19468
rect 20257 19459 20315 19465
rect 22554 19428 22560 19440
rect 16172 19400 18000 19428
rect 18064 19400 22560 19428
rect 16172 19388 16178 19400
rect 10321 19363 10379 19369
rect 5684 19332 5729 19360
rect 7944 19332 8156 19360
rect 5684 19320 5690 19332
rect 5810 19292 5816 19304
rect 5552 19264 5816 19292
rect 5810 19252 5816 19264
rect 5868 19252 5874 19304
rect 6733 19295 6791 19301
rect 6733 19261 6745 19295
rect 6779 19292 6791 19295
rect 6914 19292 6920 19304
rect 6779 19264 6920 19292
rect 6779 19261 6791 19264
rect 6733 19255 6791 19261
rect 6914 19252 6920 19264
rect 6972 19252 6978 19304
rect 7098 19292 7104 19304
rect 7059 19264 7104 19292
rect 7098 19252 7104 19264
rect 7156 19252 7162 19304
rect 8128 19292 8156 19332
rect 10321 19329 10333 19363
rect 10367 19329 10379 19363
rect 10321 19323 10379 19329
rect 10870 19320 10876 19372
rect 10928 19360 10934 19372
rect 10965 19363 11023 19369
rect 10965 19360 10977 19363
rect 10928 19332 10977 19360
rect 10928 19320 10934 19332
rect 10965 19329 10977 19332
rect 11011 19329 11023 19363
rect 10965 19323 11023 19329
rect 12253 19363 12311 19369
rect 12253 19329 12265 19363
rect 12299 19360 12311 19363
rect 14737 19363 14795 19369
rect 12299 19332 12434 19360
rect 12299 19329 12311 19332
rect 12253 19323 12311 19329
rect 8297 19295 8355 19301
rect 8297 19292 8309 19295
rect 8128 19264 8309 19292
rect 8297 19261 8309 19264
rect 8343 19261 8355 19295
rect 11238 19292 11244 19304
rect 8297 19255 8355 19261
rect 8404 19264 11244 19292
rect 4798 19184 4804 19236
rect 4856 19224 4862 19236
rect 8404 19224 8432 19264
rect 11238 19252 11244 19264
rect 11296 19252 11302 19304
rect 12406 19292 12434 19332
rect 14737 19329 14749 19363
rect 14783 19360 14795 19363
rect 15197 19363 15255 19369
rect 14783 19332 15148 19360
rect 14783 19329 14795 19332
rect 14737 19323 14795 19329
rect 12986 19292 12992 19304
rect 12406 19264 12848 19292
rect 12947 19264 12992 19292
rect 4856 19196 8432 19224
rect 4856 19184 4862 19196
rect 11054 19184 11060 19236
rect 11112 19224 11118 19236
rect 12066 19224 12072 19236
rect 11112 19196 12072 19224
rect 11112 19184 11118 19196
rect 12066 19184 12072 19196
rect 12124 19184 12130 19236
rect 5718 19156 5724 19168
rect 5679 19128 5724 19156
rect 5718 19116 5724 19128
rect 5776 19116 5782 19168
rect 11422 19116 11428 19168
rect 11480 19156 11486 19168
rect 11790 19156 11796 19168
rect 11480 19128 11796 19156
rect 11480 19116 11486 19128
rect 11790 19116 11796 19128
rect 11848 19116 11854 19168
rect 12250 19116 12256 19168
rect 12308 19156 12314 19168
rect 12345 19159 12403 19165
rect 12345 19156 12357 19159
rect 12308 19128 12357 19156
rect 12308 19116 12314 19128
rect 12345 19125 12357 19128
rect 12391 19125 12403 19159
rect 12820 19156 12848 19264
rect 12986 19252 12992 19264
rect 13044 19252 13050 19304
rect 15120 19292 15148 19332
rect 15197 19329 15209 19363
rect 15243 19360 15255 19363
rect 15746 19360 15752 19372
rect 15243 19332 15752 19360
rect 15243 19329 15255 19332
rect 15197 19323 15255 19329
rect 15746 19320 15752 19332
rect 15804 19320 15810 19372
rect 15930 19360 15936 19372
rect 15891 19332 15936 19360
rect 15930 19320 15936 19332
rect 15988 19320 15994 19372
rect 17221 19363 17279 19369
rect 17221 19329 17233 19363
rect 17267 19329 17279 19363
rect 17221 19323 17279 19329
rect 17313 19363 17371 19369
rect 17313 19329 17325 19363
rect 17359 19360 17371 19363
rect 17954 19360 17960 19372
rect 17359 19332 17960 19360
rect 17359 19329 17371 19332
rect 17313 19323 17371 19329
rect 16482 19292 16488 19304
rect 15120 19264 16488 19292
rect 16482 19252 16488 19264
rect 16540 19252 16546 19304
rect 17236 19292 17264 19323
rect 17954 19320 17960 19332
rect 18012 19320 18018 19372
rect 18064 19369 18092 19400
rect 22554 19388 22560 19400
rect 22612 19388 22618 19440
rect 22664 19428 22692 19468
rect 23014 19456 23020 19468
rect 23072 19456 23078 19508
rect 23661 19499 23719 19505
rect 23661 19465 23673 19499
rect 23707 19465 23719 19499
rect 24670 19496 24676 19508
rect 24631 19468 24676 19496
rect 23661 19459 23719 19465
rect 22922 19428 22928 19440
rect 22664 19400 22928 19428
rect 22922 19388 22928 19400
rect 22980 19388 22986 19440
rect 18049 19363 18107 19369
rect 18049 19329 18061 19363
rect 18095 19329 18107 19363
rect 18049 19323 18107 19329
rect 18506 19320 18512 19372
rect 18564 19360 18570 19372
rect 19613 19363 19671 19369
rect 19613 19360 19625 19363
rect 18564 19332 19625 19360
rect 18564 19320 18570 19332
rect 19613 19329 19625 19332
rect 19659 19329 19671 19363
rect 21082 19360 21088 19372
rect 19613 19323 19671 19329
rect 19720 19332 21088 19360
rect 18230 19292 18236 19304
rect 17236 19264 18236 19292
rect 18230 19252 18236 19264
rect 18288 19292 18294 19304
rect 19720 19292 19748 19332
rect 21082 19320 21088 19332
rect 21140 19320 21146 19372
rect 21269 19363 21327 19369
rect 21269 19329 21281 19363
rect 21315 19329 21327 19363
rect 21269 19323 21327 19329
rect 18288 19264 19748 19292
rect 19797 19295 19855 19301
rect 18288 19252 18294 19264
rect 19797 19261 19809 19295
rect 19843 19292 19855 19295
rect 20622 19292 20628 19304
rect 19843 19264 20628 19292
rect 19843 19261 19855 19264
rect 19797 19255 19855 19261
rect 20622 19252 20628 19264
rect 20680 19252 20686 19304
rect 21284 19292 21312 19323
rect 21358 19320 21364 19372
rect 21416 19360 21422 19372
rect 21726 19360 21732 19372
rect 21416 19332 21461 19360
rect 21560 19332 21732 19360
rect 21416 19320 21422 19332
rect 21560 19292 21588 19332
rect 21726 19320 21732 19332
rect 21784 19360 21790 19372
rect 23201 19363 23259 19369
rect 21784 19332 23152 19360
rect 21784 19320 21790 19332
rect 21284 19264 21588 19292
rect 23124 19292 23152 19332
rect 23201 19329 23213 19363
rect 23247 19360 23259 19363
rect 23676 19360 23704 19459
rect 24670 19456 24676 19468
rect 24728 19456 24734 19508
rect 25317 19499 25375 19505
rect 25317 19465 25329 19499
rect 25363 19496 25375 19499
rect 25774 19496 25780 19508
rect 25363 19468 25780 19496
rect 25363 19465 25375 19468
rect 25317 19459 25375 19465
rect 25774 19456 25780 19468
rect 25832 19456 25838 19508
rect 26513 19499 26571 19505
rect 26513 19465 26525 19499
rect 26559 19496 26571 19499
rect 26970 19496 26976 19508
rect 26559 19468 26976 19496
rect 26559 19465 26571 19468
rect 26513 19459 26571 19465
rect 26970 19456 26976 19468
rect 27028 19456 27034 19508
rect 28626 19496 28632 19508
rect 28587 19468 28632 19496
rect 28626 19456 28632 19468
rect 28684 19456 28690 19508
rect 28718 19456 28724 19508
rect 28776 19496 28782 19508
rect 29917 19499 29975 19505
rect 29917 19496 29929 19499
rect 28776 19468 29929 19496
rect 28776 19456 28782 19468
rect 29917 19465 29929 19468
rect 29963 19465 29975 19499
rect 29917 19459 29975 19465
rect 23845 19363 23903 19369
rect 23845 19360 23857 19363
rect 23247 19332 23704 19360
rect 23768 19332 23857 19360
rect 23247 19329 23259 19332
rect 23201 19323 23259 19329
rect 23768 19292 23796 19332
rect 23845 19329 23857 19332
rect 23891 19329 23903 19363
rect 23845 19323 23903 19329
rect 24486 19320 24492 19372
rect 24544 19360 24550 19372
rect 24581 19363 24639 19369
rect 24581 19360 24593 19363
rect 24544 19332 24593 19360
rect 24544 19320 24550 19332
rect 24581 19329 24593 19332
rect 24627 19329 24639 19363
rect 24581 19323 24639 19329
rect 25225 19363 25283 19369
rect 25225 19329 25237 19363
rect 25271 19360 25283 19363
rect 25498 19360 25504 19372
rect 25271 19332 25504 19360
rect 25271 19329 25283 19332
rect 25225 19323 25283 19329
rect 25498 19320 25504 19332
rect 25556 19320 25562 19372
rect 25869 19363 25927 19369
rect 25869 19329 25881 19363
rect 25915 19360 25927 19363
rect 26602 19360 26608 19372
rect 25915 19332 26608 19360
rect 25915 19329 25927 19332
rect 25869 19323 25927 19329
rect 26602 19320 26608 19332
rect 26660 19320 26666 19372
rect 27154 19320 27160 19372
rect 27212 19360 27218 19372
rect 27341 19363 27399 19369
rect 27341 19360 27353 19363
rect 27212 19332 27353 19360
rect 27212 19320 27218 19332
rect 27341 19329 27353 19332
rect 27387 19329 27399 19363
rect 27341 19323 27399 19329
rect 28813 19363 28871 19369
rect 28813 19329 28825 19363
rect 28859 19360 28871 19363
rect 28902 19360 28908 19372
rect 28859 19332 28908 19360
rect 28859 19329 28871 19332
rect 28813 19323 28871 19329
rect 28902 19320 28908 19332
rect 28960 19320 28966 19372
rect 29086 19320 29092 19372
rect 29144 19360 29150 19372
rect 29273 19363 29331 19369
rect 29273 19360 29285 19363
rect 29144 19332 29285 19360
rect 29144 19320 29150 19332
rect 29273 19329 29285 19332
rect 29319 19329 29331 19363
rect 30098 19360 30104 19372
rect 30059 19332 30104 19360
rect 29273 19323 29331 19329
rect 30098 19320 30104 19332
rect 30156 19320 30162 19372
rect 36906 19320 36912 19372
rect 36964 19360 36970 19372
rect 38013 19363 38071 19369
rect 38013 19360 38025 19363
rect 36964 19332 38025 19360
rect 36964 19320 36970 19332
rect 38013 19329 38025 19332
rect 38059 19329 38071 19363
rect 38013 19323 38071 19329
rect 26050 19292 26056 19304
rect 23124 19264 23796 19292
rect 26011 19264 26056 19292
rect 26050 19252 26056 19264
rect 26108 19252 26114 19304
rect 20438 19184 20444 19236
rect 20496 19224 20502 19236
rect 24578 19224 24584 19236
rect 20496 19196 24584 19224
rect 20496 19184 20502 19196
rect 24578 19184 24584 19196
rect 24636 19184 24642 19236
rect 14366 19156 14372 19168
rect 12820 19128 14372 19156
rect 12345 19119 12403 19125
rect 14366 19116 14372 19128
rect 14424 19116 14430 19168
rect 14550 19116 14556 19168
rect 14608 19156 14614 19168
rect 18138 19156 18144 19168
rect 14608 19128 18144 19156
rect 14608 19116 14614 19128
rect 18138 19116 18144 19128
rect 18196 19156 18202 19168
rect 18598 19156 18604 19168
rect 18196 19128 18604 19156
rect 18196 19116 18202 19128
rect 18598 19116 18604 19128
rect 18656 19116 18662 19168
rect 20530 19116 20536 19168
rect 20588 19156 20594 19168
rect 27062 19156 27068 19168
rect 20588 19128 27068 19156
rect 20588 19116 20594 19128
rect 27062 19116 27068 19128
rect 27120 19116 27126 19168
rect 27157 19159 27215 19165
rect 27157 19125 27169 19159
rect 27203 19156 27215 19159
rect 27522 19156 27528 19168
rect 27203 19128 27528 19156
rect 27203 19125 27215 19128
rect 27157 19119 27215 19125
rect 27522 19116 27528 19128
rect 27580 19116 27586 19168
rect 29362 19156 29368 19168
rect 29323 19128 29368 19156
rect 29362 19116 29368 19128
rect 29420 19116 29426 19168
rect 38194 19156 38200 19168
rect 38155 19128 38200 19156
rect 38194 19116 38200 19128
rect 38252 19116 38258 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 7834 18952 7840 18964
rect 7795 18924 7840 18952
rect 7834 18912 7840 18924
rect 7892 18912 7898 18964
rect 8202 18912 8208 18964
rect 8260 18952 8266 18964
rect 8481 18955 8539 18961
rect 8481 18952 8493 18955
rect 8260 18924 8493 18952
rect 8260 18912 8266 18924
rect 8481 18921 8493 18924
rect 8527 18921 8539 18955
rect 8481 18915 8539 18921
rect 11149 18955 11207 18961
rect 11149 18921 11161 18955
rect 11195 18952 11207 18955
rect 13078 18952 13084 18964
rect 11195 18924 13084 18952
rect 11195 18921 11207 18924
rect 11149 18915 11207 18921
rect 13078 18912 13084 18924
rect 13136 18912 13142 18964
rect 14366 18912 14372 18964
rect 14424 18952 14430 18964
rect 17126 18952 17132 18964
rect 14424 18924 17132 18952
rect 14424 18912 14430 18924
rect 17126 18912 17132 18924
rect 17184 18912 17190 18964
rect 17221 18955 17279 18961
rect 17221 18921 17233 18955
rect 17267 18952 17279 18955
rect 17678 18952 17684 18964
rect 17267 18924 17684 18952
rect 17267 18921 17279 18924
rect 17221 18915 17279 18921
rect 17678 18912 17684 18924
rect 17736 18912 17742 18964
rect 20622 18952 20628 18964
rect 20583 18924 20628 18952
rect 20622 18912 20628 18924
rect 20680 18912 20686 18964
rect 23842 18912 23848 18964
rect 23900 18952 23906 18964
rect 23900 18924 25636 18952
rect 23900 18912 23906 18924
rect 1581 18887 1639 18893
rect 1581 18853 1593 18887
rect 1627 18853 1639 18887
rect 1581 18847 1639 18853
rect 11793 18887 11851 18893
rect 11793 18853 11805 18887
rect 11839 18884 11851 18887
rect 11839 18856 12572 18884
rect 11839 18853 11851 18856
rect 11793 18847 11851 18853
rect 1596 18816 1624 18847
rect 8662 18816 8668 18828
rect 1596 18788 6500 18816
rect 1762 18748 1768 18760
rect 1723 18720 1768 18748
rect 1762 18708 1768 18720
rect 1820 18708 1826 18760
rect 5810 18748 5816 18760
rect 5771 18720 5816 18748
rect 5810 18708 5816 18720
rect 5868 18708 5874 18760
rect 6472 18757 6500 18788
rect 7116 18788 8668 18816
rect 7116 18757 7144 18788
rect 8662 18776 8668 18788
rect 8720 18776 8726 18828
rect 12066 18816 12072 18828
rect 10428 18788 12072 18816
rect 6457 18751 6515 18757
rect 6457 18717 6469 18751
rect 6503 18717 6515 18751
rect 6457 18711 6515 18717
rect 7101 18751 7159 18757
rect 7101 18717 7113 18751
rect 7147 18717 7159 18751
rect 7101 18711 7159 18717
rect 7745 18751 7803 18757
rect 7745 18717 7757 18751
rect 7791 18717 7803 18751
rect 7745 18711 7803 18717
rect 8389 18751 8447 18757
rect 8389 18717 8401 18751
rect 8435 18717 8447 18751
rect 8389 18711 8447 18717
rect 9125 18751 9183 18757
rect 9125 18717 9137 18751
rect 9171 18748 9183 18751
rect 9766 18748 9772 18760
rect 9171 18720 9772 18748
rect 9171 18717 9183 18720
rect 9125 18711 9183 18717
rect 5442 18572 5448 18624
rect 5500 18612 5506 18624
rect 5905 18615 5963 18621
rect 5905 18612 5917 18615
rect 5500 18584 5917 18612
rect 5500 18572 5506 18584
rect 5905 18581 5917 18584
rect 5951 18581 5963 18615
rect 5905 18575 5963 18581
rect 6549 18615 6607 18621
rect 6549 18581 6561 18615
rect 6595 18612 6607 18615
rect 7006 18612 7012 18624
rect 6595 18584 7012 18612
rect 6595 18581 6607 18584
rect 6549 18575 6607 18581
rect 7006 18572 7012 18584
rect 7064 18572 7070 18624
rect 7098 18572 7104 18624
rect 7156 18612 7162 18624
rect 7193 18615 7251 18621
rect 7193 18612 7205 18615
rect 7156 18584 7205 18612
rect 7156 18572 7162 18584
rect 7193 18581 7205 18584
rect 7239 18581 7251 18615
rect 7760 18612 7788 18711
rect 8404 18680 8432 18711
rect 9766 18708 9772 18720
rect 9824 18748 9830 18760
rect 10134 18748 10140 18760
rect 9824 18720 10140 18748
rect 9824 18708 9830 18720
rect 10134 18708 10140 18720
rect 10192 18708 10198 18760
rect 10428 18757 10456 18788
rect 12066 18776 12072 18788
rect 12124 18776 12130 18828
rect 12437 18819 12495 18825
rect 12437 18816 12449 18819
rect 12176 18788 12449 18816
rect 10413 18751 10471 18757
rect 10413 18717 10425 18751
rect 10459 18717 10471 18751
rect 10413 18711 10471 18717
rect 11057 18751 11115 18757
rect 11057 18717 11069 18751
rect 11103 18748 11115 18751
rect 11238 18748 11244 18760
rect 11103 18720 11244 18748
rect 11103 18717 11115 18720
rect 11057 18711 11115 18717
rect 11238 18708 11244 18720
rect 11296 18708 11302 18760
rect 11698 18748 11704 18760
rect 11659 18720 11704 18748
rect 11698 18708 11704 18720
rect 11756 18708 11762 18760
rect 11790 18708 11796 18760
rect 11848 18748 11854 18760
rect 12176 18748 12204 18788
rect 12437 18785 12449 18788
rect 12483 18785 12495 18819
rect 12544 18816 12572 18856
rect 12618 18844 12624 18896
rect 12676 18884 12682 18896
rect 12676 18856 16804 18884
rect 12676 18844 12682 18856
rect 13722 18816 13728 18828
rect 12544 18788 13728 18816
rect 12437 18779 12495 18785
rect 13722 18776 13728 18788
rect 13780 18776 13786 18828
rect 16025 18819 16083 18825
rect 16025 18785 16037 18819
rect 16071 18816 16083 18819
rect 16206 18816 16212 18828
rect 16071 18788 16212 18816
rect 16071 18785 16083 18788
rect 16025 18779 16083 18785
rect 16206 18776 16212 18788
rect 16264 18776 16270 18828
rect 16666 18816 16672 18828
rect 16627 18788 16672 18816
rect 16666 18776 16672 18788
rect 16724 18776 16730 18828
rect 16776 18816 16804 18856
rect 25608 18825 25636 18924
rect 26050 18912 26056 18964
rect 26108 18952 26114 18964
rect 27341 18955 27399 18961
rect 27341 18952 27353 18955
rect 26108 18924 27353 18952
rect 26108 18912 26114 18924
rect 27341 18921 27353 18924
rect 27387 18921 27399 18955
rect 27341 18915 27399 18921
rect 34977 18955 35035 18961
rect 34977 18921 34989 18955
rect 35023 18952 35035 18955
rect 36906 18952 36912 18964
rect 35023 18924 36912 18952
rect 35023 18921 35035 18924
rect 34977 18915 35035 18921
rect 36906 18912 36912 18924
rect 36964 18912 36970 18964
rect 25682 18844 25688 18896
rect 25740 18884 25746 18896
rect 31573 18887 31631 18893
rect 31573 18884 31585 18887
rect 25740 18856 31585 18884
rect 25740 18844 25746 18856
rect 31573 18853 31585 18856
rect 31619 18853 31631 18887
rect 38378 18884 38384 18896
rect 31573 18847 31631 18853
rect 31726 18856 38384 18884
rect 25593 18819 25651 18825
rect 16776 18788 25544 18816
rect 17126 18748 17132 18760
rect 11848 18720 12204 18748
rect 17087 18720 17132 18748
rect 11848 18708 11854 18720
rect 17126 18708 17132 18720
rect 17184 18708 17190 18760
rect 17957 18751 18015 18757
rect 17957 18717 17969 18751
rect 18003 18717 18015 18751
rect 17957 18711 18015 18717
rect 9398 18680 9404 18692
rect 8404 18652 9404 18680
rect 9398 18640 9404 18652
rect 9456 18640 9462 18692
rect 9861 18683 9919 18689
rect 9861 18649 9873 18683
rect 9907 18680 9919 18683
rect 9907 18652 12434 18680
rect 9907 18649 9919 18652
rect 9861 18643 9919 18649
rect 9030 18612 9036 18624
rect 7760 18584 9036 18612
rect 7193 18575 7251 18581
rect 9030 18572 9036 18584
rect 9088 18572 9094 18624
rect 9214 18612 9220 18624
rect 9175 18584 9220 18612
rect 9214 18572 9220 18584
rect 9272 18572 9278 18624
rect 10502 18612 10508 18624
rect 10463 18584 10508 18612
rect 10502 18572 10508 18584
rect 10560 18572 10566 18624
rect 10594 18572 10600 18624
rect 10652 18612 10658 18624
rect 11974 18612 11980 18624
rect 10652 18584 11980 18612
rect 10652 18572 10658 18584
rect 11974 18572 11980 18584
rect 12032 18572 12038 18624
rect 12406 18612 12434 18652
rect 12526 18640 12532 18692
rect 12584 18680 12590 18692
rect 13449 18683 13507 18689
rect 12584 18652 12629 18680
rect 12584 18640 12590 18652
rect 13449 18649 13461 18683
rect 13495 18680 13507 18683
rect 14550 18680 14556 18692
rect 13495 18652 14556 18680
rect 13495 18649 13507 18652
rect 13449 18643 13507 18649
rect 14550 18640 14556 18652
rect 14608 18640 14614 18692
rect 14734 18680 14740 18692
rect 14695 18652 14740 18680
rect 14734 18640 14740 18652
rect 14792 18640 14798 18692
rect 14829 18683 14887 18689
rect 14829 18649 14841 18683
rect 14875 18649 14887 18683
rect 14829 18643 14887 18649
rect 15381 18683 15439 18689
rect 15381 18649 15393 18683
rect 15427 18680 15439 18683
rect 15470 18680 15476 18692
rect 15427 18652 15476 18680
rect 15427 18649 15439 18652
rect 15381 18643 15439 18649
rect 14844 18612 14872 18643
rect 15470 18640 15476 18652
rect 15528 18640 15534 18692
rect 16114 18680 16120 18692
rect 16075 18652 16120 18680
rect 16114 18640 16120 18652
rect 16172 18640 16178 18692
rect 17972 18680 18000 18711
rect 20254 18708 20260 18760
rect 20312 18748 20318 18760
rect 20533 18751 20591 18757
rect 20533 18748 20545 18751
rect 20312 18720 20545 18748
rect 20312 18708 20318 18720
rect 20533 18717 20545 18720
rect 20579 18717 20591 18751
rect 20533 18711 20591 18717
rect 22738 18708 22744 18760
rect 22796 18748 22802 18760
rect 23845 18751 23903 18757
rect 23845 18748 23857 18751
rect 22796 18720 23857 18748
rect 22796 18708 22802 18720
rect 23845 18717 23857 18720
rect 23891 18717 23903 18751
rect 25516 18748 25544 18788
rect 25593 18785 25605 18819
rect 25639 18785 25651 18819
rect 25593 18779 25651 18785
rect 26237 18819 26295 18825
rect 26237 18785 26249 18819
rect 26283 18816 26295 18819
rect 26602 18816 26608 18828
rect 26283 18788 26608 18816
rect 26283 18785 26295 18788
rect 26237 18779 26295 18785
rect 26602 18776 26608 18788
rect 26660 18776 26666 18828
rect 27062 18776 27068 18828
rect 27120 18816 27126 18828
rect 29089 18819 29147 18825
rect 27120 18788 29040 18816
rect 27120 18776 27126 18788
rect 29012 18760 29040 18788
rect 29089 18785 29101 18819
rect 29135 18816 29147 18819
rect 29917 18819 29975 18825
rect 29917 18816 29929 18819
rect 29135 18788 29929 18816
rect 29135 18785 29147 18788
rect 29089 18779 29147 18785
rect 29917 18785 29929 18788
rect 29963 18785 29975 18819
rect 29917 18779 29975 18785
rect 27522 18748 27528 18760
rect 25516 18720 25820 18748
rect 27483 18720 27528 18748
rect 23845 18711 23903 18717
rect 24670 18680 24676 18692
rect 16408 18652 18000 18680
rect 24631 18652 24676 18680
rect 12406 18584 14872 18612
rect 14918 18572 14924 18624
rect 14976 18612 14982 18624
rect 16408 18612 16436 18652
rect 24670 18640 24676 18652
rect 24728 18640 24734 18692
rect 24765 18683 24823 18689
rect 24765 18649 24777 18683
rect 24811 18680 24823 18683
rect 25314 18680 25320 18692
rect 24811 18652 25320 18680
rect 24811 18649 24823 18652
rect 24765 18643 24823 18649
rect 25314 18640 25320 18652
rect 25372 18640 25378 18692
rect 25792 18680 25820 18720
rect 27522 18708 27528 18720
rect 27580 18708 27586 18760
rect 28994 18748 29000 18760
rect 28907 18720 29000 18748
rect 28994 18708 29000 18720
rect 29052 18708 29058 18760
rect 29733 18751 29791 18757
rect 29733 18717 29745 18751
rect 29779 18717 29791 18751
rect 29733 18711 29791 18717
rect 31481 18751 31539 18757
rect 31481 18717 31493 18751
rect 31527 18748 31539 18751
rect 31726 18748 31754 18856
rect 38378 18844 38384 18856
rect 38436 18844 38442 18896
rect 31527 18720 31754 18748
rect 33505 18751 33563 18757
rect 31527 18717 31539 18720
rect 31481 18711 31539 18717
rect 33505 18717 33517 18751
rect 33551 18748 33563 18751
rect 34698 18748 34704 18760
rect 33551 18720 34704 18748
rect 33551 18717 33563 18720
rect 33505 18711 33563 18717
rect 26329 18683 26387 18689
rect 25792 18652 26280 18680
rect 14976 18584 16436 18612
rect 14976 18572 14982 18584
rect 16482 18572 16488 18624
rect 16540 18612 16546 18624
rect 17773 18615 17831 18621
rect 17773 18612 17785 18615
rect 16540 18584 17785 18612
rect 16540 18572 16546 18584
rect 17773 18581 17785 18584
rect 17819 18581 17831 18615
rect 17773 18575 17831 18581
rect 23937 18615 23995 18621
rect 23937 18581 23949 18615
rect 23983 18612 23995 18615
rect 25958 18612 25964 18624
rect 23983 18584 25964 18612
rect 23983 18581 23995 18584
rect 23937 18575 23995 18581
rect 25958 18572 25964 18584
rect 26016 18572 26022 18624
rect 26252 18612 26280 18652
rect 26329 18649 26341 18683
rect 26375 18680 26387 18683
rect 26510 18680 26516 18692
rect 26375 18652 26516 18680
rect 26375 18649 26387 18652
rect 26329 18643 26387 18649
rect 26510 18640 26516 18652
rect 26568 18640 26574 18692
rect 26878 18680 26884 18692
rect 26791 18652 26884 18680
rect 26878 18640 26884 18652
rect 26936 18640 26942 18692
rect 26970 18640 26976 18692
rect 27028 18680 27034 18692
rect 29748 18680 29776 18711
rect 34698 18708 34704 18720
rect 34756 18708 34762 18760
rect 35158 18748 35164 18760
rect 35119 18720 35164 18748
rect 35158 18708 35164 18720
rect 35216 18708 35222 18760
rect 27028 18652 29776 18680
rect 27028 18640 27034 18652
rect 26896 18612 26924 18640
rect 26252 18584 26924 18612
rect 30190 18572 30196 18624
rect 30248 18612 30254 18624
rect 30377 18615 30435 18621
rect 30377 18612 30389 18615
rect 30248 18584 30389 18612
rect 30248 18572 30254 18584
rect 30377 18581 30389 18584
rect 30423 18581 30435 18615
rect 33594 18612 33600 18624
rect 33555 18584 33600 18612
rect 30377 18575 30435 18581
rect 33594 18572 33600 18584
rect 33652 18572 33658 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 8754 18408 8760 18420
rect 1872 18380 8760 18408
rect 1872 18281 1900 18380
rect 8754 18368 8760 18380
rect 8812 18368 8818 18420
rect 11790 18408 11796 18420
rect 9048 18380 11796 18408
rect 4249 18343 4307 18349
rect 4249 18309 4261 18343
rect 4295 18340 4307 18343
rect 4614 18340 4620 18352
rect 4295 18312 4620 18340
rect 4295 18309 4307 18312
rect 4249 18303 4307 18309
rect 4614 18300 4620 18312
rect 4672 18300 4678 18352
rect 4798 18340 4804 18352
rect 4759 18312 4804 18340
rect 4798 18300 4804 18312
rect 4856 18300 4862 18352
rect 5442 18340 5448 18352
rect 5403 18312 5448 18340
rect 5442 18300 5448 18312
rect 5500 18300 5506 18352
rect 6638 18300 6644 18352
rect 6696 18340 6702 18352
rect 6917 18343 6975 18349
rect 6917 18340 6929 18343
rect 6696 18312 6929 18340
rect 6696 18300 6702 18312
rect 6917 18309 6929 18312
rect 6963 18309 6975 18343
rect 6917 18303 6975 18309
rect 7009 18343 7067 18349
rect 7009 18309 7021 18343
rect 7055 18340 7067 18343
rect 7926 18340 7932 18352
rect 7055 18312 7932 18340
rect 7055 18309 7067 18312
rect 7009 18303 7067 18309
rect 7926 18300 7932 18312
rect 7984 18300 7990 18352
rect 1857 18275 1915 18281
rect 1857 18241 1869 18275
rect 1903 18241 1915 18275
rect 1857 18235 1915 18241
rect 8389 18275 8447 18281
rect 8389 18241 8401 18275
rect 8435 18272 8447 18275
rect 8662 18272 8668 18284
rect 8435 18244 8668 18272
rect 8435 18241 8447 18244
rect 8389 18235 8447 18241
rect 8662 18232 8668 18244
rect 8720 18232 8726 18284
rect 9048 18281 9076 18380
rect 11790 18368 11796 18380
rect 11848 18368 11854 18420
rect 11974 18368 11980 18420
rect 12032 18408 12038 18420
rect 12434 18408 12440 18420
rect 12032 18380 12440 18408
rect 12032 18368 12038 18380
rect 12434 18368 12440 18380
rect 12492 18368 12498 18420
rect 13446 18368 13452 18420
rect 13504 18368 13510 18420
rect 13541 18411 13599 18417
rect 13541 18377 13553 18411
rect 13587 18408 13599 18411
rect 14458 18408 14464 18420
rect 13587 18380 14464 18408
rect 13587 18377 13599 18380
rect 13541 18371 13599 18377
rect 14458 18368 14464 18380
rect 14516 18368 14522 18420
rect 18141 18411 18199 18417
rect 14568 18380 18092 18408
rect 10502 18300 10508 18352
rect 10560 18340 10566 18352
rect 11885 18343 11943 18349
rect 11885 18340 11897 18343
rect 10560 18312 11897 18340
rect 10560 18300 10566 18312
rect 11885 18309 11897 18312
rect 11931 18309 11943 18343
rect 11885 18303 11943 18309
rect 12805 18343 12863 18349
rect 12805 18309 12817 18343
rect 12851 18340 12863 18343
rect 13464 18340 13492 18368
rect 14568 18340 14596 18380
rect 12851 18312 13492 18340
rect 14016 18312 14596 18340
rect 12851 18309 12863 18312
rect 12805 18303 12863 18309
rect 9033 18275 9091 18281
rect 9033 18241 9045 18275
rect 9079 18241 9091 18275
rect 9033 18235 9091 18241
rect 9677 18275 9735 18281
rect 9677 18241 9689 18275
rect 9723 18272 9735 18275
rect 9950 18272 9956 18284
rect 9723 18244 9956 18272
rect 9723 18241 9735 18244
rect 9677 18235 9735 18241
rect 9950 18232 9956 18244
rect 10008 18232 10014 18284
rect 10318 18272 10324 18284
rect 10279 18244 10324 18272
rect 10318 18232 10324 18244
rect 10376 18232 10382 18284
rect 10989 18275 11047 18281
rect 10989 18241 11001 18275
rect 11035 18272 11047 18275
rect 11330 18272 11336 18284
rect 11035 18244 11336 18272
rect 11035 18241 11047 18244
rect 10989 18235 11047 18241
rect 11330 18232 11336 18244
rect 11388 18232 11394 18284
rect 13449 18275 13507 18281
rect 13449 18241 13461 18275
rect 13495 18272 13507 18275
rect 14016 18272 14044 18312
rect 14642 18300 14648 18352
rect 14700 18340 14706 18352
rect 14921 18343 14979 18349
rect 14921 18340 14933 18343
rect 14700 18312 14933 18340
rect 14700 18300 14706 18312
rect 14921 18309 14933 18312
rect 14967 18309 14979 18343
rect 17034 18340 17040 18352
rect 16995 18312 17040 18340
rect 14921 18303 14979 18309
rect 17034 18300 17040 18312
rect 17092 18300 17098 18352
rect 18064 18340 18092 18380
rect 18141 18377 18153 18411
rect 18187 18408 18199 18411
rect 18322 18408 18328 18420
rect 18187 18380 18328 18408
rect 18187 18377 18199 18380
rect 18141 18371 18199 18377
rect 18322 18368 18328 18380
rect 18380 18368 18386 18420
rect 18414 18368 18420 18420
rect 18472 18408 18478 18420
rect 18785 18411 18843 18417
rect 18785 18408 18797 18411
rect 18472 18380 18797 18408
rect 18472 18368 18478 18380
rect 18785 18377 18797 18380
rect 18831 18377 18843 18411
rect 20254 18408 20260 18420
rect 18785 18371 18843 18377
rect 19306 18380 20260 18408
rect 19306 18340 19334 18380
rect 20254 18368 20260 18380
rect 20312 18368 20318 18420
rect 29549 18411 29607 18417
rect 24872 18380 29500 18408
rect 18064 18312 19334 18340
rect 19429 18343 19487 18349
rect 19429 18309 19441 18343
rect 19475 18340 19487 18343
rect 20346 18340 20352 18352
rect 19475 18312 20352 18340
rect 19475 18309 19487 18312
rect 19429 18303 19487 18309
rect 20346 18300 20352 18312
rect 20404 18340 20410 18352
rect 22370 18340 22376 18352
rect 20404 18312 22376 18340
rect 20404 18300 20410 18312
rect 22370 18300 22376 18312
rect 22428 18300 22434 18352
rect 23566 18300 23572 18352
rect 23624 18340 23630 18352
rect 24872 18349 24900 18380
rect 24673 18343 24731 18349
rect 24673 18340 24685 18343
rect 23624 18312 24685 18340
rect 23624 18300 23630 18312
rect 24673 18309 24685 18312
rect 24719 18309 24731 18343
rect 24673 18303 24731 18309
rect 24857 18343 24915 18349
rect 24857 18309 24869 18343
rect 24903 18309 24915 18343
rect 27798 18340 27804 18352
rect 27759 18312 27804 18340
rect 24857 18303 24915 18309
rect 27798 18300 27804 18312
rect 27856 18300 27862 18352
rect 27893 18343 27951 18349
rect 27893 18309 27905 18343
rect 27939 18340 27951 18343
rect 29362 18340 29368 18352
rect 27939 18312 29368 18340
rect 27939 18309 27951 18312
rect 27893 18303 27951 18309
rect 29362 18300 29368 18312
rect 29420 18300 29426 18352
rect 29472 18340 29500 18380
rect 29549 18377 29561 18411
rect 29595 18408 29607 18411
rect 30098 18408 30104 18420
rect 29595 18380 30104 18408
rect 29595 18377 29607 18380
rect 29549 18371 29607 18377
rect 30098 18368 30104 18380
rect 30156 18368 30162 18420
rect 30285 18411 30343 18417
rect 30285 18377 30297 18411
rect 30331 18408 30343 18411
rect 35158 18408 35164 18420
rect 30331 18380 35164 18408
rect 30331 18377 30343 18380
rect 30285 18371 30343 18377
rect 35158 18368 35164 18380
rect 35216 18368 35222 18420
rect 35342 18340 35348 18352
rect 29472 18312 35348 18340
rect 35342 18300 35348 18312
rect 35400 18300 35406 18352
rect 13495 18244 14044 18272
rect 14093 18275 14151 18281
rect 13495 18241 13507 18244
rect 13449 18235 13507 18241
rect 14093 18241 14105 18275
rect 14139 18272 14151 18275
rect 14182 18272 14188 18284
rect 14139 18244 14188 18272
rect 14139 18241 14151 18244
rect 14093 18235 14151 18241
rect 14182 18232 14188 18244
rect 14240 18232 14246 18284
rect 18046 18272 18052 18284
rect 18007 18244 18052 18272
rect 18046 18232 18052 18244
rect 18104 18232 18110 18284
rect 18693 18275 18751 18281
rect 18693 18241 18705 18275
rect 18739 18272 18751 18275
rect 18782 18272 18788 18284
rect 18739 18244 18788 18272
rect 18739 18241 18751 18244
rect 18693 18235 18751 18241
rect 18782 18232 18788 18244
rect 18840 18232 18846 18284
rect 20530 18272 20536 18284
rect 20491 18244 20536 18272
rect 20530 18232 20536 18244
rect 20588 18232 20594 18284
rect 20625 18275 20683 18281
rect 20625 18241 20637 18275
rect 20671 18272 20683 18275
rect 23658 18272 23664 18284
rect 20671 18244 23664 18272
rect 20671 18241 20683 18244
rect 20625 18235 20683 18241
rect 23658 18232 23664 18244
rect 23716 18232 23722 18284
rect 24762 18232 24768 18284
rect 24820 18272 24826 18284
rect 25501 18275 25559 18281
rect 25501 18272 25513 18275
rect 24820 18244 25513 18272
rect 24820 18232 24826 18244
rect 25501 18241 25513 18244
rect 25547 18241 25559 18275
rect 28902 18272 28908 18284
rect 28863 18244 28908 18272
rect 25501 18235 25559 18241
rect 28902 18232 28908 18244
rect 28960 18232 28966 18284
rect 28994 18232 29000 18284
rect 29052 18272 29058 18284
rect 29733 18275 29791 18281
rect 29733 18272 29745 18275
rect 29052 18244 29745 18272
rect 29052 18232 29058 18244
rect 29733 18241 29745 18244
rect 29779 18241 29791 18275
rect 30190 18272 30196 18284
rect 30151 18244 30196 18272
rect 29733 18235 29791 18241
rect 30190 18232 30196 18244
rect 30248 18232 30254 18284
rect 1578 18204 1584 18216
rect 1539 18176 1584 18204
rect 1578 18164 1584 18176
rect 1636 18164 1642 18216
rect 4157 18207 4215 18213
rect 4157 18173 4169 18207
rect 4203 18204 4215 18207
rect 5353 18207 5411 18213
rect 5353 18204 5365 18207
rect 4203 18176 5365 18204
rect 4203 18173 4215 18176
rect 4157 18167 4215 18173
rect 5353 18173 5365 18176
rect 5399 18204 5411 18207
rect 5718 18204 5724 18216
rect 5399 18176 5724 18204
rect 5399 18173 5411 18176
rect 5353 18167 5411 18173
rect 5718 18164 5724 18176
rect 5776 18164 5782 18216
rect 5997 18207 6055 18213
rect 5997 18173 6009 18207
rect 6043 18204 6055 18207
rect 6914 18204 6920 18216
rect 6043 18176 6920 18204
rect 6043 18173 6055 18176
rect 5997 18167 6055 18173
rect 6914 18164 6920 18176
rect 6972 18164 6978 18216
rect 7929 18207 7987 18213
rect 7929 18173 7941 18207
rect 7975 18204 7987 18207
rect 8570 18204 8576 18216
rect 7975 18176 8576 18204
rect 7975 18173 7987 18176
rect 7929 18167 7987 18173
rect 8570 18164 8576 18176
rect 8628 18164 8634 18216
rect 10413 18207 10471 18213
rect 10413 18173 10425 18207
rect 10459 18204 10471 18207
rect 10594 18204 10600 18216
rect 10459 18176 10600 18204
rect 10459 18173 10471 18176
rect 10413 18167 10471 18173
rect 10594 18164 10600 18176
rect 10652 18164 10658 18216
rect 11514 18164 11520 18216
rect 11572 18204 11578 18216
rect 11793 18207 11851 18213
rect 11793 18204 11805 18207
rect 11572 18176 11805 18204
rect 11572 18164 11578 18176
rect 11793 18173 11805 18176
rect 11839 18173 11851 18207
rect 11793 18167 11851 18173
rect 12066 18164 12072 18216
rect 12124 18204 12130 18216
rect 13170 18204 13176 18216
rect 12124 18176 13176 18204
rect 12124 18164 12130 18176
rect 13170 18164 13176 18176
rect 13228 18164 13234 18216
rect 13722 18164 13728 18216
rect 13780 18204 13786 18216
rect 14829 18207 14887 18213
rect 14829 18204 14841 18207
rect 13780 18176 14841 18204
rect 13780 18164 13786 18176
rect 14829 18173 14841 18176
rect 14875 18204 14887 18207
rect 15194 18204 15200 18216
rect 14875 18176 15200 18204
rect 14875 18173 14887 18176
rect 14829 18167 14887 18173
rect 15194 18164 15200 18176
rect 15252 18164 15258 18216
rect 15378 18204 15384 18216
rect 15339 18176 15384 18204
rect 15378 18164 15384 18176
rect 15436 18164 15442 18216
rect 15838 18164 15844 18216
rect 15896 18204 15902 18216
rect 16206 18204 16212 18216
rect 15896 18176 16212 18204
rect 15896 18164 15902 18176
rect 16206 18164 16212 18176
rect 16264 18164 16270 18216
rect 16945 18207 17003 18213
rect 16945 18173 16957 18207
rect 16991 18173 17003 18207
rect 16945 18167 17003 18173
rect 19613 18207 19671 18213
rect 19613 18173 19625 18207
rect 19659 18204 19671 18207
rect 23382 18204 23388 18216
rect 19659 18176 23388 18204
rect 19659 18173 19671 18176
rect 19613 18167 19671 18173
rect 8481 18139 8539 18145
rect 8481 18105 8493 18139
rect 8527 18136 8539 18139
rect 9674 18136 9680 18148
rect 8527 18108 9680 18136
rect 8527 18105 8539 18108
rect 8481 18099 8539 18105
rect 9674 18096 9680 18108
rect 9732 18096 9738 18148
rect 9769 18139 9827 18145
rect 9769 18105 9781 18139
rect 9815 18105 9827 18139
rect 9769 18099 9827 18105
rect 11057 18139 11115 18145
rect 11057 18105 11069 18139
rect 11103 18136 11115 18139
rect 14185 18139 14243 18145
rect 11103 18108 14136 18136
rect 11103 18105 11115 18108
rect 11057 18099 11115 18105
rect 9125 18071 9183 18077
rect 9125 18037 9137 18071
rect 9171 18068 9183 18071
rect 9582 18068 9588 18080
rect 9171 18040 9588 18068
rect 9171 18037 9183 18040
rect 9125 18031 9183 18037
rect 9582 18028 9588 18040
rect 9640 18028 9646 18080
rect 9784 18068 9812 18099
rect 12802 18068 12808 18080
rect 9784 18040 12808 18068
rect 12802 18028 12808 18040
rect 12860 18028 12866 18080
rect 14108 18068 14136 18108
rect 14185 18105 14197 18139
rect 14231 18136 14243 18139
rect 16114 18136 16120 18148
rect 14231 18108 16120 18136
rect 14231 18105 14243 18108
rect 14185 18099 14243 18105
rect 16114 18096 16120 18108
rect 16172 18096 16178 18148
rect 14642 18068 14648 18080
rect 14108 18040 14648 18068
rect 14642 18028 14648 18040
rect 14700 18028 14706 18080
rect 14734 18028 14740 18080
rect 14792 18068 14798 18080
rect 16960 18068 16988 18167
rect 23382 18164 23388 18176
rect 23440 18164 23446 18216
rect 24670 18164 24676 18216
rect 24728 18204 24734 18216
rect 25317 18207 25375 18213
rect 25317 18204 25329 18207
rect 24728 18176 25329 18204
rect 24728 18164 24734 18176
rect 25317 18173 25329 18176
rect 25363 18204 25375 18207
rect 25682 18204 25688 18216
rect 25363 18176 25688 18204
rect 25363 18173 25375 18176
rect 25317 18167 25375 18173
rect 25682 18164 25688 18176
rect 25740 18164 25746 18216
rect 28077 18207 28135 18213
rect 28077 18173 28089 18207
rect 28123 18173 28135 18207
rect 28077 18167 28135 18173
rect 17497 18139 17555 18145
rect 17497 18105 17509 18139
rect 17543 18136 17555 18139
rect 27982 18136 27988 18148
rect 17543 18108 27988 18136
rect 17543 18105 17555 18108
rect 17497 18099 17555 18105
rect 27982 18096 27988 18108
rect 28040 18136 28046 18148
rect 28092 18136 28120 18167
rect 28040 18108 28120 18136
rect 28040 18096 28046 18108
rect 14792 18040 16988 18068
rect 14792 18028 14798 18040
rect 21082 18028 21088 18080
rect 21140 18068 21146 18080
rect 25685 18071 25743 18077
rect 25685 18068 25697 18071
rect 21140 18040 25697 18068
rect 21140 18028 21146 18040
rect 25685 18037 25697 18040
rect 25731 18068 25743 18071
rect 26970 18068 26976 18080
rect 25731 18040 26976 18068
rect 25731 18037 25743 18040
rect 25685 18031 25743 18037
rect 26970 18028 26976 18040
rect 27028 18028 27034 18080
rect 28534 18028 28540 18080
rect 28592 18068 28598 18080
rect 28997 18071 29055 18077
rect 28997 18068 29009 18071
rect 28592 18040 29009 18068
rect 28592 18028 28598 18040
rect 28997 18037 29009 18040
rect 29043 18037 29055 18071
rect 28997 18031 29055 18037
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 4341 17867 4399 17873
rect 4341 17833 4353 17867
rect 4387 17864 4399 17867
rect 4614 17864 4620 17876
rect 4387 17836 4620 17864
rect 4387 17833 4399 17836
rect 4341 17827 4399 17833
rect 4614 17824 4620 17836
rect 4672 17824 4678 17876
rect 5166 17824 5172 17876
rect 5224 17864 5230 17876
rect 5224 17836 13676 17864
rect 5224 17824 5230 17836
rect 9401 17799 9459 17805
rect 9401 17765 9413 17799
rect 9447 17796 9459 17799
rect 10226 17796 10232 17808
rect 9447 17768 10232 17796
rect 9447 17765 9459 17768
rect 9401 17759 9459 17765
rect 10226 17756 10232 17768
rect 10284 17756 10290 17808
rect 10318 17756 10324 17808
rect 10376 17796 10382 17808
rect 11974 17796 11980 17808
rect 10376 17768 11980 17796
rect 10376 17756 10382 17768
rect 11974 17756 11980 17768
rect 12032 17756 12038 17808
rect 12360 17768 13584 17796
rect 1854 17688 1860 17740
rect 1912 17728 1918 17740
rect 8481 17731 8539 17737
rect 1912 17700 7788 17728
rect 1912 17688 1918 17700
rect 4246 17660 4252 17672
rect 4207 17632 4252 17660
rect 4246 17620 4252 17632
rect 4304 17620 4310 17672
rect 4893 17663 4951 17669
rect 4893 17629 4905 17663
rect 4939 17660 4951 17663
rect 5442 17660 5448 17672
rect 4939 17632 5448 17660
rect 4939 17629 4951 17632
rect 4893 17623 4951 17629
rect 5442 17620 5448 17632
rect 5500 17620 5506 17672
rect 7760 17669 7788 17700
rect 8481 17697 8493 17731
rect 8527 17728 8539 17731
rect 10778 17728 10784 17740
rect 8527 17700 10784 17728
rect 8527 17697 8539 17700
rect 8481 17691 8539 17697
rect 10778 17688 10784 17700
rect 10836 17688 10842 17740
rect 11333 17731 11391 17737
rect 11333 17697 11345 17731
rect 11379 17728 11391 17731
rect 11422 17728 11428 17740
rect 11379 17700 11428 17728
rect 11379 17697 11391 17700
rect 11333 17691 11391 17697
rect 11422 17688 11428 17700
rect 11480 17688 11486 17740
rect 12360 17737 12388 17768
rect 12345 17731 12403 17737
rect 12345 17697 12357 17731
rect 12391 17697 12403 17731
rect 12345 17691 12403 17697
rect 7745 17663 7803 17669
rect 7745 17629 7757 17663
rect 7791 17629 7803 17663
rect 7745 17623 7803 17629
rect 8389 17663 8447 17669
rect 8389 17629 8401 17663
rect 8435 17660 8447 17663
rect 8662 17660 8668 17672
rect 8435 17632 8668 17660
rect 8435 17629 8447 17632
rect 8389 17623 8447 17629
rect 8662 17620 8668 17632
rect 8720 17620 8726 17672
rect 9309 17663 9367 17669
rect 9309 17629 9321 17663
rect 9355 17629 9367 17663
rect 9309 17623 9367 17629
rect 9953 17663 10011 17669
rect 9953 17629 9965 17663
rect 9999 17660 10011 17663
rect 10318 17660 10324 17672
rect 9999 17632 10324 17660
rect 9999 17629 10011 17632
rect 9953 17623 10011 17629
rect 9324 17592 9352 17623
rect 10318 17620 10324 17632
rect 10376 17620 10382 17672
rect 10594 17660 10600 17672
rect 10555 17632 10600 17660
rect 10594 17620 10600 17632
rect 10652 17620 10658 17672
rect 12805 17663 12863 17669
rect 12805 17629 12817 17663
rect 12851 17629 12863 17663
rect 13556 17660 13584 17768
rect 13648 17728 13676 17836
rect 13722 17824 13728 17876
rect 13780 17864 13786 17876
rect 18509 17867 18567 17873
rect 13780 17836 17908 17864
rect 13780 17824 13786 17836
rect 14090 17728 14096 17740
rect 13648 17700 14096 17728
rect 14090 17688 14096 17700
rect 14148 17688 14154 17740
rect 15194 17728 15200 17740
rect 15155 17700 15200 17728
rect 15194 17688 15200 17700
rect 15252 17688 15258 17740
rect 16758 17728 16764 17740
rect 16719 17700 16764 17728
rect 16758 17688 16764 17700
rect 16816 17688 16822 17740
rect 17880 17737 17908 17836
rect 18509 17833 18521 17867
rect 18555 17864 18567 17867
rect 21082 17864 21088 17876
rect 18555 17836 21088 17864
rect 18555 17833 18567 17836
rect 18509 17827 18567 17833
rect 21082 17824 21088 17836
rect 21140 17824 21146 17876
rect 21174 17824 21180 17876
rect 21232 17864 21238 17876
rect 21269 17867 21327 17873
rect 21269 17864 21281 17867
rect 21232 17836 21281 17864
rect 21232 17824 21238 17836
rect 21269 17833 21281 17836
rect 21315 17833 21327 17867
rect 21910 17864 21916 17876
rect 21871 17836 21916 17864
rect 21269 17827 21327 17833
rect 21910 17824 21916 17836
rect 21968 17824 21974 17876
rect 21358 17796 21364 17808
rect 18156 17768 21364 17796
rect 17865 17731 17923 17737
rect 17865 17697 17877 17731
rect 17911 17697 17923 17731
rect 17865 17691 17923 17697
rect 17954 17688 17960 17740
rect 18012 17728 18018 17740
rect 18049 17731 18107 17737
rect 18049 17728 18061 17731
rect 18012 17700 18061 17728
rect 18012 17688 18018 17700
rect 18049 17697 18061 17700
rect 18095 17697 18107 17731
rect 18049 17691 18107 17697
rect 13814 17660 13820 17672
rect 13556 17632 13820 17660
rect 12805 17623 12863 17629
rect 10045 17595 10103 17601
rect 9324 17564 10003 17592
rect 4246 17484 4252 17536
rect 4304 17524 4310 17536
rect 4985 17527 5043 17533
rect 4985 17524 4997 17527
rect 4304 17496 4997 17524
rect 4304 17484 4310 17496
rect 4985 17493 4997 17496
rect 5031 17493 5043 17527
rect 4985 17487 5043 17493
rect 7837 17527 7895 17533
rect 7837 17493 7849 17527
rect 7883 17524 7895 17527
rect 9858 17524 9864 17536
rect 7883 17496 9864 17524
rect 7883 17493 7895 17496
rect 7837 17487 7895 17493
rect 9858 17484 9864 17496
rect 9916 17484 9922 17536
rect 9975 17524 10003 17564
rect 10045 17561 10057 17595
rect 10091 17592 10103 17595
rect 11425 17595 11483 17601
rect 10091 17564 11284 17592
rect 10091 17561 10103 17564
rect 10045 17555 10103 17561
rect 10502 17524 10508 17536
rect 9975 17496 10508 17524
rect 10502 17484 10508 17496
rect 10560 17484 10566 17536
rect 10686 17524 10692 17536
rect 10647 17496 10692 17524
rect 10686 17484 10692 17496
rect 10744 17484 10750 17536
rect 11256 17524 11284 17564
rect 11425 17561 11437 17595
rect 11471 17561 11483 17595
rect 11425 17555 11483 17561
rect 11440 17524 11468 17555
rect 11514 17552 11520 17604
rect 11572 17592 11578 17604
rect 12820 17592 12848 17623
rect 13814 17620 13820 17632
rect 13872 17620 13878 17672
rect 14461 17663 14519 17669
rect 14461 17629 14473 17663
rect 14507 17660 14519 17663
rect 14826 17660 14832 17672
rect 14507 17632 14832 17660
rect 14507 17629 14519 17632
rect 14461 17623 14519 17629
rect 14826 17620 14832 17632
rect 14884 17620 14890 17672
rect 11572 17564 12848 17592
rect 11572 17552 11578 17564
rect 12986 17552 12992 17604
rect 13044 17592 13050 17604
rect 13081 17595 13139 17601
rect 13081 17592 13093 17595
rect 13044 17564 13093 17592
rect 13044 17552 13050 17564
rect 13081 17561 13093 17564
rect 13127 17561 13139 17595
rect 13081 17555 13139 17561
rect 15286 17552 15292 17604
rect 15344 17592 15350 17604
rect 15838 17592 15844 17604
rect 15344 17564 15389 17592
rect 15799 17564 15844 17592
rect 15344 17552 15350 17564
rect 15838 17552 15844 17564
rect 15896 17552 15902 17604
rect 16393 17595 16451 17601
rect 16393 17561 16405 17595
rect 16439 17561 16451 17595
rect 16393 17555 16451 17561
rect 11256 17496 11468 17524
rect 14553 17527 14611 17533
rect 14553 17493 14565 17527
rect 14599 17524 14611 17527
rect 15654 17524 15660 17536
rect 14599 17496 15660 17524
rect 14599 17493 14611 17496
rect 14553 17487 14611 17493
rect 15654 17484 15660 17496
rect 15712 17484 15718 17536
rect 16408 17524 16436 17555
rect 16482 17552 16488 17604
rect 16540 17592 16546 17604
rect 16540 17564 16585 17592
rect 16540 17552 16546 17564
rect 18156 17524 18184 17768
rect 21358 17756 21364 17768
rect 21416 17756 21422 17808
rect 30558 17796 30564 17808
rect 24228 17768 30564 17796
rect 18414 17688 18420 17740
rect 18472 17728 18478 17740
rect 22462 17728 22468 17740
rect 18472 17700 22468 17728
rect 18472 17688 18478 17700
rect 22462 17688 22468 17700
rect 22520 17688 22526 17740
rect 23290 17688 23296 17740
rect 23348 17728 23354 17740
rect 24228 17728 24256 17768
rect 30558 17756 30564 17768
rect 30616 17756 30622 17808
rect 23348 17700 24256 17728
rect 25869 17731 25927 17737
rect 23348 17688 23354 17700
rect 25869 17697 25881 17731
rect 25915 17728 25927 17731
rect 27798 17728 27804 17740
rect 25915 17700 27804 17728
rect 25915 17697 25927 17700
rect 25869 17691 25927 17697
rect 27798 17688 27804 17700
rect 27856 17688 27862 17740
rect 18230 17620 18236 17672
rect 18288 17660 18294 17672
rect 20073 17663 20131 17669
rect 20073 17660 20085 17663
rect 18288 17632 20085 17660
rect 18288 17620 18294 17632
rect 20073 17629 20085 17632
rect 20119 17629 20131 17663
rect 20073 17623 20131 17629
rect 20162 17620 20168 17672
rect 20220 17620 20226 17672
rect 21177 17663 21235 17669
rect 21177 17629 21189 17663
rect 21223 17660 21235 17663
rect 21634 17660 21640 17672
rect 21223 17632 21640 17660
rect 21223 17629 21235 17632
rect 21177 17623 21235 17629
rect 21634 17620 21640 17632
rect 21692 17620 21698 17672
rect 21821 17663 21879 17669
rect 21821 17629 21833 17663
rect 21867 17629 21879 17663
rect 21821 17623 21879 17629
rect 20180 17592 20208 17620
rect 21836 17592 21864 17623
rect 27614 17620 27620 17672
rect 27672 17660 27678 17672
rect 28537 17663 28595 17669
rect 28537 17660 28549 17663
rect 27672 17632 28549 17660
rect 27672 17620 27678 17632
rect 28537 17629 28549 17632
rect 28583 17629 28595 17663
rect 28537 17623 28595 17629
rect 23842 17592 23848 17604
rect 20180 17564 21864 17592
rect 22066 17564 23848 17592
rect 16408 17496 18184 17524
rect 18874 17484 18880 17536
rect 18932 17524 18938 17536
rect 19429 17527 19487 17533
rect 19429 17524 19441 17527
rect 18932 17496 19441 17524
rect 18932 17484 18938 17496
rect 19429 17493 19441 17496
rect 19475 17493 19487 17527
rect 19429 17487 19487 17493
rect 19978 17484 19984 17536
rect 20036 17524 20042 17536
rect 20165 17527 20223 17533
rect 20165 17524 20177 17527
rect 20036 17496 20177 17524
rect 20036 17484 20042 17496
rect 20165 17493 20177 17496
rect 20211 17493 20223 17527
rect 20165 17487 20223 17493
rect 20254 17484 20260 17536
rect 20312 17524 20318 17536
rect 22066 17524 22094 17564
rect 23842 17552 23848 17564
rect 23900 17552 23906 17604
rect 25958 17552 25964 17604
rect 26016 17592 26022 17604
rect 26881 17595 26939 17601
rect 26016 17564 26061 17592
rect 26016 17552 26022 17564
rect 26881 17561 26893 17595
rect 26927 17561 26939 17595
rect 26881 17555 26939 17561
rect 20312 17496 22094 17524
rect 20312 17484 20318 17496
rect 22186 17484 22192 17536
rect 22244 17524 22250 17536
rect 22465 17527 22523 17533
rect 22465 17524 22477 17527
rect 22244 17496 22477 17524
rect 22244 17484 22250 17496
rect 22465 17493 22477 17496
rect 22511 17493 22523 17527
rect 22465 17487 22523 17493
rect 24762 17484 24768 17536
rect 24820 17524 24826 17536
rect 26896 17524 26924 17555
rect 24820 17496 26924 17524
rect 27893 17527 27951 17533
rect 24820 17484 24826 17496
rect 27893 17493 27905 17527
rect 27939 17524 27951 17527
rect 28166 17524 28172 17536
rect 27939 17496 28172 17524
rect 27939 17493 27951 17496
rect 27893 17487 27951 17493
rect 28166 17484 28172 17496
rect 28224 17484 28230 17536
rect 28629 17527 28687 17533
rect 28629 17493 28641 17527
rect 28675 17524 28687 17527
rect 31294 17524 31300 17536
rect 28675 17496 31300 17524
rect 28675 17493 28687 17496
rect 28629 17487 28687 17493
rect 31294 17484 31300 17496
rect 31352 17484 31358 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 7926 17320 7932 17332
rect 7887 17292 7932 17320
rect 7926 17280 7932 17292
rect 7984 17280 7990 17332
rect 11514 17320 11520 17332
rect 9140 17292 11520 17320
rect 4246 17252 4252 17264
rect 4207 17224 4252 17252
rect 4246 17212 4252 17224
rect 4304 17212 4310 17264
rect 5166 17252 5172 17264
rect 5127 17224 5172 17252
rect 5166 17212 5172 17224
rect 5224 17212 5230 17264
rect 6362 17212 6368 17264
rect 6420 17252 6426 17264
rect 6420 17224 7236 17252
rect 6420 17212 6426 17224
rect 1762 17184 1768 17196
rect 1723 17156 1768 17184
rect 1762 17144 1768 17156
rect 1820 17144 1826 17196
rect 7208 17193 7236 17224
rect 6549 17187 6607 17193
rect 6549 17153 6561 17187
rect 6595 17153 6607 17187
rect 6549 17147 6607 17153
rect 7193 17187 7251 17193
rect 7193 17153 7205 17187
rect 7239 17153 7251 17187
rect 7834 17184 7840 17196
rect 7795 17156 7840 17184
rect 7193 17147 7251 17153
rect 4157 17119 4215 17125
rect 4157 17085 4169 17119
rect 4203 17116 4215 17119
rect 4798 17116 4804 17128
rect 4203 17088 4804 17116
rect 4203 17085 4215 17088
rect 4157 17079 4215 17085
rect 4798 17076 4804 17088
rect 4856 17076 4862 17128
rect 1946 17008 1952 17060
rect 2004 17048 2010 17060
rect 6564 17048 6592 17147
rect 7834 17144 7840 17156
rect 7892 17144 7898 17196
rect 8294 17144 8300 17196
rect 8352 17184 8358 17196
rect 9140 17193 9168 17292
rect 11514 17280 11520 17292
rect 11572 17280 11578 17332
rect 11606 17280 11612 17332
rect 11664 17320 11670 17332
rect 15197 17323 15255 17329
rect 15197 17320 15209 17323
rect 11664 17292 15209 17320
rect 11664 17280 11670 17292
rect 15197 17289 15209 17292
rect 15243 17289 15255 17323
rect 15197 17283 15255 17289
rect 16209 17323 16267 17329
rect 16209 17289 16221 17323
rect 16255 17320 16267 17323
rect 16482 17320 16488 17332
rect 16255 17292 16488 17320
rect 16255 17289 16267 17292
rect 16209 17283 16267 17289
rect 16482 17280 16488 17292
rect 16540 17280 16546 17332
rect 20254 17320 20260 17332
rect 16960 17292 20260 17320
rect 9582 17212 9588 17264
rect 9640 17252 9646 17264
rect 10597 17255 10655 17261
rect 10597 17252 10609 17255
rect 9640 17224 10609 17252
rect 9640 17212 9646 17224
rect 10597 17221 10609 17224
rect 10643 17221 10655 17255
rect 10597 17215 10655 17221
rect 10870 17212 10876 17264
rect 10928 17252 10934 17264
rect 10928 17224 12204 17252
rect 10928 17212 10934 17224
rect 8481 17187 8539 17193
rect 8481 17184 8493 17187
rect 8352 17156 8493 17184
rect 8352 17144 8358 17156
rect 8481 17153 8493 17156
rect 8527 17153 8539 17187
rect 8481 17147 8539 17153
rect 9125 17187 9183 17193
rect 9125 17153 9137 17187
rect 9171 17153 9183 17187
rect 9766 17184 9772 17196
rect 9727 17156 9772 17184
rect 9125 17147 9183 17153
rect 9766 17144 9772 17156
rect 9824 17144 9830 17196
rect 9858 17144 9864 17196
rect 9916 17184 9922 17196
rect 10226 17184 10232 17196
rect 9916 17156 10232 17184
rect 9916 17144 9922 17156
rect 10226 17144 10232 17156
rect 10284 17144 10290 17196
rect 11422 17144 11428 17196
rect 11480 17184 11486 17196
rect 11885 17187 11943 17193
rect 11885 17184 11897 17187
rect 11480 17156 11897 17184
rect 11480 17144 11486 17156
rect 11885 17153 11897 17156
rect 11931 17153 11943 17187
rect 12176 17184 12204 17224
rect 12250 17212 12256 17264
rect 12308 17252 12314 17264
rect 13173 17255 13231 17261
rect 13173 17252 13185 17255
rect 12308 17224 13185 17252
rect 12308 17212 12314 17224
rect 13173 17221 13185 17224
rect 13219 17221 13231 17255
rect 13173 17215 13231 17221
rect 14093 17255 14151 17261
rect 14093 17221 14105 17255
rect 14139 17252 14151 17255
rect 16960 17252 16988 17292
rect 20254 17280 20260 17292
rect 20312 17280 20318 17332
rect 23290 17320 23296 17332
rect 20824 17292 23296 17320
rect 17126 17252 17132 17264
rect 14139 17224 16988 17252
rect 17087 17224 17132 17252
rect 14139 17221 14151 17224
rect 14093 17215 14151 17221
rect 17126 17212 17132 17224
rect 17184 17212 17190 17264
rect 18874 17252 18880 17264
rect 18835 17224 18880 17252
rect 18874 17212 18880 17224
rect 18932 17212 18938 17264
rect 18966 17212 18972 17264
rect 19024 17252 19030 17264
rect 19024 17224 19069 17252
rect 19024 17212 19030 17224
rect 19150 17212 19156 17264
rect 19208 17252 19214 17264
rect 20824 17261 20852 17292
rect 23290 17280 23296 17292
rect 23348 17280 23354 17332
rect 23382 17280 23388 17332
rect 23440 17320 23446 17332
rect 28813 17323 28871 17329
rect 23440 17292 24348 17320
rect 23440 17280 23446 17292
rect 20809 17255 20867 17261
rect 19208 17224 20300 17252
rect 19208 17212 19214 17224
rect 20272 17196 20300 17224
rect 20809 17221 20821 17255
rect 20855 17221 20867 17255
rect 20809 17215 20867 17221
rect 20901 17255 20959 17261
rect 20901 17221 20913 17255
rect 20947 17252 20959 17255
rect 22186 17252 22192 17264
rect 20947 17224 21496 17252
rect 22147 17224 22192 17252
rect 20947 17221 20959 17224
rect 20901 17215 20959 17221
rect 12176 17156 12434 17184
rect 11885 17147 11943 17153
rect 6641 17119 6699 17125
rect 6641 17085 6653 17119
rect 6687 17116 6699 17119
rect 10505 17119 10563 17125
rect 10505 17116 10517 17119
rect 6687 17088 10517 17116
rect 6687 17085 6699 17088
rect 6641 17079 6699 17085
rect 10505 17085 10517 17088
rect 10551 17085 10563 17119
rect 10505 17079 10563 17085
rect 10686 17076 10692 17128
rect 10744 17116 10750 17128
rect 10744 17088 11560 17116
rect 10744 17076 10750 17088
rect 2004 17020 6592 17048
rect 9217 17051 9275 17057
rect 2004 17008 2010 17020
rect 9217 17017 9229 17051
rect 9263 17048 9275 17051
rect 11054 17048 11060 17060
rect 9263 17020 10824 17048
rect 11015 17020 11060 17048
rect 9263 17017 9275 17020
rect 9217 17011 9275 17017
rect 1578 16980 1584 16992
rect 1539 16952 1584 16980
rect 1578 16940 1584 16952
rect 1636 16940 1642 16992
rect 7285 16983 7343 16989
rect 7285 16949 7297 16983
rect 7331 16980 7343 16983
rect 7650 16980 7656 16992
rect 7331 16952 7656 16980
rect 7331 16949 7343 16952
rect 7285 16943 7343 16949
rect 7650 16940 7656 16952
rect 7708 16940 7714 16992
rect 8570 16980 8576 16992
rect 8531 16952 8576 16980
rect 8570 16940 8576 16952
rect 8628 16940 8634 16992
rect 9858 16980 9864 16992
rect 9819 16952 9864 16980
rect 9858 16940 9864 16952
rect 9916 16940 9922 16992
rect 10318 16940 10324 16992
rect 10376 16980 10382 16992
rect 10686 16980 10692 16992
rect 10376 16952 10692 16980
rect 10376 16940 10382 16952
rect 10686 16940 10692 16952
rect 10744 16940 10750 16992
rect 10796 16980 10824 17020
rect 11054 17008 11060 17020
rect 11112 17008 11118 17060
rect 11532 17048 11560 17088
rect 11790 17076 11796 17128
rect 11848 17116 11854 17128
rect 12069 17119 12127 17125
rect 12069 17116 12081 17119
rect 11848 17088 12081 17116
rect 11848 17076 11854 17088
rect 12069 17085 12081 17088
rect 12115 17085 12127 17119
rect 12406 17116 12434 17156
rect 14274 17144 14280 17196
rect 14332 17184 14338 17196
rect 15105 17187 15163 17193
rect 14332 17156 15056 17184
rect 14332 17144 14338 17156
rect 13081 17119 13139 17125
rect 13081 17116 13093 17119
rect 12406 17088 13093 17116
rect 12069 17079 12127 17085
rect 13081 17085 13093 17088
rect 13127 17085 13139 17119
rect 13081 17079 13139 17085
rect 13538 17076 13544 17128
rect 13596 17116 13602 17128
rect 14918 17116 14924 17128
rect 13596 17088 14924 17116
rect 13596 17076 13602 17088
rect 14918 17076 14924 17088
rect 14976 17076 14982 17128
rect 15028 17116 15056 17156
rect 15105 17153 15117 17187
rect 15151 17184 15163 17187
rect 15930 17184 15936 17196
rect 15151 17156 15936 17184
rect 15151 17153 15163 17156
rect 15105 17147 15163 17153
rect 15930 17144 15936 17156
rect 15988 17144 15994 17196
rect 16114 17184 16120 17196
rect 16075 17156 16120 17184
rect 16114 17144 16120 17156
rect 16172 17144 16178 17196
rect 16758 17184 16764 17196
rect 16211 17156 16764 17184
rect 16211 17116 16239 17156
rect 16758 17144 16764 17156
rect 16816 17144 16822 17196
rect 19981 17187 20039 17193
rect 19981 17153 19993 17187
rect 20027 17153 20039 17187
rect 19981 17147 20039 17153
rect 15028 17088 16239 17116
rect 16666 17076 16672 17128
rect 16724 17116 16730 17128
rect 17037 17119 17095 17125
rect 17037 17116 17049 17119
rect 16724 17088 17049 17116
rect 16724 17076 16730 17088
rect 17037 17085 17049 17088
rect 17083 17085 17095 17119
rect 17037 17079 17095 17085
rect 17865 17119 17923 17125
rect 17865 17085 17877 17119
rect 17911 17116 17923 17119
rect 17954 17116 17960 17128
rect 17911 17088 17960 17116
rect 17911 17085 17923 17088
rect 17865 17079 17923 17085
rect 17954 17076 17960 17088
rect 18012 17076 18018 17128
rect 19521 17119 19579 17125
rect 19521 17085 19533 17119
rect 19567 17116 19579 17119
rect 19610 17116 19616 17128
rect 19567 17088 19616 17116
rect 19567 17085 19579 17088
rect 19521 17079 19579 17085
rect 19610 17076 19616 17088
rect 19668 17076 19674 17128
rect 19996 17116 20024 17147
rect 20254 17144 20260 17196
rect 20312 17144 20318 17196
rect 20806 17116 20812 17128
rect 19996 17088 20812 17116
rect 20806 17076 20812 17088
rect 20864 17076 20870 17128
rect 21085 17119 21143 17125
rect 21085 17085 21097 17119
rect 21131 17085 21143 17119
rect 21085 17079 21143 17085
rect 14642 17048 14648 17060
rect 11532 17020 14648 17048
rect 14642 17008 14648 17020
rect 14700 17008 14706 17060
rect 15102 17008 15108 17060
rect 15160 17048 15166 17060
rect 18230 17048 18236 17060
rect 15160 17020 18236 17048
rect 15160 17008 15166 17020
rect 18230 17008 18236 17020
rect 18288 17008 18294 17060
rect 19536 17020 20208 17048
rect 13446 16980 13452 16992
rect 10796 16952 13452 16980
rect 13446 16940 13452 16952
rect 13504 16940 13510 16992
rect 14090 16940 14096 16992
rect 14148 16980 14154 16992
rect 19536 16980 19564 17020
rect 20070 16980 20076 16992
rect 14148 16952 19564 16980
rect 20031 16952 20076 16980
rect 14148 16940 14154 16952
rect 20070 16940 20076 16952
rect 20128 16940 20134 16992
rect 20180 16980 20208 17020
rect 20530 17008 20536 17060
rect 20588 17048 20594 17060
rect 21100 17048 21128 17079
rect 20588 17020 21128 17048
rect 21468 17048 21496 17224
rect 22186 17212 22192 17224
rect 22244 17212 22250 17264
rect 22278 17212 22284 17264
rect 22336 17252 22342 17264
rect 22336 17224 22381 17252
rect 22336 17212 22342 17224
rect 22830 17212 22836 17264
rect 22888 17252 22894 17264
rect 23198 17252 23204 17264
rect 22888 17224 23204 17252
rect 22888 17212 22894 17224
rect 23198 17212 23204 17224
rect 23256 17212 23262 17264
rect 24210 17252 24216 17264
rect 24171 17224 24216 17252
rect 24210 17212 24216 17224
rect 24268 17212 24274 17264
rect 24320 17252 24348 17292
rect 28813 17289 28825 17323
rect 28859 17320 28871 17323
rect 30190 17320 30196 17332
rect 28859 17292 30196 17320
rect 28859 17289 28871 17292
rect 28813 17283 28871 17289
rect 30190 17280 30196 17292
rect 30248 17280 30254 17332
rect 37918 17252 37924 17264
rect 24320 17224 37924 17252
rect 37918 17212 37924 17224
rect 37976 17212 37982 17264
rect 28166 17184 28172 17196
rect 28127 17156 28172 17184
rect 28166 17144 28172 17156
rect 28224 17144 28230 17196
rect 28353 17187 28411 17193
rect 28353 17153 28365 17187
rect 28399 17184 28411 17187
rect 28718 17184 28724 17196
rect 28399 17156 28724 17184
rect 28399 17153 28411 17156
rect 28353 17147 28411 17153
rect 28718 17144 28724 17156
rect 28776 17144 28782 17196
rect 32582 17144 32588 17196
rect 32640 17184 32646 17196
rect 32953 17187 33011 17193
rect 32953 17184 32965 17187
rect 32640 17156 32965 17184
rect 32640 17144 32646 17156
rect 32953 17153 32965 17156
rect 32999 17153 33011 17187
rect 38013 17187 38071 17193
rect 38013 17184 38025 17187
rect 32953 17147 33011 17153
rect 35866 17156 38025 17184
rect 24121 17119 24179 17125
rect 24121 17085 24133 17119
rect 24167 17085 24179 17119
rect 24394 17116 24400 17128
rect 24355 17088 24400 17116
rect 24121 17079 24179 17085
rect 22554 17048 22560 17060
rect 21468 17020 22560 17048
rect 20588 17008 20594 17020
rect 22554 17008 22560 17020
rect 22612 17008 22618 17060
rect 24136 17048 24164 17079
rect 24394 17076 24400 17088
rect 24452 17076 24458 17128
rect 29273 17119 29331 17125
rect 29273 17085 29285 17119
rect 29319 17116 29331 17119
rect 29822 17116 29828 17128
rect 29319 17088 29828 17116
rect 29319 17085 29331 17088
rect 29273 17079 29331 17085
rect 29822 17076 29828 17088
rect 29880 17076 29886 17128
rect 24946 17048 24952 17060
rect 24136 17020 24952 17048
rect 24946 17008 24952 17020
rect 25004 17008 25010 17060
rect 32769 17051 32827 17057
rect 32769 17017 32781 17051
rect 32815 17048 32827 17051
rect 35866 17048 35894 17156
rect 38013 17153 38025 17156
rect 38059 17153 38071 17187
rect 38013 17147 38071 17153
rect 38194 17048 38200 17060
rect 32815 17020 35894 17048
rect 38155 17020 38200 17048
rect 32815 17017 32827 17020
rect 32769 17011 32827 17017
rect 38194 17008 38200 17020
rect 38252 17008 38258 17060
rect 24578 16980 24584 16992
rect 20180 16952 24584 16980
rect 24578 16940 24584 16952
rect 24636 16980 24642 16992
rect 24762 16980 24768 16992
rect 24636 16952 24768 16980
rect 24636 16940 24642 16952
rect 24762 16940 24768 16952
rect 24820 16940 24826 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 3694 16736 3700 16788
rect 3752 16776 3758 16788
rect 9674 16776 9680 16788
rect 3752 16748 9680 16776
rect 3752 16736 3758 16748
rect 9674 16736 9680 16748
rect 9732 16736 9738 16788
rect 9858 16736 9864 16788
rect 9916 16776 9922 16788
rect 14458 16776 14464 16788
rect 9916 16748 14464 16776
rect 9916 16736 9922 16748
rect 14458 16736 14464 16748
rect 14516 16736 14522 16788
rect 16022 16736 16028 16788
rect 16080 16776 16086 16788
rect 16298 16776 16304 16788
rect 16080 16748 16304 16776
rect 16080 16736 16086 16748
rect 16298 16736 16304 16748
rect 16356 16736 16362 16788
rect 17037 16779 17095 16785
rect 17037 16745 17049 16779
rect 17083 16776 17095 16779
rect 17126 16776 17132 16788
rect 17083 16748 17132 16776
rect 17083 16745 17095 16748
rect 17037 16739 17095 16745
rect 17126 16736 17132 16748
rect 17184 16736 17190 16788
rect 18601 16779 18659 16785
rect 18601 16745 18613 16779
rect 18647 16776 18659 16779
rect 18966 16776 18972 16788
rect 18647 16748 18972 16776
rect 18647 16745 18659 16748
rect 18601 16739 18659 16745
rect 18966 16736 18972 16748
rect 19024 16736 19030 16788
rect 23477 16779 23535 16785
rect 19306 16748 20392 16776
rect 6822 16668 6828 16720
rect 6880 16708 6886 16720
rect 6880 16680 7144 16708
rect 6880 16668 6886 16680
rect 1578 16600 1584 16652
rect 1636 16640 1642 16652
rect 7006 16640 7012 16652
rect 1636 16612 6316 16640
rect 6967 16612 7012 16640
rect 1636 16600 1642 16612
rect 6288 16581 6316 16612
rect 7006 16600 7012 16612
rect 7064 16600 7070 16652
rect 7116 16640 7144 16680
rect 8570 16668 8576 16720
rect 8628 16708 8634 16720
rect 14734 16708 14740 16720
rect 8628 16680 14740 16708
rect 8628 16668 8634 16680
rect 14734 16668 14740 16680
rect 14792 16668 14798 16720
rect 14918 16668 14924 16720
rect 14976 16708 14982 16720
rect 14976 16680 18644 16708
rect 14976 16668 14982 16680
rect 10229 16643 10287 16649
rect 10229 16640 10241 16643
rect 7116 16612 10241 16640
rect 10229 16609 10241 16612
rect 10275 16609 10287 16643
rect 10870 16640 10876 16652
rect 10831 16612 10876 16640
rect 10229 16603 10287 16609
rect 10870 16600 10876 16612
rect 10928 16600 10934 16652
rect 11514 16600 11520 16652
rect 11572 16640 11578 16652
rect 12066 16640 12072 16652
rect 11572 16612 12072 16640
rect 11572 16600 11578 16612
rect 12066 16600 12072 16612
rect 12124 16600 12130 16652
rect 12621 16643 12679 16649
rect 12621 16609 12633 16643
rect 12667 16640 12679 16643
rect 15562 16640 15568 16652
rect 12667 16612 15568 16640
rect 12667 16609 12679 16612
rect 12621 16603 12679 16609
rect 15562 16600 15568 16612
rect 15620 16600 15626 16652
rect 16482 16600 16488 16652
rect 16540 16640 16546 16652
rect 18616 16640 18644 16680
rect 19306 16640 19334 16748
rect 20364 16708 20392 16748
rect 23477 16745 23489 16779
rect 23523 16776 23535 16779
rect 24210 16776 24216 16788
rect 23523 16748 24216 16776
rect 23523 16745 23535 16748
rect 23477 16739 23535 16745
rect 24210 16736 24216 16748
rect 24268 16736 24274 16788
rect 24394 16708 24400 16720
rect 20364 16680 24400 16708
rect 24394 16668 24400 16680
rect 24452 16668 24458 16720
rect 28736 16680 30144 16708
rect 23106 16640 23112 16652
rect 16540 16612 18552 16640
rect 18616 16612 19334 16640
rect 21468 16612 23112 16640
rect 16540 16600 16546 16612
rect 6273 16575 6331 16581
rect 6273 16541 6285 16575
rect 6319 16541 6331 16575
rect 6273 16535 6331 16541
rect 9674 16532 9680 16584
rect 9732 16572 9738 16584
rect 10042 16572 10048 16584
rect 9732 16544 10048 16572
rect 9732 16532 9738 16544
rect 10042 16532 10048 16544
rect 10100 16532 10106 16584
rect 11422 16572 11428 16584
rect 11335 16544 11428 16572
rect 11422 16532 11428 16544
rect 11480 16572 11486 16584
rect 11606 16572 11612 16584
rect 11480 16544 11612 16572
rect 11480 16532 11486 16544
rect 11606 16532 11612 16544
rect 11664 16532 11670 16584
rect 15470 16572 15476 16584
rect 15431 16544 15476 16572
rect 15470 16532 15476 16544
rect 15528 16532 15534 16584
rect 16666 16572 16672 16584
rect 15764 16544 16672 16572
rect 7098 16464 7104 16516
rect 7156 16504 7162 16516
rect 8018 16504 8024 16516
rect 7156 16476 7201 16504
rect 7979 16476 8024 16504
rect 7156 16464 7162 16476
rect 8018 16464 8024 16476
rect 8076 16464 8082 16516
rect 9214 16464 9220 16516
rect 9272 16504 9278 16516
rect 10321 16507 10379 16513
rect 10321 16504 10333 16507
rect 9272 16476 10333 16504
rect 9272 16464 9278 16476
rect 10321 16473 10333 16476
rect 10367 16473 10379 16507
rect 10321 16467 10379 16473
rect 10594 16464 10600 16516
rect 10652 16504 10658 16516
rect 11793 16507 11851 16513
rect 11793 16504 11805 16507
rect 10652 16476 11805 16504
rect 10652 16464 10658 16476
rect 11793 16473 11805 16476
rect 11839 16504 11851 16507
rect 12618 16504 12624 16516
rect 11839 16476 12624 16504
rect 11839 16473 11851 16476
rect 11793 16467 11851 16473
rect 12618 16464 12624 16476
rect 12676 16464 12682 16516
rect 12713 16507 12771 16513
rect 12713 16473 12725 16507
rect 12759 16504 12771 16507
rect 12894 16504 12900 16516
rect 12759 16476 12900 16504
rect 12759 16473 12771 16476
rect 12713 16467 12771 16473
rect 12894 16464 12900 16476
rect 12952 16464 12958 16516
rect 13633 16507 13691 16513
rect 13633 16473 13645 16507
rect 13679 16504 13691 16507
rect 14090 16504 14096 16516
rect 13679 16476 14096 16504
rect 13679 16473 13691 16476
rect 13633 16467 13691 16473
rect 14090 16464 14096 16476
rect 14148 16464 14154 16516
rect 14369 16507 14427 16513
rect 14369 16473 14381 16507
rect 14415 16473 14427 16507
rect 14369 16467 14427 16473
rect 6365 16439 6423 16445
rect 6365 16405 6377 16439
rect 6411 16436 6423 16439
rect 8478 16436 8484 16448
rect 6411 16408 8484 16436
rect 6411 16405 6423 16408
rect 6365 16399 6423 16405
rect 8478 16396 8484 16408
rect 8536 16396 8542 16448
rect 9493 16439 9551 16445
rect 9493 16405 9505 16439
rect 9539 16436 9551 16439
rect 14384 16436 14412 16467
rect 14458 16464 14464 16516
rect 14516 16504 14522 16516
rect 14516 16476 14561 16504
rect 14516 16464 14522 16476
rect 15286 16464 15292 16516
rect 15344 16504 15350 16516
rect 15764 16513 15792 16544
rect 16666 16532 16672 16544
rect 16724 16532 16730 16584
rect 16758 16532 16764 16584
rect 16816 16572 16822 16584
rect 16945 16575 17003 16581
rect 16945 16572 16957 16575
rect 16816 16544 16957 16572
rect 16816 16532 16822 16544
rect 16945 16541 16957 16544
rect 16991 16541 17003 16575
rect 16945 16535 17003 16541
rect 17589 16575 17647 16581
rect 17589 16541 17601 16575
rect 17635 16572 17647 16575
rect 17678 16572 17684 16584
rect 17635 16544 17684 16572
rect 17635 16541 17647 16544
rect 17589 16535 17647 16541
rect 17678 16532 17684 16544
rect 17736 16532 17742 16584
rect 18524 16581 18552 16612
rect 18509 16575 18567 16581
rect 18509 16541 18521 16575
rect 18555 16541 18567 16575
rect 18509 16535 18567 16541
rect 20165 16575 20223 16581
rect 20165 16541 20177 16575
rect 20211 16572 20223 16575
rect 20714 16572 20720 16584
rect 20211 16544 20720 16572
rect 20211 16541 20223 16544
rect 20165 16535 20223 16541
rect 20714 16532 20720 16544
rect 20772 16572 20778 16584
rect 21468 16572 21496 16612
rect 23106 16600 23112 16612
rect 23164 16600 23170 16652
rect 23492 16612 24624 16640
rect 20772 16544 21496 16572
rect 21729 16575 21787 16581
rect 20772 16532 20778 16544
rect 21729 16541 21741 16575
rect 21775 16541 21787 16575
rect 22462 16572 22468 16584
rect 22375 16544 22468 16572
rect 21729 16535 21787 16541
rect 15749 16507 15807 16513
rect 15749 16504 15761 16507
rect 15344 16476 15761 16504
rect 15344 16464 15350 16476
rect 15749 16473 15761 16476
rect 15795 16473 15807 16507
rect 15749 16467 15807 16473
rect 15930 16464 15936 16516
rect 15988 16504 15994 16516
rect 19518 16504 19524 16516
rect 15988 16476 17816 16504
rect 19479 16476 19524 16504
rect 15988 16464 15994 16476
rect 9539 16408 14412 16436
rect 9539 16405 9551 16408
rect 9493 16399 9551 16405
rect 14550 16396 14556 16448
rect 14608 16436 14614 16448
rect 17681 16439 17739 16445
rect 17681 16436 17693 16439
rect 14608 16408 17693 16436
rect 14608 16396 14614 16408
rect 17681 16405 17693 16408
rect 17727 16405 17739 16439
rect 17788 16436 17816 16476
rect 19518 16464 19524 16476
rect 19576 16464 19582 16516
rect 19613 16507 19671 16513
rect 19613 16473 19625 16507
rect 19659 16504 19671 16507
rect 19978 16504 19984 16516
rect 19659 16476 19984 16504
rect 19659 16473 19671 16476
rect 19613 16467 19671 16473
rect 19978 16464 19984 16476
rect 20036 16464 20042 16516
rect 20254 16464 20260 16516
rect 20312 16504 20318 16516
rect 21744 16504 21772 16535
rect 22462 16532 22468 16544
rect 22520 16532 22526 16584
rect 22554 16532 22560 16584
rect 22612 16572 22618 16584
rect 23382 16572 23388 16584
rect 22612 16544 22657 16572
rect 23343 16544 23388 16572
rect 22612 16532 22618 16544
rect 23382 16532 23388 16544
rect 23440 16532 23446 16584
rect 20312 16476 21772 16504
rect 21821 16507 21879 16513
rect 20312 16464 20318 16476
rect 21821 16473 21833 16507
rect 21867 16504 21879 16507
rect 22278 16504 22284 16516
rect 21867 16476 22284 16504
rect 21867 16473 21879 16476
rect 21821 16467 21879 16473
rect 22278 16464 22284 16476
rect 22336 16464 22342 16516
rect 22480 16504 22508 16532
rect 23492 16504 23520 16612
rect 24596 16581 24624 16612
rect 27430 16600 27436 16652
rect 27488 16640 27494 16652
rect 28736 16649 28764 16680
rect 28721 16643 28779 16649
rect 28721 16640 28733 16643
rect 27488 16612 28733 16640
rect 27488 16600 27494 16612
rect 28721 16609 28733 16612
rect 28767 16609 28779 16643
rect 29822 16640 29828 16652
rect 29783 16612 29828 16640
rect 28721 16603 28779 16609
rect 29822 16600 29828 16612
rect 29880 16600 29886 16652
rect 30116 16649 30144 16680
rect 30101 16643 30159 16649
rect 30101 16609 30113 16643
rect 30147 16609 30159 16643
rect 30101 16603 30159 16609
rect 24581 16575 24639 16581
rect 24581 16541 24593 16575
rect 24627 16541 24639 16575
rect 24581 16535 24639 16541
rect 26326 16532 26332 16584
rect 26384 16572 26390 16584
rect 27525 16575 27583 16581
rect 27525 16572 27537 16575
rect 26384 16544 27537 16572
rect 26384 16532 26390 16544
rect 27525 16541 27537 16544
rect 27571 16541 27583 16575
rect 27525 16535 27583 16541
rect 22480 16476 23520 16504
rect 28166 16464 28172 16516
rect 28224 16504 28230 16516
rect 28445 16507 28503 16513
rect 28445 16504 28457 16507
rect 28224 16476 28457 16504
rect 28224 16464 28230 16476
rect 28445 16473 28457 16476
rect 28491 16473 28503 16507
rect 28445 16467 28503 16473
rect 28534 16464 28540 16516
rect 28592 16504 28598 16516
rect 29914 16504 29920 16516
rect 28592 16476 28637 16504
rect 29875 16476 29920 16504
rect 28592 16464 28598 16476
rect 29914 16464 29920 16476
rect 29972 16464 29978 16516
rect 21082 16436 21088 16448
rect 17788 16408 21088 16436
rect 17681 16399 17739 16405
rect 21082 16396 21088 16408
rect 21140 16396 21146 16448
rect 24486 16396 24492 16448
rect 24544 16436 24550 16448
rect 24673 16439 24731 16445
rect 24673 16436 24685 16439
rect 24544 16408 24685 16436
rect 24544 16396 24550 16408
rect 24673 16405 24685 16408
rect 24719 16405 24731 16439
rect 24673 16399 24731 16405
rect 27341 16439 27399 16445
rect 27341 16405 27353 16439
rect 27387 16436 27399 16439
rect 38010 16436 38016 16448
rect 27387 16408 38016 16436
rect 27387 16405 27399 16408
rect 27341 16399 27399 16405
rect 38010 16396 38016 16408
rect 38068 16396 38074 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 3881 16235 3939 16241
rect 3881 16232 3893 16235
rect 2746 16204 3893 16232
rect 2746 16164 2774 16204
rect 3881 16201 3893 16204
rect 3927 16201 3939 16235
rect 3881 16195 3939 16201
rect 5169 16235 5227 16241
rect 5169 16201 5181 16235
rect 5215 16232 5227 16235
rect 7558 16232 7564 16244
rect 5215 16204 7564 16232
rect 5215 16201 5227 16204
rect 5169 16195 5227 16201
rect 7558 16192 7564 16204
rect 7616 16192 7622 16244
rect 8496 16204 9720 16232
rect 8496 16176 8524 16204
rect 1596 16136 2774 16164
rect 1596 16105 1624 16136
rect 7374 16124 7380 16176
rect 7432 16164 7438 16176
rect 8202 16164 8208 16176
rect 7432 16136 8208 16164
rect 7432 16124 7438 16136
rect 8202 16124 8208 16136
rect 8260 16124 8266 16176
rect 8478 16164 8484 16176
rect 8439 16136 8484 16164
rect 8478 16124 8484 16136
rect 8536 16124 8542 16176
rect 8573 16167 8631 16173
rect 8573 16133 8585 16167
rect 8619 16164 8631 16167
rect 9490 16164 9496 16176
rect 8619 16136 9496 16164
rect 8619 16133 8631 16136
rect 8573 16127 8631 16133
rect 9490 16124 9496 16136
rect 9548 16124 9554 16176
rect 9692 16173 9720 16204
rect 16114 16192 16120 16244
rect 16172 16232 16178 16244
rect 16172 16204 19288 16232
rect 16172 16192 16178 16204
rect 9677 16167 9735 16173
rect 9677 16133 9689 16167
rect 9723 16133 9735 16167
rect 9677 16127 9735 16133
rect 9766 16124 9772 16176
rect 9824 16164 9830 16176
rect 9824 16136 9869 16164
rect 9824 16124 9830 16136
rect 10778 16124 10784 16176
rect 10836 16164 10842 16176
rect 12253 16167 12311 16173
rect 12253 16164 12265 16167
rect 10836 16136 12265 16164
rect 10836 16124 10842 16136
rect 12253 16133 12265 16136
rect 12299 16133 12311 16167
rect 13446 16164 13452 16176
rect 13407 16136 13452 16164
rect 12253 16127 12311 16133
rect 13446 16124 13452 16136
rect 13504 16124 13510 16176
rect 14366 16164 14372 16176
rect 14279 16136 14372 16164
rect 14366 16124 14372 16136
rect 14424 16164 14430 16176
rect 15010 16164 15016 16176
rect 14424 16136 15016 16164
rect 14424 16124 14430 16136
rect 15010 16124 15016 16136
rect 15068 16124 15074 16176
rect 15654 16164 15660 16176
rect 15615 16136 15660 16164
rect 15654 16124 15660 16136
rect 15712 16124 15718 16176
rect 16666 16124 16672 16176
rect 16724 16164 16730 16176
rect 18506 16164 18512 16176
rect 16724 16136 17724 16164
rect 18467 16136 18512 16164
rect 16724 16124 16730 16136
rect 1581 16099 1639 16105
rect 1581 16065 1593 16099
rect 1627 16065 1639 16099
rect 2498 16096 2504 16108
rect 2459 16068 2504 16096
rect 1581 16059 1639 16065
rect 2498 16056 2504 16068
rect 2556 16056 2562 16108
rect 4062 16096 4068 16108
rect 4023 16068 4068 16096
rect 4062 16056 4068 16068
rect 4120 16056 4126 16108
rect 5077 16099 5135 16105
rect 5077 16065 5089 16099
rect 5123 16065 5135 16099
rect 5077 16059 5135 16065
rect 1486 15988 1492 16040
rect 1544 16028 1550 16040
rect 5092 16028 5120 16059
rect 5626 16056 5632 16108
rect 5684 16096 5690 16108
rect 5813 16099 5871 16105
rect 5813 16096 5825 16099
rect 5684 16068 5825 16096
rect 5684 16056 5690 16068
rect 5813 16065 5825 16068
rect 5859 16065 5871 16099
rect 5813 16059 5871 16065
rect 6730 16056 6736 16108
rect 6788 16096 6794 16108
rect 7101 16099 7159 16105
rect 7101 16096 7113 16099
rect 6788 16068 7113 16096
rect 6788 16056 6794 16068
rect 7101 16065 7113 16068
rect 7147 16065 7159 16099
rect 7101 16059 7159 16065
rect 1544 16000 5120 16028
rect 1544 15988 1550 16000
rect 7116 15960 7144 16059
rect 7282 16056 7288 16108
rect 7340 16096 7346 16108
rect 7745 16099 7803 16105
rect 7745 16096 7757 16099
rect 7340 16068 7757 16096
rect 7340 16056 7346 16068
rect 7745 16065 7757 16068
rect 7791 16065 7803 16099
rect 7745 16059 7803 16065
rect 9125 16099 9183 16105
rect 9125 16065 9137 16099
rect 9171 16096 9183 16099
rect 9214 16096 9220 16108
rect 9171 16068 9220 16096
rect 9171 16065 9183 16068
rect 9125 16059 9183 16065
rect 9214 16056 9220 16068
rect 9272 16056 9278 16108
rect 10962 16096 10968 16108
rect 10612 16068 10968 16096
rect 7837 16031 7895 16037
rect 7837 15997 7849 16031
rect 7883 16028 7895 16031
rect 10612 16028 10640 16068
rect 10962 16056 10968 16068
rect 11020 16056 11026 16108
rect 14826 16096 14832 16108
rect 14787 16068 14832 16096
rect 14826 16056 14832 16068
rect 14884 16056 14890 16108
rect 17696 16105 17724 16136
rect 18506 16124 18512 16136
rect 18564 16124 18570 16176
rect 17037 16099 17095 16105
rect 17037 16065 17049 16099
rect 17083 16065 17095 16099
rect 17037 16059 17095 16065
rect 17681 16099 17739 16105
rect 17681 16065 17693 16099
rect 17727 16065 17739 16099
rect 17681 16059 17739 16065
rect 7883 16000 10640 16028
rect 10689 16031 10747 16037
rect 7883 15997 7895 16000
rect 7837 15991 7895 15997
rect 10689 15997 10701 16031
rect 10735 15997 10747 16031
rect 10689 15991 10747 15997
rect 12161 16031 12219 16037
rect 12161 15997 12173 16031
rect 12207 16028 12219 16031
rect 12342 16028 12348 16040
rect 12207 16000 12348 16028
rect 12207 15997 12219 16000
rect 12161 15991 12219 15997
rect 10594 15960 10600 15972
rect 7116 15932 10600 15960
rect 10594 15920 10600 15932
rect 10652 15920 10658 15972
rect 10704 15960 10732 15991
rect 12342 15988 12348 16000
rect 12400 15988 12406 16040
rect 12802 16028 12808 16040
rect 12763 16000 12808 16028
rect 12802 15988 12808 16000
rect 12860 15988 12866 16040
rect 13357 16031 13415 16037
rect 13357 15997 13369 16031
rect 13403 16028 13415 16031
rect 13446 16028 13452 16040
rect 13403 16000 13452 16028
rect 13403 15997 13415 16000
rect 13357 15991 13415 15997
rect 13446 15988 13452 16000
rect 13504 15988 13510 16040
rect 13722 15988 13728 16040
rect 13780 16028 13786 16040
rect 15286 16028 15292 16040
rect 13780 16000 15292 16028
rect 13780 15988 13786 16000
rect 15286 15988 15292 16000
rect 15344 15988 15350 16040
rect 15562 16028 15568 16040
rect 15523 16000 15568 16028
rect 15562 15988 15568 16000
rect 15620 15988 15626 16040
rect 17052 16028 17080 16059
rect 17126 16028 17132 16040
rect 17052 16000 17132 16028
rect 17126 15988 17132 16000
rect 17184 15988 17190 16040
rect 18414 16028 18420 16040
rect 18375 16000 18420 16028
rect 18414 15988 18420 16000
rect 18472 15988 18478 16040
rect 18690 16028 18696 16040
rect 18651 16000 18696 16028
rect 18690 15988 18696 16000
rect 18748 15988 18754 16040
rect 15194 15960 15200 15972
rect 10704 15932 15200 15960
rect 15194 15920 15200 15932
rect 15252 15920 15258 15972
rect 15838 15920 15844 15972
rect 15896 15960 15902 15972
rect 16114 15960 16120 15972
rect 15896 15932 16120 15960
rect 15896 15920 15902 15932
rect 16114 15920 16120 15932
rect 16172 15920 16178 15972
rect 17310 15960 17316 15972
rect 17060 15932 17316 15960
rect 1762 15892 1768 15904
rect 1723 15864 1768 15892
rect 1762 15852 1768 15864
rect 1820 15852 1826 15904
rect 2317 15895 2375 15901
rect 2317 15861 2329 15895
rect 2363 15892 2375 15895
rect 2590 15892 2596 15904
rect 2363 15864 2596 15892
rect 2363 15861 2375 15864
rect 2317 15855 2375 15861
rect 2590 15852 2596 15864
rect 2648 15852 2654 15904
rect 5905 15895 5963 15901
rect 5905 15861 5917 15895
rect 5951 15892 5963 15895
rect 6546 15892 6552 15904
rect 5951 15864 6552 15892
rect 5951 15861 5963 15864
rect 5905 15855 5963 15861
rect 6546 15852 6552 15864
rect 6604 15852 6610 15904
rect 7193 15895 7251 15901
rect 7193 15861 7205 15895
rect 7239 15892 7251 15895
rect 8570 15892 8576 15904
rect 7239 15864 8576 15892
rect 7239 15861 7251 15864
rect 7193 15855 7251 15861
rect 8570 15852 8576 15864
rect 8628 15852 8634 15904
rect 9214 15852 9220 15904
rect 9272 15892 9278 15904
rect 13538 15892 13544 15904
rect 9272 15864 13544 15892
rect 9272 15852 9278 15864
rect 13538 15852 13544 15864
rect 13596 15852 13602 15904
rect 14921 15895 14979 15901
rect 14921 15861 14933 15895
rect 14967 15892 14979 15895
rect 17060 15892 17088 15932
rect 17310 15920 17316 15932
rect 17368 15920 17374 15972
rect 14967 15864 17088 15892
rect 17129 15895 17187 15901
rect 14967 15861 14979 15864
rect 14921 15855 14979 15861
rect 17129 15861 17141 15895
rect 17175 15892 17187 15895
rect 17586 15892 17592 15904
rect 17175 15864 17592 15892
rect 17175 15861 17187 15864
rect 17129 15855 17187 15861
rect 17586 15852 17592 15864
rect 17644 15852 17650 15904
rect 17773 15895 17831 15901
rect 17773 15861 17785 15895
rect 17819 15892 17831 15895
rect 17862 15892 17868 15904
rect 17819 15864 17868 15892
rect 17819 15861 17831 15864
rect 17773 15855 17831 15861
rect 17862 15852 17868 15864
rect 17920 15852 17926 15904
rect 19260 15892 19288 16204
rect 19978 16192 19984 16244
rect 20036 16232 20042 16244
rect 25685 16235 25743 16241
rect 25685 16232 25697 16235
rect 20036 16204 25697 16232
rect 20036 16192 20042 16204
rect 25685 16201 25697 16204
rect 25731 16201 25743 16235
rect 28166 16232 28172 16244
rect 28127 16204 28172 16232
rect 25685 16195 25743 16201
rect 28166 16192 28172 16204
rect 28224 16192 28230 16244
rect 28258 16192 28264 16244
rect 28316 16232 28322 16244
rect 30650 16232 30656 16244
rect 28316 16204 30656 16232
rect 28316 16192 28322 16204
rect 30650 16192 30656 16204
rect 30708 16192 30714 16244
rect 20070 16164 20076 16176
rect 20031 16136 20076 16164
rect 20070 16124 20076 16136
rect 20128 16124 20134 16176
rect 20346 16124 20352 16176
rect 20404 16164 20410 16176
rect 20714 16164 20720 16176
rect 20404 16136 20720 16164
rect 20404 16124 20410 16136
rect 20714 16124 20720 16136
rect 20772 16124 20778 16176
rect 21177 16167 21235 16173
rect 21177 16133 21189 16167
rect 21223 16164 21235 16167
rect 22833 16167 22891 16173
rect 22833 16164 22845 16167
rect 21223 16136 22845 16164
rect 21223 16133 21235 16136
rect 21177 16127 21235 16133
rect 22833 16133 22845 16136
rect 22879 16133 22891 16167
rect 33594 16164 33600 16176
rect 22833 16127 22891 16133
rect 27540 16136 33600 16164
rect 21082 16096 21088 16108
rect 21043 16068 21088 16096
rect 21082 16056 21088 16068
rect 21140 16056 21146 16108
rect 21910 16056 21916 16108
rect 21968 16096 21974 16108
rect 22005 16099 22063 16105
rect 22005 16096 22017 16099
rect 21968 16068 22017 16096
rect 21968 16056 21974 16068
rect 22005 16065 22017 16068
rect 22051 16065 22063 16099
rect 22005 16059 22063 16065
rect 23658 16056 23664 16108
rect 23716 16096 23722 16108
rect 27540 16105 27568 16136
rect 33594 16124 33600 16136
rect 33652 16124 33658 16176
rect 25225 16099 25283 16105
rect 25225 16096 25237 16099
rect 23716 16068 25237 16096
rect 23716 16056 23722 16068
rect 25225 16065 25237 16068
rect 25271 16065 25283 16099
rect 25225 16059 25283 16065
rect 27525 16099 27583 16105
rect 27525 16065 27537 16099
rect 27571 16065 27583 16099
rect 28813 16099 28871 16105
rect 28813 16096 28825 16099
rect 27525 16059 27583 16065
rect 27632 16068 28825 16096
rect 19981 16031 20039 16037
rect 19981 15997 19993 16031
rect 20027 16028 20039 16031
rect 22094 16028 22100 16040
rect 20027 16000 22100 16028
rect 20027 15997 20039 16000
rect 19981 15991 20039 15997
rect 22094 15988 22100 16000
rect 22152 15988 22158 16040
rect 22741 16031 22799 16037
rect 22741 15997 22753 16031
rect 22787 16028 22799 16031
rect 22922 16028 22928 16040
rect 22787 16000 22928 16028
rect 22787 15997 22799 16000
rect 22741 15991 22799 15997
rect 22922 15988 22928 16000
rect 22980 15988 22986 16040
rect 23106 16028 23112 16040
rect 23067 16000 23112 16028
rect 23106 15988 23112 16000
rect 23164 15988 23170 16040
rect 25041 16031 25099 16037
rect 25041 15997 25053 16031
rect 25087 15997 25099 16031
rect 25041 15991 25099 15997
rect 20070 15920 20076 15972
rect 20128 15960 20134 15972
rect 20530 15960 20536 15972
rect 20128 15932 20536 15960
rect 20128 15920 20134 15932
rect 20530 15920 20536 15932
rect 20588 15920 20594 15972
rect 23198 15960 23204 15972
rect 20640 15932 23204 15960
rect 20640 15892 20668 15932
rect 23198 15920 23204 15932
rect 23256 15920 23262 15972
rect 25056 15960 25084 15991
rect 27154 15988 27160 16040
rect 27212 16028 27218 16040
rect 27632 16028 27660 16068
rect 28813 16065 28825 16068
rect 28859 16065 28871 16099
rect 30285 16099 30343 16105
rect 30285 16096 30297 16099
rect 28813 16059 28871 16065
rect 29012 16068 30297 16096
rect 27212 16000 27660 16028
rect 27709 16031 27767 16037
rect 27212 15988 27218 16000
rect 27709 15997 27721 16031
rect 27755 16028 27767 16031
rect 28534 16028 28540 16040
rect 27755 16000 28540 16028
rect 27755 15997 27767 16000
rect 27709 15991 27767 15997
rect 28534 15988 28540 16000
rect 28592 15988 28598 16040
rect 27430 15960 27436 15972
rect 25056 15932 27436 15960
rect 27430 15920 27436 15932
rect 27488 15920 27494 15972
rect 28350 15920 28356 15972
rect 28408 15960 28414 15972
rect 29012 15960 29040 16068
rect 30285 16065 30297 16068
rect 30331 16065 30343 16099
rect 30285 16059 30343 16065
rect 30929 16099 30987 16105
rect 30929 16065 30941 16099
rect 30975 16065 30987 16099
rect 38010 16096 38016 16108
rect 37971 16068 38016 16096
rect 30929 16059 30987 16065
rect 29270 16028 29276 16040
rect 29231 16000 29276 16028
rect 29270 15988 29276 16000
rect 29328 15988 29334 16040
rect 30944 16028 30972 16059
rect 38010 16056 38016 16068
rect 38068 16056 38074 16108
rect 30116 16000 30972 16028
rect 30116 15969 30144 16000
rect 28408 15932 29040 15960
rect 30101 15963 30159 15969
rect 28408 15920 28414 15932
rect 30101 15929 30113 15963
rect 30147 15929 30159 15963
rect 30101 15923 30159 15929
rect 30190 15920 30196 15972
rect 30248 15960 30254 15972
rect 34790 15960 34796 15972
rect 30248 15932 34796 15960
rect 30248 15920 30254 15932
rect 34790 15920 34796 15932
rect 34848 15920 34854 15972
rect 19260 15864 20668 15892
rect 22094 15852 22100 15904
rect 22152 15892 22158 15904
rect 22152 15864 22197 15892
rect 22152 15852 22158 15864
rect 24210 15852 24216 15904
rect 24268 15892 24274 15904
rect 28258 15892 28264 15904
rect 24268 15864 28264 15892
rect 24268 15852 24274 15864
rect 28258 15852 28264 15864
rect 28316 15852 28322 15904
rect 28629 15895 28687 15901
rect 28629 15861 28641 15895
rect 28675 15892 28687 15895
rect 29914 15892 29920 15904
rect 28675 15864 29920 15892
rect 28675 15861 28687 15864
rect 28629 15855 28687 15861
rect 29914 15852 29920 15864
rect 29972 15852 29978 15904
rect 30742 15892 30748 15904
rect 30703 15864 30748 15892
rect 30742 15852 30748 15864
rect 30800 15852 30806 15904
rect 38194 15892 38200 15904
rect 38155 15864 38200 15892
rect 38194 15852 38200 15864
rect 38252 15852 38258 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 1765 15691 1823 15697
rect 1765 15657 1777 15691
rect 1811 15688 1823 15691
rect 2498 15688 2504 15700
rect 1811 15660 2504 15688
rect 1811 15657 1823 15660
rect 1765 15651 1823 15657
rect 2498 15648 2504 15660
rect 2556 15648 2562 15700
rect 6454 15648 6460 15700
rect 6512 15688 6518 15700
rect 12526 15688 12532 15700
rect 6512 15660 12532 15688
rect 6512 15648 6518 15660
rect 12526 15648 12532 15660
rect 12584 15648 12590 15700
rect 12618 15648 12624 15700
rect 12676 15688 12682 15700
rect 15286 15688 15292 15700
rect 12676 15660 15292 15688
rect 12676 15648 12682 15660
rect 15286 15648 15292 15660
rect 15344 15648 15350 15700
rect 15838 15648 15844 15700
rect 15896 15688 15902 15700
rect 16114 15688 16120 15700
rect 15896 15660 16120 15688
rect 15896 15648 15902 15660
rect 16114 15648 16120 15660
rect 16172 15648 16178 15700
rect 23106 15688 23112 15700
rect 16684 15660 23112 15688
rect 5258 15580 5264 15632
rect 5316 15620 5322 15632
rect 8478 15620 8484 15632
rect 5316 15592 8484 15620
rect 5316 15580 5322 15592
rect 8478 15580 8484 15592
rect 8536 15580 8542 15632
rect 9582 15580 9588 15632
rect 9640 15620 9646 15632
rect 12342 15620 12348 15632
rect 9640 15592 12348 15620
rect 9640 15580 9646 15592
rect 12342 15580 12348 15592
rect 12400 15580 12406 15632
rect 12452 15592 15608 15620
rect 6549 15555 6607 15561
rect 6549 15521 6561 15555
rect 6595 15552 6607 15555
rect 8018 15552 8024 15564
rect 6595 15524 8024 15552
rect 6595 15521 6607 15524
rect 6549 15515 6607 15521
rect 8018 15512 8024 15524
rect 8076 15512 8082 15564
rect 8846 15552 8852 15564
rect 8312 15524 8852 15552
rect 1670 15444 1676 15496
rect 1728 15484 1734 15496
rect 1949 15487 2007 15493
rect 1949 15484 1961 15487
rect 1728 15456 1961 15484
rect 1728 15444 1734 15456
rect 1949 15453 1961 15456
rect 1995 15453 2007 15487
rect 1949 15447 2007 15453
rect 4525 15487 4583 15493
rect 4525 15453 4537 15487
rect 4571 15484 4583 15487
rect 4890 15484 4896 15496
rect 4571 15456 4896 15484
rect 4571 15453 4583 15456
rect 4525 15447 4583 15453
rect 4890 15444 4896 15456
rect 4948 15444 4954 15496
rect 5074 15444 5080 15496
rect 5132 15484 5138 15496
rect 5169 15487 5227 15493
rect 5169 15484 5181 15487
rect 5132 15456 5181 15484
rect 5132 15444 5138 15456
rect 5169 15453 5181 15456
rect 5215 15453 5227 15487
rect 5810 15484 5816 15496
rect 5771 15456 5816 15484
rect 5169 15447 5227 15453
rect 5810 15444 5816 15456
rect 5868 15444 5874 15496
rect 6454 15484 6460 15496
rect 6415 15456 6460 15484
rect 6454 15444 6460 15456
rect 6512 15444 6518 15496
rect 7285 15487 7343 15493
rect 7285 15453 7297 15487
rect 7331 15484 7343 15487
rect 7374 15484 7380 15496
rect 7331 15456 7380 15484
rect 7331 15453 7343 15456
rect 7285 15447 7343 15453
rect 7374 15444 7380 15456
rect 7432 15444 7438 15496
rect 7745 15487 7803 15493
rect 7745 15453 7757 15487
rect 7791 15484 7803 15487
rect 8312 15484 8340 15524
rect 8846 15512 8852 15524
rect 8904 15512 8910 15564
rect 9214 15552 9220 15564
rect 9175 15524 9220 15552
rect 9214 15512 9220 15524
rect 9272 15512 9278 15564
rect 9766 15552 9772 15564
rect 9727 15524 9772 15552
rect 9766 15512 9772 15524
rect 9824 15512 9830 15564
rect 9858 15512 9864 15564
rect 9916 15552 9922 15564
rect 11885 15555 11943 15561
rect 9916 15524 11744 15552
rect 9916 15512 9922 15524
rect 7791 15456 8340 15484
rect 8389 15487 8447 15493
rect 7791 15453 7803 15456
rect 7745 15447 7803 15453
rect 8389 15453 8401 15487
rect 8435 15484 8447 15487
rect 8478 15484 8484 15496
rect 8435 15456 8484 15484
rect 8435 15453 8447 15456
rect 8389 15447 8447 15453
rect 8478 15444 8484 15456
rect 8536 15444 8542 15496
rect 11716 15484 11744 15524
rect 11885 15521 11897 15555
rect 11931 15552 11943 15555
rect 12452 15552 12480 15592
rect 11931 15524 12480 15552
rect 12713 15555 12771 15561
rect 11931 15521 11943 15524
rect 11885 15515 11943 15521
rect 12713 15521 12725 15555
rect 12759 15552 12771 15555
rect 13814 15552 13820 15564
rect 12759 15524 13820 15552
rect 12759 15521 12771 15524
rect 12713 15515 12771 15521
rect 13814 15512 13820 15524
rect 13872 15512 13878 15564
rect 13906 15512 13912 15564
rect 13964 15552 13970 15564
rect 15580 15561 15608 15592
rect 14553 15555 14611 15561
rect 14553 15552 14565 15555
rect 13964 15524 14565 15552
rect 13964 15512 13970 15524
rect 14553 15521 14565 15524
rect 14599 15521 14611 15555
rect 14553 15515 14611 15521
rect 15565 15555 15623 15561
rect 15565 15521 15577 15555
rect 15611 15552 15623 15555
rect 16684 15552 16712 15660
rect 23106 15648 23112 15660
rect 23164 15648 23170 15700
rect 24394 15648 24400 15700
rect 24452 15688 24458 15700
rect 27985 15691 28043 15697
rect 24452 15660 26280 15688
rect 24452 15648 24458 15660
rect 18230 15620 18236 15632
rect 15611 15524 16712 15552
rect 17512 15592 18236 15620
rect 15611 15521 15623 15524
rect 15565 15515 15623 15521
rect 17512 15493 17540 15592
rect 18230 15580 18236 15592
rect 18288 15580 18294 15632
rect 18414 15580 18420 15632
rect 18472 15620 18478 15632
rect 20622 15620 20628 15632
rect 18472 15592 20628 15620
rect 18472 15580 18478 15592
rect 20622 15580 20628 15592
rect 20680 15620 20686 15632
rect 24210 15620 24216 15632
rect 20680 15592 24216 15620
rect 20680 15580 20686 15592
rect 24210 15580 24216 15592
rect 24268 15580 24274 15632
rect 26142 15620 26148 15632
rect 24688 15592 26148 15620
rect 18141 15555 18199 15561
rect 18141 15521 18153 15555
rect 18187 15552 18199 15555
rect 19978 15552 19984 15564
rect 18187 15524 19984 15552
rect 18187 15521 18199 15524
rect 18141 15515 18199 15521
rect 19978 15512 19984 15524
rect 20036 15512 20042 15564
rect 20438 15552 20444 15564
rect 20351 15524 20444 15552
rect 20438 15512 20444 15524
rect 20496 15552 20502 15564
rect 20714 15552 20720 15564
rect 20496 15524 20720 15552
rect 20496 15512 20502 15524
rect 20714 15512 20720 15524
rect 20772 15512 20778 15564
rect 22094 15512 22100 15564
rect 22152 15552 22158 15564
rect 24581 15555 24639 15561
rect 24581 15552 24593 15555
rect 22152 15524 24593 15552
rect 22152 15512 22158 15524
rect 24581 15521 24593 15524
rect 24627 15521 24639 15555
rect 24581 15515 24639 15521
rect 17497 15487 17555 15493
rect 11716 15456 12007 15484
rect 3602 15376 3608 15428
rect 3660 15416 3666 15428
rect 7558 15416 7564 15428
rect 3660 15388 7564 15416
rect 3660 15376 3666 15388
rect 7558 15376 7564 15388
rect 7616 15376 7622 15428
rect 7837 15419 7895 15425
rect 7837 15385 7849 15419
rect 7883 15416 7895 15419
rect 9309 15419 9367 15425
rect 9309 15416 9321 15419
rect 7883 15388 8156 15416
rect 7883 15385 7895 15388
rect 7837 15379 7895 15385
rect 2406 15348 2412 15360
rect 2367 15320 2412 15348
rect 2406 15308 2412 15320
rect 2464 15308 2470 15360
rect 4617 15351 4675 15357
rect 4617 15317 4629 15351
rect 4663 15348 4675 15351
rect 5166 15348 5172 15360
rect 4663 15320 5172 15348
rect 4663 15317 4675 15320
rect 4617 15311 4675 15317
rect 5166 15308 5172 15320
rect 5224 15308 5230 15360
rect 5261 15351 5319 15357
rect 5261 15317 5273 15351
rect 5307 15348 5319 15351
rect 5350 15348 5356 15360
rect 5307 15320 5356 15348
rect 5307 15317 5319 15320
rect 5261 15311 5319 15317
rect 5350 15308 5356 15320
rect 5408 15308 5414 15360
rect 5905 15351 5963 15357
rect 5905 15317 5917 15351
rect 5951 15348 5963 15351
rect 6822 15348 6828 15360
rect 5951 15320 6828 15348
rect 5951 15317 5963 15320
rect 5905 15311 5963 15317
rect 6822 15308 6828 15320
rect 6880 15308 6886 15360
rect 7101 15351 7159 15357
rect 7101 15317 7113 15351
rect 7147 15348 7159 15351
rect 7190 15348 7196 15360
rect 7147 15320 7196 15348
rect 7147 15317 7159 15320
rect 7101 15311 7159 15317
rect 7190 15308 7196 15320
rect 7248 15308 7254 15360
rect 8128 15348 8156 15388
rect 8404 15388 9321 15416
rect 8404 15348 8432 15388
rect 9309 15385 9321 15388
rect 9355 15385 9367 15419
rect 9309 15379 9367 15385
rect 9766 15376 9772 15428
rect 9824 15416 9830 15428
rect 10870 15416 10876 15428
rect 9824 15388 10876 15416
rect 9824 15376 9830 15388
rect 10870 15376 10876 15388
rect 10928 15376 10934 15428
rect 10962 15376 10968 15428
rect 11020 15416 11026 15428
rect 11020 15388 11065 15416
rect 11020 15376 11026 15388
rect 8128 15320 8432 15348
rect 8481 15351 8539 15357
rect 8481 15317 8493 15351
rect 8527 15348 8539 15351
rect 11882 15348 11888 15360
rect 8527 15320 11888 15348
rect 8527 15317 8539 15320
rect 8481 15311 8539 15317
rect 11882 15308 11888 15320
rect 11940 15308 11946 15360
rect 11979 15348 12007 15456
rect 17497 15453 17509 15487
rect 17543 15453 17555 15487
rect 17497 15447 17555 15453
rect 17681 15487 17739 15493
rect 17681 15453 17693 15487
rect 17727 15453 17739 15487
rect 18690 15484 18696 15496
rect 18651 15456 18696 15484
rect 17681 15447 17739 15453
rect 12805 15419 12863 15425
rect 12805 15416 12817 15419
rect 12801 15385 12817 15416
rect 12851 15385 12863 15419
rect 12801 15379 12863 15385
rect 13725 15419 13783 15425
rect 13725 15385 13737 15419
rect 13771 15416 13783 15419
rect 14366 15416 14372 15428
rect 13771 15388 14372 15416
rect 13771 15385 13783 15388
rect 13725 15379 13783 15385
rect 12801 15348 12829 15379
rect 14366 15376 14372 15388
rect 14424 15376 14430 15428
rect 14642 15416 14648 15428
rect 14603 15388 14648 15416
rect 14642 15376 14648 15388
rect 14700 15376 14706 15428
rect 15562 15376 15568 15428
rect 15620 15416 15626 15428
rect 16117 15419 16175 15425
rect 16117 15416 16129 15419
rect 15620 15388 16129 15416
rect 15620 15376 15626 15388
rect 16117 15385 16129 15388
rect 16163 15385 16175 15419
rect 16117 15379 16175 15385
rect 16945 15419 17003 15425
rect 16945 15385 16957 15419
rect 16991 15416 17003 15419
rect 17126 15416 17132 15428
rect 16991 15388 17132 15416
rect 16991 15385 17003 15388
rect 16945 15379 17003 15385
rect 17126 15376 17132 15388
rect 17184 15376 17190 15428
rect 17696 15416 17724 15447
rect 18690 15444 18696 15456
rect 18748 15444 18754 15496
rect 19334 15444 19340 15496
rect 19392 15484 19398 15496
rect 19705 15487 19763 15493
rect 19705 15484 19717 15487
rect 19392 15456 19717 15484
rect 19392 15444 19398 15456
rect 19705 15453 19717 15456
rect 19751 15453 19763 15487
rect 19705 15447 19763 15453
rect 21913 15487 21971 15493
rect 21913 15453 21925 15487
rect 21959 15484 21971 15487
rect 22002 15484 22008 15496
rect 21959 15456 22008 15484
rect 21959 15453 21971 15456
rect 21913 15447 21971 15453
rect 22002 15444 22008 15456
rect 22060 15444 22066 15496
rect 22370 15444 22376 15496
rect 22428 15484 22434 15496
rect 22557 15487 22615 15493
rect 22557 15484 22569 15487
rect 22428 15456 22569 15484
rect 22428 15444 22434 15456
rect 22557 15453 22569 15456
rect 22603 15453 22615 15487
rect 22557 15447 22615 15453
rect 23845 15487 23903 15493
rect 23845 15453 23857 15487
rect 23891 15484 23903 15487
rect 24688 15484 24716 15592
rect 26142 15580 26148 15592
rect 26200 15580 26206 15632
rect 26252 15620 26280 15660
rect 27985 15657 27997 15691
rect 28031 15688 28043 15691
rect 28166 15688 28172 15700
rect 28031 15660 28172 15688
rect 28031 15657 28043 15660
rect 27985 15651 28043 15657
rect 28166 15648 28172 15660
rect 28224 15648 28230 15700
rect 28534 15688 28540 15700
rect 28495 15660 28540 15688
rect 28534 15648 28540 15660
rect 28592 15648 28598 15700
rect 30190 15620 30196 15632
rect 26252 15592 30196 15620
rect 30190 15580 30196 15592
rect 30248 15580 30254 15632
rect 25225 15555 25283 15561
rect 25225 15521 25237 15555
rect 25271 15552 25283 15555
rect 26418 15552 26424 15564
rect 25271 15524 26424 15552
rect 25271 15521 25283 15524
rect 25225 15515 25283 15521
rect 26418 15512 26424 15524
rect 26476 15512 26482 15564
rect 27525 15555 27583 15561
rect 27525 15521 27537 15555
rect 27571 15552 27583 15555
rect 30742 15552 30748 15564
rect 27571 15524 30748 15552
rect 27571 15521 27583 15524
rect 27525 15515 27583 15521
rect 30742 15512 30748 15524
rect 30800 15512 30806 15564
rect 23891 15456 24716 15484
rect 24765 15487 24823 15493
rect 23891 15453 23903 15456
rect 23845 15447 23903 15453
rect 24765 15453 24777 15487
rect 24811 15484 24823 15487
rect 26050 15484 26056 15496
rect 24811 15456 26056 15484
rect 24811 15453 24823 15456
rect 24765 15447 24823 15453
rect 26050 15444 26056 15456
rect 26108 15444 26114 15496
rect 26510 15484 26516 15496
rect 26471 15456 26516 15484
rect 26510 15444 26516 15456
rect 26568 15444 26574 15496
rect 27341 15487 27399 15493
rect 27341 15453 27353 15487
rect 27387 15484 27399 15487
rect 27430 15484 27436 15496
rect 27387 15456 27436 15484
rect 27387 15453 27399 15456
rect 27341 15447 27399 15453
rect 27430 15444 27436 15456
rect 27488 15444 27494 15496
rect 28350 15444 28356 15496
rect 28408 15484 28414 15496
rect 28445 15487 28503 15493
rect 28445 15484 28457 15487
rect 28408 15456 28457 15484
rect 28408 15444 28414 15456
rect 28445 15453 28457 15456
rect 28491 15453 28503 15487
rect 29914 15484 29920 15496
rect 29875 15456 29920 15484
rect 28445 15447 28503 15453
rect 29914 15444 29920 15456
rect 29972 15444 29978 15496
rect 17236 15388 17724 15416
rect 11979 15320 12829 15348
rect 13078 15308 13084 15360
rect 13136 15348 13142 15360
rect 13446 15348 13452 15360
rect 13136 15320 13452 15348
rect 13136 15308 13142 15320
rect 13446 15308 13452 15320
rect 13504 15308 13510 15360
rect 15010 15308 15016 15360
rect 15068 15348 15074 15360
rect 17236 15348 17264 15388
rect 17954 15376 17960 15428
rect 18012 15416 18018 15428
rect 20070 15416 20076 15428
rect 18012 15388 20076 15416
rect 18012 15376 18018 15388
rect 20070 15376 20076 15388
rect 20128 15376 20134 15428
rect 20533 15419 20591 15425
rect 20533 15385 20545 15419
rect 20579 15385 20591 15419
rect 20533 15379 20591 15385
rect 21453 15419 21511 15425
rect 21453 15385 21465 15419
rect 21499 15416 21511 15419
rect 23658 15416 23664 15428
rect 21499 15388 23664 15416
rect 21499 15385 21511 15388
rect 21453 15379 21511 15385
rect 15068 15320 17264 15348
rect 18785 15351 18843 15357
rect 15068 15308 15074 15320
rect 18785 15317 18797 15351
rect 18831 15348 18843 15351
rect 19518 15348 19524 15360
rect 18831 15320 19524 15348
rect 18831 15317 18843 15320
rect 18785 15311 18843 15317
rect 19518 15308 19524 15320
rect 19576 15308 19582 15360
rect 19797 15351 19855 15357
rect 19797 15317 19809 15351
rect 19843 15348 19855 15351
rect 20548 15348 20576 15379
rect 23658 15376 23664 15388
rect 23716 15416 23722 15428
rect 24394 15416 24400 15428
rect 23716 15388 24400 15416
rect 23716 15376 23722 15388
rect 24394 15376 24400 15388
rect 24452 15376 24458 15428
rect 25685 15419 25743 15425
rect 25685 15416 25697 15419
rect 24780 15388 25697 15416
rect 24780 15360 24808 15388
rect 25685 15385 25697 15388
rect 25731 15385 25743 15419
rect 38102 15416 38108 15428
rect 38063 15388 38108 15416
rect 25685 15379 25743 15385
rect 38102 15376 38108 15388
rect 38160 15376 38166 15428
rect 19843 15320 20576 15348
rect 19843 15317 19855 15320
rect 19797 15311 19855 15317
rect 21174 15308 21180 15360
rect 21232 15348 21238 15360
rect 22005 15351 22063 15357
rect 22005 15348 22017 15351
rect 21232 15320 22017 15348
rect 21232 15308 21238 15320
rect 22005 15317 22017 15320
rect 22051 15317 22063 15351
rect 22005 15311 22063 15317
rect 22649 15351 22707 15357
rect 22649 15317 22661 15351
rect 22695 15348 22707 15351
rect 23290 15348 23296 15360
rect 22695 15320 23296 15348
rect 22695 15317 22707 15320
rect 22649 15311 22707 15317
rect 23290 15308 23296 15320
rect 23348 15308 23354 15360
rect 23937 15351 23995 15357
rect 23937 15317 23949 15351
rect 23983 15348 23995 15351
rect 24670 15348 24676 15360
rect 23983 15320 24676 15348
rect 23983 15317 23995 15320
rect 23937 15311 23995 15317
rect 24670 15308 24676 15320
rect 24728 15308 24734 15360
rect 24762 15308 24768 15360
rect 24820 15308 24826 15360
rect 26234 15308 26240 15360
rect 26292 15348 26298 15360
rect 26329 15351 26387 15357
rect 26329 15348 26341 15351
rect 26292 15320 26341 15348
rect 26292 15308 26298 15320
rect 26329 15317 26341 15320
rect 26375 15317 26387 15351
rect 26329 15311 26387 15317
rect 28994 15308 29000 15360
rect 29052 15348 29058 15360
rect 29733 15351 29791 15357
rect 29733 15348 29745 15351
rect 29052 15320 29745 15348
rect 29052 15308 29058 15320
rect 29733 15317 29745 15320
rect 29779 15317 29791 15351
rect 38194 15348 38200 15360
rect 38155 15320 38200 15348
rect 29733 15311 29791 15317
rect 38194 15308 38200 15320
rect 38252 15308 38258 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 6917 15147 6975 15153
rect 6917 15113 6929 15147
rect 6963 15144 6975 15147
rect 17770 15144 17776 15156
rect 6963 15116 11284 15144
rect 6963 15113 6975 15116
rect 6917 15107 6975 15113
rect 5074 15076 5080 15088
rect 3896 15048 5080 15076
rect 1670 14968 1676 15020
rect 1728 15008 1734 15020
rect 1765 15011 1823 15017
rect 1765 15008 1777 15011
rect 1728 14980 1777 15008
rect 1728 14968 1734 14980
rect 1765 14977 1777 14980
rect 1811 14977 1823 15011
rect 2406 15008 2412 15020
rect 2367 14980 2412 15008
rect 1765 14971 1823 14977
rect 2406 14968 2412 14980
rect 2464 14968 2470 15020
rect 2590 15008 2596 15020
rect 2551 14980 2596 15008
rect 2590 14968 2596 14980
rect 2648 14968 2654 15020
rect 3896 15017 3924 15048
rect 5074 15036 5080 15048
rect 5132 15036 5138 15088
rect 5261 15079 5319 15085
rect 5261 15045 5273 15079
rect 5307 15076 5319 15079
rect 8849 15079 8907 15085
rect 8849 15076 8861 15079
rect 5307 15048 8861 15076
rect 5307 15045 5319 15048
rect 5261 15039 5319 15045
rect 8849 15045 8861 15048
rect 8895 15045 8907 15079
rect 10594 15076 10600 15088
rect 10555 15048 10600 15076
rect 8849 15039 8907 15045
rect 10594 15036 10600 15048
rect 10652 15036 10658 15088
rect 3881 15011 3939 15017
rect 3881 14977 3893 15011
rect 3927 14977 3939 15011
rect 3881 14971 3939 14977
rect 4982 14968 4988 15020
rect 5040 15008 5046 15020
rect 5169 15011 5227 15017
rect 5169 15008 5181 15011
rect 5040 14980 5181 15008
rect 5040 14968 5046 14980
rect 5169 14977 5181 14980
rect 5215 14977 5227 15011
rect 5810 15008 5816 15020
rect 5771 14980 5816 15008
rect 5169 14971 5227 14977
rect 5810 14968 5816 14980
rect 5868 14968 5874 15020
rect 5994 14968 6000 15020
rect 6052 15008 6058 15020
rect 6641 15011 6699 15017
rect 6641 15008 6653 15011
rect 6052 14980 6653 15008
rect 6052 14968 6058 14980
rect 6641 14977 6653 14980
rect 6687 14977 6699 15011
rect 6641 14971 6699 14977
rect 7466 14968 7472 15020
rect 7524 15008 7530 15020
rect 8018 15008 8024 15020
rect 7524 14980 8024 15008
rect 7524 14968 7530 14980
rect 8018 14968 8024 14980
rect 8076 14968 8082 15020
rect 11256 15008 11284 15116
rect 12728 15116 14688 15144
rect 12526 15036 12532 15088
rect 12584 15076 12590 15088
rect 12728 15085 12756 15116
rect 12713 15079 12771 15085
rect 12713 15076 12725 15079
rect 12584 15048 12725 15076
rect 12584 15036 12590 15048
rect 12713 15045 12725 15048
rect 12759 15045 12771 15079
rect 12713 15039 12771 15045
rect 13078 15036 13084 15088
rect 13136 15076 13142 15088
rect 13357 15079 13415 15085
rect 13357 15076 13369 15079
rect 13136 15048 13369 15076
rect 13136 15036 13142 15048
rect 13357 15045 13369 15048
rect 13403 15045 13415 15079
rect 13357 15039 13415 15045
rect 13449 15079 13507 15085
rect 13449 15045 13461 15079
rect 13495 15076 13507 15079
rect 14550 15076 14556 15088
rect 13495 15048 14556 15076
rect 13495 15045 13507 15048
rect 13449 15039 13507 15045
rect 14550 15036 14556 15048
rect 14608 15036 14614 15088
rect 14660 15076 14688 15116
rect 16211 15116 17776 15144
rect 14660 15048 16160 15076
rect 11606 15008 11612 15020
rect 11256 14980 11612 15008
rect 11606 14968 11612 14980
rect 11664 15008 11670 15020
rect 12161 15011 12219 15017
rect 12161 15008 12173 15011
rect 11664 14980 12173 15008
rect 11664 14968 11670 14980
rect 12161 14977 12173 14980
rect 12207 14977 12219 15011
rect 14918 15008 14924 15020
rect 14831 14980 14924 15008
rect 12161 14971 12219 14977
rect 4525 14943 4583 14949
rect 4525 14909 4537 14943
rect 4571 14940 4583 14943
rect 7558 14940 7564 14952
rect 4571 14912 7564 14940
rect 4571 14909 4583 14912
rect 4525 14903 4583 14909
rect 7558 14900 7564 14912
rect 7616 14900 7622 14952
rect 8386 14900 8392 14952
rect 8444 14940 8450 14952
rect 8758 14943 8816 14949
rect 8444 14928 8708 14940
rect 8758 14928 8770 14943
rect 8444 14912 8770 14928
rect 8444 14900 8450 14912
rect 8680 14909 8770 14912
rect 8804 14909 8816 14943
rect 9122 14940 9128 14952
rect 9083 14912 9128 14940
rect 8680 14903 8816 14909
rect 8680 14900 8800 14903
rect 9122 14900 9128 14912
rect 9180 14940 9186 14952
rect 9674 14940 9680 14952
rect 9180 14912 9680 14940
rect 9180 14900 9186 14912
rect 9674 14900 9680 14912
rect 9732 14900 9738 14952
rect 10226 14900 10232 14952
rect 10284 14940 10290 14952
rect 10505 14943 10563 14949
rect 10505 14940 10517 14943
rect 10284 14912 10517 14940
rect 10284 14900 10290 14912
rect 10505 14909 10517 14912
rect 10551 14909 10563 14943
rect 10505 14903 10563 14909
rect 11330 14900 11336 14952
rect 11388 14940 11394 14952
rect 11698 14940 11704 14952
rect 11388 14912 11704 14940
rect 11388 14900 11394 14912
rect 11698 14900 11704 14912
rect 11756 14900 11762 14952
rect 12176 14940 12204 14971
rect 14918 14968 14924 14980
rect 14976 15008 14982 15020
rect 15378 15008 15384 15020
rect 14976 14980 15384 15008
rect 14976 14968 14982 14980
rect 15378 14968 15384 14980
rect 15436 14968 15442 15020
rect 16132 15017 16160 15048
rect 16117 15011 16175 15017
rect 16117 14977 16129 15011
rect 16163 14977 16175 15011
rect 16117 14971 16175 14977
rect 12618 14940 12624 14952
rect 12176 14912 12624 14940
rect 12618 14900 12624 14912
rect 12676 14900 12682 14952
rect 14366 14940 14372 14952
rect 14327 14912 14372 14940
rect 14366 14900 14372 14912
rect 14424 14900 14430 14952
rect 15194 14940 15200 14952
rect 15155 14912 15200 14940
rect 15194 14900 15200 14912
rect 15252 14900 15258 14952
rect 16211 14940 16239 15116
rect 17770 15104 17776 15116
rect 17828 15144 17834 15156
rect 19518 15144 19524 15156
rect 17828 15116 19524 15144
rect 17828 15104 17834 15116
rect 19518 15104 19524 15116
rect 19576 15104 19582 15156
rect 20070 15104 20076 15156
rect 20128 15144 20134 15156
rect 22830 15144 22836 15156
rect 20128 15116 22836 15144
rect 20128 15104 20134 15116
rect 22830 15104 22836 15116
rect 22888 15104 22894 15156
rect 23198 15104 23204 15156
rect 23256 15144 23262 15156
rect 26050 15144 26056 15156
rect 23256 15116 24808 15144
rect 26011 15116 26056 15144
rect 23256 15104 23262 15116
rect 17586 15076 17592 15088
rect 17547 15048 17592 15076
rect 17586 15036 17592 15048
rect 17644 15036 17650 15088
rect 19797 15079 19855 15085
rect 19797 15045 19809 15079
rect 19843 15076 19855 15079
rect 20530 15076 20536 15088
rect 19843 15048 20536 15076
rect 19843 15045 19855 15048
rect 19797 15039 19855 15045
rect 20530 15036 20536 15048
rect 20588 15036 20594 15088
rect 22189 15079 22247 15085
rect 22189 15076 22201 15079
rect 20824 15048 22201 15076
rect 18966 15008 18972 15020
rect 18927 14980 18972 15008
rect 18966 14968 18972 14980
rect 19024 14968 19030 15020
rect 16040 14912 16239 14940
rect 5626 14832 5632 14884
rect 5684 14872 5690 14884
rect 10778 14872 10784 14884
rect 5684 14844 10784 14872
rect 5684 14832 5690 14844
rect 10778 14832 10784 14844
rect 10836 14872 10842 14884
rect 10962 14872 10968 14884
rect 10836 14844 10968 14872
rect 10836 14832 10842 14844
rect 10962 14832 10968 14844
rect 11020 14832 11026 14884
rect 11057 14875 11115 14881
rect 11057 14841 11069 14875
rect 11103 14872 11115 14875
rect 16040 14872 16068 14912
rect 16298 14900 16304 14952
rect 16356 14940 16362 14952
rect 17497 14943 17555 14949
rect 17497 14940 17509 14943
rect 16356 14912 17509 14940
rect 16356 14900 16362 14912
rect 17497 14909 17509 14912
rect 17543 14909 17555 14943
rect 18138 14940 18144 14952
rect 18099 14912 18144 14940
rect 17497 14903 17555 14909
rect 18138 14900 18144 14912
rect 18196 14900 18202 14952
rect 19705 14943 19763 14949
rect 19705 14909 19717 14943
rect 19751 14940 19763 14943
rect 19978 14940 19984 14952
rect 19751 14912 19984 14940
rect 19751 14909 19763 14912
rect 19705 14903 19763 14909
rect 19978 14900 19984 14912
rect 20036 14900 20042 14952
rect 20070 14900 20076 14952
rect 20128 14940 20134 14952
rect 20128 14912 20173 14940
rect 20128 14900 20134 14912
rect 20530 14900 20536 14952
rect 20588 14940 20594 14952
rect 20824 14940 20852 15048
rect 22189 15045 22201 15048
rect 22235 15045 22247 15079
rect 24670 15076 24676 15088
rect 24631 15048 24676 15076
rect 22189 15039 22247 15045
rect 24670 15036 24676 15048
rect 24728 15036 24734 15088
rect 24780 15076 24808 15116
rect 26050 15104 26056 15116
rect 26108 15104 26114 15156
rect 24780 15048 27200 15076
rect 26234 15008 26240 15020
rect 26195 14980 26240 15008
rect 26234 14968 26240 14980
rect 26292 14968 26298 15020
rect 27172 15017 27200 15048
rect 27157 15011 27215 15017
rect 27157 14977 27169 15011
rect 27203 14977 27215 15011
rect 27157 14971 27215 14977
rect 28629 15011 28687 15017
rect 28629 14977 28641 15011
rect 28675 15008 28687 15011
rect 28994 15008 29000 15020
rect 28675 14980 29000 15008
rect 28675 14977 28687 14980
rect 28629 14971 28687 14977
rect 28994 14968 29000 14980
rect 29052 14968 29058 15020
rect 29086 14968 29092 15020
rect 29144 15008 29150 15020
rect 29733 15011 29791 15017
rect 29733 15008 29745 15011
rect 29144 14980 29745 15008
rect 29144 14968 29150 14980
rect 29733 14977 29745 14980
rect 29779 14977 29791 15011
rect 29733 14971 29791 14977
rect 30466 14968 30472 15020
rect 30524 15008 30530 15020
rect 31205 15011 31263 15017
rect 31205 15008 31217 15011
rect 30524 14980 31217 15008
rect 30524 14968 30530 14980
rect 31205 14977 31217 14980
rect 31251 14977 31263 15011
rect 31205 14971 31263 14977
rect 31294 14968 31300 15020
rect 31352 15008 31358 15020
rect 33137 15011 33195 15017
rect 33137 15008 33149 15011
rect 31352 14980 33149 15008
rect 31352 14968 31358 14980
rect 33137 14977 33149 14980
rect 33183 14977 33195 15011
rect 33137 14971 33195 14977
rect 20588 14912 20852 14940
rect 20588 14900 20594 14912
rect 21450 14900 21456 14952
rect 21508 14940 21514 14952
rect 21910 14940 21916 14952
rect 21508 14912 21916 14940
rect 21508 14900 21514 14912
rect 21910 14900 21916 14912
rect 21968 14940 21974 14952
rect 22097 14943 22155 14949
rect 22097 14940 22109 14943
rect 21968 14912 22109 14940
rect 21968 14900 21974 14912
rect 22097 14909 22109 14912
rect 22143 14909 22155 14943
rect 23106 14940 23112 14952
rect 23067 14912 23112 14940
rect 22097 14903 22155 14909
rect 23106 14900 23112 14912
rect 23164 14900 23170 14952
rect 24581 14943 24639 14949
rect 24581 14909 24593 14943
rect 24627 14940 24639 14943
rect 24762 14940 24768 14952
rect 24627 14912 24768 14940
rect 24627 14909 24639 14912
rect 24581 14903 24639 14909
rect 24762 14900 24768 14912
rect 24820 14900 24826 14952
rect 24857 14943 24915 14949
rect 24857 14909 24869 14943
rect 24903 14909 24915 14943
rect 27338 14940 27344 14952
rect 27299 14912 27344 14940
rect 24857 14903 24915 14909
rect 24872 14872 24900 14903
rect 27338 14900 27344 14912
rect 27396 14900 27402 14952
rect 28445 14943 28503 14949
rect 28445 14909 28457 14943
rect 28491 14940 28503 14943
rect 29270 14940 29276 14952
rect 28491 14912 29276 14940
rect 28491 14909 28503 14912
rect 28445 14903 28503 14909
rect 29270 14900 29276 14912
rect 29328 14900 29334 14952
rect 25222 14872 25228 14884
rect 11103 14844 16068 14872
rect 16132 14844 25228 14872
rect 11103 14841 11115 14844
rect 11057 14835 11115 14841
rect 1857 14807 1915 14813
rect 1857 14773 1869 14807
rect 1903 14804 1915 14807
rect 2682 14804 2688 14816
rect 1903 14776 2688 14804
rect 1903 14773 1915 14776
rect 1857 14767 1915 14773
rect 2682 14764 2688 14776
rect 2740 14764 2746 14816
rect 3050 14804 3056 14816
rect 3011 14776 3056 14804
rect 3050 14764 3056 14776
rect 3108 14764 3114 14816
rect 3786 14764 3792 14816
rect 3844 14804 3850 14816
rect 3973 14807 4031 14813
rect 3973 14804 3985 14807
rect 3844 14776 3985 14804
rect 3844 14764 3850 14776
rect 3973 14773 3985 14776
rect 4019 14773 4031 14807
rect 5902 14804 5908 14816
rect 5863 14776 5908 14804
rect 3973 14767 4031 14773
rect 5902 14764 5908 14776
rect 5960 14764 5966 14816
rect 8113 14807 8171 14813
rect 8113 14773 8125 14807
rect 8159 14804 8171 14807
rect 15010 14804 15016 14816
rect 8159 14776 15016 14804
rect 8159 14773 8171 14776
rect 8113 14767 8171 14773
rect 15010 14764 15016 14776
rect 15068 14764 15074 14816
rect 15102 14764 15108 14816
rect 15160 14804 15166 14816
rect 16132 14804 16160 14844
rect 25222 14832 25228 14844
rect 25280 14832 25286 14884
rect 15160 14776 16160 14804
rect 16209 14807 16267 14813
rect 15160 14764 15166 14776
rect 16209 14773 16221 14807
rect 16255 14804 16267 14807
rect 16666 14804 16672 14816
rect 16255 14776 16672 14804
rect 16255 14773 16267 14776
rect 16209 14767 16267 14773
rect 16666 14764 16672 14776
rect 16724 14764 16730 14816
rect 17954 14764 17960 14816
rect 18012 14804 18018 14816
rect 19061 14807 19119 14813
rect 19061 14804 19073 14807
rect 18012 14776 19073 14804
rect 18012 14764 18018 14776
rect 19061 14773 19073 14776
rect 19107 14773 19119 14807
rect 19061 14767 19119 14773
rect 19426 14764 19432 14816
rect 19484 14804 19490 14816
rect 20438 14804 20444 14816
rect 19484 14776 20444 14804
rect 19484 14764 19490 14776
rect 20438 14764 20444 14776
rect 20496 14764 20502 14816
rect 21082 14764 21088 14816
rect 21140 14804 21146 14816
rect 22738 14804 22744 14816
rect 21140 14776 22744 14804
rect 21140 14764 21146 14776
rect 22738 14764 22744 14776
rect 22796 14764 22802 14816
rect 23106 14764 23112 14816
rect 23164 14804 23170 14816
rect 26878 14804 26884 14816
rect 23164 14776 26884 14804
rect 23164 14764 23170 14776
rect 26878 14764 26884 14776
rect 26936 14764 26942 14816
rect 27801 14807 27859 14813
rect 27801 14773 27813 14807
rect 27847 14804 27859 14807
rect 28810 14804 28816 14816
rect 27847 14776 28816 14804
rect 27847 14773 27859 14776
rect 27801 14767 27859 14773
rect 28810 14764 28816 14776
rect 28868 14764 28874 14816
rect 29549 14807 29607 14813
rect 29549 14773 29561 14807
rect 29595 14804 29607 14807
rect 29914 14804 29920 14816
rect 29595 14776 29920 14804
rect 29595 14773 29607 14776
rect 29549 14767 29607 14773
rect 29914 14764 29920 14776
rect 29972 14764 29978 14816
rect 31021 14807 31079 14813
rect 31021 14773 31033 14807
rect 31067 14804 31079 14807
rect 31478 14804 31484 14816
rect 31067 14776 31484 14804
rect 31067 14773 31079 14776
rect 31021 14767 31079 14773
rect 31478 14764 31484 14776
rect 31536 14764 31542 14816
rect 32953 14807 33011 14813
rect 32953 14773 32965 14807
rect 32999 14804 33011 14807
rect 34422 14804 34428 14816
rect 32999 14776 34428 14804
rect 32999 14773 33011 14776
rect 32953 14767 33011 14773
rect 34422 14764 34428 14776
rect 34480 14764 34486 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 1581 14603 1639 14609
rect 1581 14569 1593 14603
rect 1627 14600 1639 14603
rect 1854 14600 1860 14612
rect 1627 14572 1860 14600
rect 1627 14569 1639 14572
rect 1581 14563 1639 14569
rect 1854 14560 1860 14572
rect 1912 14560 1918 14612
rect 3050 14600 3056 14612
rect 3011 14572 3056 14600
rect 3050 14560 3056 14572
rect 3108 14560 3114 14612
rect 6273 14603 6331 14609
rect 6273 14569 6285 14603
rect 6319 14600 6331 14603
rect 10594 14600 10600 14612
rect 6319 14572 10600 14600
rect 6319 14569 6331 14572
rect 6273 14563 6331 14569
rect 10594 14560 10600 14572
rect 10652 14560 10658 14612
rect 12805 14603 12863 14609
rect 11164 14572 12388 14600
rect 8386 14532 8392 14544
rect 6104 14504 8392 14532
rect 2682 14464 2688 14476
rect 2643 14436 2688 14464
rect 2682 14424 2688 14436
rect 2740 14424 2746 14476
rect 1762 14396 1768 14408
rect 1723 14368 1768 14396
rect 1762 14356 1768 14368
rect 1820 14356 1826 14408
rect 2498 14396 2504 14408
rect 2459 14368 2504 14396
rect 2498 14356 2504 14368
rect 2556 14356 2562 14408
rect 3973 14399 4031 14405
rect 3973 14365 3985 14399
rect 4019 14396 4031 14399
rect 4706 14396 4712 14408
rect 4019 14368 4712 14396
rect 4019 14365 4031 14368
rect 3973 14359 4031 14365
rect 4706 14356 4712 14368
rect 4764 14356 4770 14408
rect 4890 14396 4896 14408
rect 4851 14368 4896 14396
rect 4890 14356 4896 14368
rect 4948 14356 4954 14408
rect 5537 14399 5595 14405
rect 5537 14365 5549 14399
rect 5583 14396 5595 14399
rect 5626 14396 5632 14408
rect 5583 14368 5632 14396
rect 5583 14365 5595 14368
rect 5537 14359 5595 14365
rect 5626 14356 5632 14368
rect 5684 14356 5690 14408
rect 6104 14396 6132 14504
rect 8386 14492 8392 14504
rect 8444 14492 8450 14544
rect 8478 14492 8484 14544
rect 8536 14532 8542 14544
rect 9582 14532 9588 14544
rect 8536 14504 9588 14532
rect 8536 14492 8542 14504
rect 9582 14492 9588 14504
rect 9640 14532 9646 14544
rect 11164 14532 11192 14572
rect 9640 14504 11192 14532
rect 12360 14532 12388 14572
rect 12805 14569 12817 14603
rect 12851 14600 12863 14603
rect 15746 14600 15752 14612
rect 12851 14572 15752 14600
rect 12851 14569 12863 14572
rect 12805 14563 12863 14569
rect 15746 14560 15752 14572
rect 15804 14600 15810 14612
rect 16850 14600 16856 14612
rect 15804 14572 16856 14600
rect 15804 14560 15810 14572
rect 16850 14560 16856 14572
rect 16908 14560 16914 14612
rect 17034 14560 17040 14612
rect 17092 14600 17098 14612
rect 19426 14600 19432 14612
rect 17092 14572 19432 14600
rect 17092 14560 17098 14572
rect 19426 14560 19432 14572
rect 19484 14560 19490 14612
rect 20530 14600 20536 14612
rect 20491 14572 20536 14600
rect 20530 14560 20536 14572
rect 20588 14560 20594 14612
rect 22002 14600 22008 14612
rect 20640 14572 22008 14600
rect 14274 14532 14280 14544
rect 12360 14504 14280 14532
rect 9640 14492 9646 14504
rect 7834 14464 7840 14476
rect 7795 14436 7840 14464
rect 7834 14424 7840 14436
rect 7892 14424 7898 14476
rect 12342 14464 12348 14476
rect 8588 14436 12348 14464
rect 6181 14399 6239 14405
rect 6181 14396 6193 14399
rect 6104 14368 6193 14396
rect 6181 14365 6193 14368
rect 6227 14365 6239 14399
rect 6181 14359 6239 14365
rect 6270 14356 6276 14408
rect 6328 14396 6334 14408
rect 6454 14396 6460 14408
rect 6328 14368 6460 14396
rect 6328 14356 6334 14368
rect 6454 14356 6460 14368
rect 6512 14396 6518 14408
rect 6825 14399 6883 14405
rect 6825 14396 6837 14399
rect 6512 14368 6837 14396
rect 6512 14356 6518 14368
rect 6825 14365 6837 14368
rect 6871 14365 6883 14399
rect 6825 14359 6883 14365
rect 6917 14399 6975 14405
rect 6917 14365 6929 14399
rect 6963 14396 6975 14399
rect 7374 14396 7380 14408
rect 6963 14368 7380 14396
rect 6963 14365 6975 14368
rect 6917 14359 6975 14365
rect 7374 14356 7380 14368
rect 7432 14356 7438 14408
rect 4985 14331 5043 14337
rect 4985 14297 4997 14331
rect 5031 14328 5043 14331
rect 7098 14328 7104 14340
rect 5031 14300 7104 14328
rect 5031 14297 5043 14300
rect 4985 14291 5043 14297
rect 7098 14288 7104 14300
rect 7156 14288 7162 14340
rect 7558 14328 7564 14340
rect 7519 14300 7564 14328
rect 7558 14288 7564 14300
rect 7616 14288 7622 14340
rect 7650 14288 7656 14340
rect 7708 14328 7714 14340
rect 7708 14300 7753 14328
rect 7708 14288 7714 14300
rect 4065 14263 4123 14269
rect 4065 14229 4077 14263
rect 4111 14260 4123 14263
rect 4706 14260 4712 14272
rect 4111 14232 4712 14260
rect 4111 14229 4123 14232
rect 4065 14223 4123 14229
rect 4706 14220 4712 14232
rect 4764 14220 4770 14272
rect 5626 14260 5632 14272
rect 5587 14232 5632 14260
rect 5626 14220 5632 14232
rect 5684 14220 5690 14272
rect 6914 14220 6920 14272
rect 6972 14260 6978 14272
rect 8588 14260 8616 14436
rect 12342 14424 12348 14436
rect 12400 14424 12406 14476
rect 13556 14473 13584 14504
rect 14274 14492 14280 14504
rect 14332 14492 14338 14544
rect 14458 14492 14464 14544
rect 14516 14532 14522 14544
rect 20640 14532 20668 14572
rect 22002 14560 22008 14572
rect 22060 14560 22066 14612
rect 25516 14572 31754 14600
rect 23198 14532 23204 14544
rect 14516 14504 20668 14532
rect 23159 14504 23204 14532
rect 14516 14492 14522 14504
rect 23198 14492 23204 14504
rect 23256 14492 23262 14544
rect 13541 14467 13599 14473
rect 13541 14433 13553 14467
rect 13587 14433 13599 14467
rect 13541 14427 13599 14433
rect 16025 14467 16083 14473
rect 16025 14433 16037 14467
rect 16071 14464 16083 14467
rect 16114 14464 16120 14476
rect 16071 14436 16120 14464
rect 16071 14433 16083 14436
rect 16025 14427 16083 14433
rect 16114 14424 16120 14436
rect 16172 14424 16178 14476
rect 18230 14424 18236 14476
rect 18288 14464 18294 14476
rect 21453 14467 21511 14473
rect 21453 14464 21465 14467
rect 18288 14436 21465 14464
rect 18288 14424 18294 14436
rect 21453 14433 21465 14436
rect 21499 14464 21511 14467
rect 21818 14464 21824 14476
rect 21499 14436 21824 14464
rect 21499 14433 21511 14436
rect 21453 14427 21511 14433
rect 21818 14424 21824 14436
rect 21876 14424 21882 14476
rect 22097 14467 22155 14473
rect 22097 14433 22109 14467
rect 22143 14464 22155 14467
rect 25406 14464 25412 14476
rect 22143 14436 25412 14464
rect 22143 14433 22155 14436
rect 22097 14427 22155 14433
rect 25406 14424 25412 14436
rect 25464 14424 25470 14476
rect 9125 14399 9183 14405
rect 9125 14365 9137 14399
rect 9171 14396 9183 14399
rect 10226 14396 10232 14408
rect 9171 14368 10232 14396
rect 9171 14365 9183 14368
rect 9125 14359 9183 14365
rect 10226 14356 10232 14368
rect 10284 14356 10290 14408
rect 11054 14396 11060 14408
rect 11015 14368 11060 14396
rect 11054 14356 11060 14368
rect 11112 14356 11118 14408
rect 12618 14356 12624 14408
rect 12676 14396 12682 14408
rect 13265 14399 13323 14405
rect 13265 14396 13277 14399
rect 12676 14368 13277 14396
rect 12676 14356 12682 14368
rect 13265 14365 13277 14368
rect 13311 14396 13323 14399
rect 14277 14399 14335 14405
rect 14277 14396 14289 14399
rect 13311 14368 14289 14396
rect 13311 14365 13323 14368
rect 13265 14359 13323 14365
rect 14277 14365 14289 14368
rect 14323 14396 14335 14399
rect 14918 14396 14924 14408
rect 14323 14368 14924 14396
rect 14323 14365 14335 14368
rect 14277 14359 14335 14365
rect 14918 14356 14924 14368
rect 14976 14356 14982 14408
rect 15286 14396 15292 14408
rect 15247 14368 15292 14396
rect 15286 14356 15292 14368
rect 15344 14356 15350 14408
rect 16942 14356 16948 14408
rect 17000 14396 17006 14408
rect 18049 14399 18107 14405
rect 18049 14396 18061 14399
rect 17000 14368 18061 14396
rect 17000 14356 17006 14368
rect 18049 14365 18061 14368
rect 18095 14396 18107 14399
rect 18693 14399 18751 14405
rect 18693 14396 18705 14399
rect 18095 14368 18705 14396
rect 18095 14365 18107 14368
rect 18049 14359 18107 14365
rect 18693 14365 18705 14368
rect 18739 14396 18751 14399
rect 18966 14396 18972 14408
rect 18739 14368 18972 14396
rect 18739 14365 18751 14368
rect 18693 14359 18751 14365
rect 18966 14356 18972 14368
rect 19024 14396 19030 14408
rect 19797 14399 19855 14405
rect 19797 14396 19809 14399
rect 19024 14368 19809 14396
rect 19024 14356 19030 14368
rect 19797 14365 19809 14368
rect 19843 14365 19855 14399
rect 20438 14396 20444 14408
rect 20399 14368 20444 14396
rect 19797 14359 19855 14365
rect 20438 14356 20444 14368
rect 20496 14356 20502 14408
rect 23566 14356 23572 14408
rect 23624 14396 23630 14408
rect 23753 14399 23811 14405
rect 23753 14396 23765 14399
rect 23624 14368 23765 14396
rect 23624 14356 23630 14368
rect 23753 14365 23765 14368
rect 23799 14365 23811 14399
rect 23753 14359 23811 14365
rect 24302 14356 24308 14408
rect 24360 14396 24366 14408
rect 24581 14399 24639 14405
rect 24581 14396 24593 14399
rect 24360 14368 24593 14396
rect 24360 14356 24366 14368
rect 24581 14365 24593 14368
rect 24627 14396 24639 14399
rect 25516 14396 25544 14572
rect 28813 14535 28871 14541
rect 28813 14532 28825 14535
rect 25700 14504 28825 14532
rect 25700 14476 25728 14504
rect 28813 14501 28825 14504
rect 28859 14501 28871 14535
rect 31726 14532 31754 14572
rect 31726 14504 35894 14532
rect 28813 14495 28871 14501
rect 25682 14464 25688 14476
rect 25595 14436 25688 14464
rect 25682 14424 25688 14436
rect 25740 14424 25746 14476
rect 35866 14464 35894 14504
rect 38194 14464 38200 14476
rect 35866 14436 38200 14464
rect 38194 14424 38200 14436
rect 38252 14424 38258 14476
rect 24627 14368 25544 14396
rect 28721 14399 28779 14405
rect 24627 14365 24639 14368
rect 24581 14359 24639 14365
rect 28721 14365 28733 14399
rect 28767 14365 28779 14399
rect 28721 14359 28779 14365
rect 9214 14288 9220 14340
rect 9272 14328 9278 14340
rect 9861 14331 9919 14337
rect 9861 14328 9873 14331
rect 9272 14300 9873 14328
rect 9272 14288 9278 14300
rect 9861 14297 9873 14300
rect 9907 14297 9919 14331
rect 11330 14328 11336 14340
rect 11291 14300 11336 14328
rect 9861 14291 9919 14297
rect 11330 14288 11336 14300
rect 11388 14288 11394 14340
rect 11440 14300 11822 14328
rect 6972 14232 8616 14260
rect 6972 14220 6978 14232
rect 8754 14220 8760 14272
rect 8812 14260 8818 14272
rect 11440 14260 11468 14300
rect 14366 14288 14372 14340
rect 14424 14328 14430 14340
rect 14553 14331 14611 14337
rect 14553 14328 14565 14331
rect 14424 14300 14565 14328
rect 14424 14288 14430 14300
rect 14553 14297 14565 14300
rect 14599 14297 14611 14331
rect 16117 14331 16175 14337
rect 16117 14328 16129 14331
rect 14553 14291 14611 14297
rect 14660 14300 16129 14328
rect 8812 14232 11468 14260
rect 8812 14220 8818 14232
rect 13078 14220 13084 14272
rect 13136 14260 13142 14272
rect 14660 14260 14688 14300
rect 16117 14297 16129 14300
rect 16163 14297 16175 14331
rect 17034 14328 17040 14340
rect 16995 14300 17040 14328
rect 16117 14291 16175 14297
rect 17034 14288 17040 14300
rect 17092 14288 17098 14340
rect 17770 14288 17776 14340
rect 17828 14328 17834 14340
rect 21266 14328 21272 14340
rect 17828 14300 21272 14328
rect 17828 14288 17834 14300
rect 21266 14288 21272 14300
rect 21324 14288 21330 14340
rect 21542 14288 21548 14340
rect 21600 14328 21606 14340
rect 22646 14328 22652 14340
rect 21600 14300 21645 14328
rect 22607 14300 22652 14328
rect 21600 14288 21606 14300
rect 22646 14288 22652 14300
rect 22704 14288 22710 14340
rect 22741 14331 22799 14337
rect 22741 14297 22753 14331
rect 22787 14297 22799 14331
rect 22741 14291 22799 14297
rect 13136 14232 14688 14260
rect 15381 14263 15439 14269
rect 13136 14220 13142 14232
rect 15381 14229 15393 14263
rect 15427 14260 15439 14263
rect 17310 14260 17316 14272
rect 15427 14232 17316 14260
rect 15427 14229 15439 14232
rect 15381 14223 15439 14229
rect 17310 14220 17316 14232
rect 17368 14220 17374 14272
rect 17586 14220 17592 14272
rect 17644 14260 17650 14272
rect 18141 14263 18199 14269
rect 18141 14260 18153 14263
rect 17644 14232 18153 14260
rect 17644 14220 17650 14232
rect 18141 14229 18153 14232
rect 18187 14229 18199 14263
rect 18141 14223 18199 14229
rect 18322 14220 18328 14272
rect 18380 14260 18386 14272
rect 18785 14263 18843 14269
rect 18785 14260 18797 14263
rect 18380 14232 18797 14260
rect 18380 14220 18386 14232
rect 18785 14229 18797 14232
rect 18831 14229 18843 14263
rect 18785 14223 18843 14229
rect 19150 14220 19156 14272
rect 19208 14260 19214 14272
rect 19889 14263 19947 14269
rect 19889 14260 19901 14263
rect 19208 14232 19901 14260
rect 19208 14220 19214 14232
rect 19889 14229 19901 14232
rect 19935 14229 19947 14263
rect 19889 14223 19947 14229
rect 19978 14220 19984 14272
rect 20036 14260 20042 14272
rect 22756 14260 22784 14291
rect 25774 14288 25780 14340
rect 25832 14328 25838 14340
rect 26697 14331 26755 14337
rect 26697 14328 26709 14331
rect 25832 14300 25877 14328
rect 26252 14300 26709 14328
rect 25832 14288 25838 14300
rect 20036 14232 22784 14260
rect 23845 14263 23903 14269
rect 20036 14220 20042 14232
rect 23845 14229 23857 14263
rect 23891 14260 23903 14263
rect 24302 14260 24308 14272
rect 23891 14232 24308 14260
rect 23891 14229 23903 14232
rect 23845 14223 23903 14229
rect 24302 14220 24308 14232
rect 24360 14220 24366 14272
rect 24670 14260 24676 14272
rect 24631 14232 24676 14260
rect 24670 14220 24676 14232
rect 24728 14220 24734 14272
rect 24762 14220 24768 14272
rect 24820 14260 24826 14272
rect 26252 14260 26280 14300
rect 26697 14297 26709 14300
rect 26743 14297 26755 14331
rect 27246 14328 27252 14340
rect 27207 14300 27252 14328
rect 26697 14291 26755 14297
rect 27246 14288 27252 14300
rect 27304 14288 27310 14340
rect 27341 14331 27399 14337
rect 27341 14297 27353 14331
rect 27387 14297 27399 14331
rect 28258 14328 28264 14340
rect 28219 14300 28264 14328
rect 27341 14291 27399 14297
rect 24820 14232 26280 14260
rect 24820 14220 24826 14232
rect 26326 14220 26332 14272
rect 26384 14260 26390 14272
rect 27356 14260 27384 14291
rect 28258 14288 28264 14300
rect 28316 14288 28322 14340
rect 28736 14328 28764 14359
rect 28810 14356 28816 14408
rect 28868 14396 28874 14408
rect 29733 14399 29791 14405
rect 29733 14396 29745 14399
rect 28868 14368 29745 14396
rect 28868 14356 28874 14368
rect 29733 14365 29745 14368
rect 29779 14365 29791 14399
rect 29733 14359 29791 14365
rect 29825 14399 29883 14405
rect 29825 14365 29837 14399
rect 29871 14396 29883 14399
rect 35069 14399 35127 14405
rect 35069 14396 35081 14399
rect 29871 14368 35081 14396
rect 29871 14365 29883 14368
rect 29825 14359 29883 14365
rect 35069 14365 35081 14368
rect 35115 14365 35127 14399
rect 35069 14359 35127 14365
rect 32582 14328 32588 14340
rect 28736 14300 32588 14328
rect 32582 14288 32588 14300
rect 32640 14288 32646 14340
rect 26384 14232 27384 14260
rect 34885 14263 34943 14269
rect 26384 14220 26390 14232
rect 34885 14229 34897 14263
rect 34931 14260 34943 14263
rect 38010 14260 38016 14272
rect 34931 14232 38016 14260
rect 34931 14229 34943 14232
rect 34885 14223 34943 14229
rect 38010 14220 38016 14232
rect 38068 14220 38074 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 2961 14059 3019 14065
rect 2961 14025 2973 14059
rect 3007 14056 3019 14059
rect 3510 14056 3516 14068
rect 3007 14028 3516 14056
rect 3007 14025 3019 14028
rect 2961 14019 3019 14025
rect 3510 14016 3516 14028
rect 3568 14016 3574 14068
rect 3697 14059 3755 14065
rect 3697 14025 3709 14059
rect 3743 14056 3755 14059
rect 4062 14056 4068 14068
rect 3743 14028 4068 14056
rect 3743 14025 3755 14028
rect 3697 14019 3755 14025
rect 4062 14016 4068 14028
rect 4120 14016 4126 14068
rect 5534 14056 5540 14068
rect 4172 14028 5540 14056
rect 3050 13948 3056 14000
rect 3108 13988 3114 14000
rect 3108 13960 3648 13988
rect 3108 13948 3114 13960
rect 1578 13920 1584 13932
rect 1539 13892 1584 13920
rect 1578 13880 1584 13892
rect 1636 13880 1642 13932
rect 3620 13929 3648 13960
rect 3145 13923 3203 13929
rect 3145 13889 3157 13923
rect 3191 13889 3203 13923
rect 3145 13883 3203 13889
rect 3605 13923 3663 13929
rect 3605 13889 3617 13923
rect 3651 13889 3663 13923
rect 3605 13883 3663 13889
rect 3160 13852 3188 13883
rect 4172 13852 4200 14028
rect 5534 14016 5540 14028
rect 5592 14016 5598 14068
rect 6914 14056 6920 14068
rect 6875 14028 6920 14056
rect 6914 14016 6920 14028
rect 6972 14016 6978 14068
rect 7466 14016 7472 14068
rect 7524 14056 7530 14068
rect 9217 14059 9275 14065
rect 7524 14028 9168 14056
rect 7524 14016 7530 14028
rect 4341 13991 4399 13997
rect 4341 13957 4353 13991
rect 4387 13988 4399 13991
rect 7374 13988 7380 14000
rect 4387 13960 7380 13988
rect 4387 13957 4399 13960
rect 4341 13951 4399 13957
rect 7374 13948 7380 13960
rect 7432 13948 7438 14000
rect 7742 13948 7748 14000
rect 7800 13988 7806 14000
rect 7800 13960 7845 13988
rect 7800 13948 7806 13960
rect 8294 13948 8300 14000
rect 8352 13948 8358 14000
rect 4249 13923 4307 13929
rect 4249 13889 4261 13923
rect 4295 13920 4307 13923
rect 4614 13920 4620 13932
rect 4295 13892 4620 13920
rect 4295 13889 4307 13892
rect 4249 13883 4307 13889
rect 4614 13880 4620 13892
rect 4672 13880 4678 13932
rect 4893 13923 4951 13929
rect 4893 13889 4905 13923
rect 4939 13920 4951 13923
rect 5813 13923 5871 13929
rect 4939 13892 5764 13920
rect 4939 13889 4951 13892
rect 4893 13883 4951 13889
rect 3160 13824 4200 13852
rect 4985 13855 5043 13861
rect 4985 13821 4997 13855
rect 5031 13852 5043 13855
rect 5442 13852 5448 13864
rect 5031 13824 5448 13852
rect 5031 13821 5043 13824
rect 4985 13815 5043 13821
rect 5442 13812 5448 13824
rect 5500 13812 5506 13864
rect 1762 13716 1768 13728
rect 1723 13688 1768 13716
rect 1762 13676 1768 13688
rect 1820 13676 1826 13728
rect 5736 13716 5764 13892
rect 5813 13889 5825 13923
rect 5859 13920 5871 13923
rect 6086 13920 6092 13932
rect 5859 13892 6092 13920
rect 5859 13890 5880 13892
rect 5859 13889 5871 13890
rect 5813 13883 5871 13889
rect 6086 13880 6092 13892
rect 6144 13880 6150 13932
rect 6825 13923 6883 13929
rect 6825 13889 6837 13923
rect 6871 13920 6883 13923
rect 6914 13920 6920 13932
rect 6871 13892 6920 13920
rect 6871 13889 6883 13892
rect 6825 13883 6883 13889
rect 6914 13880 6920 13892
rect 6972 13880 6978 13932
rect 5905 13855 5963 13861
rect 5905 13821 5917 13855
rect 5951 13852 5963 13855
rect 7374 13852 7380 13864
rect 5951 13824 7380 13852
rect 5951 13821 5963 13824
rect 5905 13815 5963 13821
rect 7374 13812 7380 13824
rect 7432 13812 7438 13864
rect 7469 13855 7527 13861
rect 7469 13821 7481 13855
rect 7515 13852 7527 13855
rect 7834 13852 7840 13864
rect 7515 13824 7840 13852
rect 7515 13821 7527 13824
rect 7469 13815 7527 13821
rect 7834 13812 7840 13824
rect 7892 13852 7898 13864
rect 9140 13852 9168 14028
rect 9217 14025 9229 14059
rect 9263 14025 9275 14059
rect 18233 14059 18291 14065
rect 9217 14019 9275 14025
rect 11256 14028 14964 14056
rect 9232 13988 9260 14019
rect 9766 13988 9772 14000
rect 9232 13960 9772 13988
rect 9766 13948 9772 13960
rect 9824 13948 9830 14000
rect 10226 13920 10232 13932
rect 10139 13892 10232 13920
rect 10226 13880 10232 13892
rect 10284 13920 10290 13932
rect 11256 13920 11284 14028
rect 11977 13991 12035 13997
rect 11977 13957 11989 13991
rect 12023 13988 12035 13991
rect 13078 13988 13084 14000
rect 12023 13960 13084 13988
rect 12023 13957 12035 13960
rect 11977 13951 12035 13957
rect 13078 13948 13084 13960
rect 13136 13948 13142 14000
rect 13814 13948 13820 14000
rect 13872 13948 13878 14000
rect 14936 13997 14964 14028
rect 18233 14025 18245 14059
rect 18279 14056 18291 14059
rect 19978 14056 19984 14068
rect 18279 14028 19984 14056
rect 18279 14025 18291 14028
rect 18233 14019 18291 14025
rect 19978 14016 19984 14028
rect 20036 14016 20042 14068
rect 20070 14016 20076 14068
rect 20128 14056 20134 14068
rect 20346 14056 20352 14068
rect 20128 14028 20352 14056
rect 20128 14016 20134 14028
rect 20346 14016 20352 14028
rect 20404 14056 20410 14068
rect 20533 14059 20591 14065
rect 20533 14056 20545 14059
rect 20404 14028 20545 14056
rect 20404 14016 20410 14028
rect 20533 14025 20545 14028
rect 20579 14025 20591 14059
rect 20533 14019 20591 14025
rect 21177 14059 21235 14065
rect 21177 14025 21189 14059
rect 21223 14056 21235 14059
rect 21542 14056 21548 14068
rect 21223 14028 21548 14056
rect 21223 14025 21235 14028
rect 21177 14019 21235 14025
rect 21542 14016 21548 14028
rect 21600 14016 21606 14068
rect 21910 14016 21916 14068
rect 21968 14056 21974 14068
rect 25685 14059 25743 14065
rect 21968 14028 23428 14056
rect 21968 14016 21974 14028
rect 14921 13991 14979 13997
rect 14921 13957 14933 13991
rect 14967 13957 14979 13991
rect 14921 13951 14979 13957
rect 15378 13948 15384 14000
rect 15436 13988 15442 14000
rect 19334 13988 19340 14000
rect 15436 13960 16804 13988
rect 15436 13948 15442 13960
rect 11882 13920 11888 13932
rect 10284 13892 11284 13920
rect 11843 13892 11888 13920
rect 10284 13880 10290 13892
rect 11882 13880 11888 13892
rect 11940 13880 11946 13932
rect 16776 13918 16804 13960
rect 18800 13960 19340 13988
rect 16853 13923 16911 13929
rect 16853 13918 16865 13923
rect 16776 13890 16865 13918
rect 16853 13889 16865 13890
rect 16899 13889 16911 13923
rect 18141 13923 18199 13929
rect 18141 13920 18153 13923
rect 16853 13883 16911 13889
rect 16960 13892 18153 13920
rect 10502 13852 10508 13864
rect 7892 13824 8800 13852
rect 9140 13824 10508 13852
rect 7892 13812 7898 13824
rect 8772 13784 8800 13824
rect 10502 13812 10508 13824
rect 10560 13812 10566 13864
rect 11054 13852 11060 13864
rect 11015 13824 11060 13852
rect 11054 13812 11060 13824
rect 11112 13852 11118 13864
rect 12529 13855 12587 13861
rect 12529 13852 12541 13855
rect 11112 13824 12541 13852
rect 11112 13812 11118 13824
rect 12529 13821 12541 13824
rect 12575 13821 12587 13855
rect 12529 13815 12587 13821
rect 13998 13812 14004 13864
rect 14056 13852 14062 13864
rect 15657 13855 15715 13861
rect 15657 13852 15669 13855
rect 14056 13824 15669 13852
rect 14056 13812 14062 13824
rect 15657 13821 15669 13824
rect 15703 13821 15715 13855
rect 15657 13815 15715 13821
rect 16114 13812 16120 13864
rect 16172 13852 16178 13864
rect 16960 13852 16988 13892
rect 18141 13889 18153 13892
rect 18187 13889 18199 13923
rect 18141 13883 18199 13889
rect 16172 13824 16988 13852
rect 17129 13855 17187 13861
rect 16172 13812 16178 13824
rect 17129 13821 17141 13855
rect 17175 13852 17187 13855
rect 17770 13852 17776 13864
rect 17175 13824 17776 13852
rect 17175 13821 17187 13824
rect 17129 13815 17187 13821
rect 17770 13812 17776 13824
rect 17828 13812 17834 13864
rect 18800 13861 18828 13960
rect 19334 13948 19340 13960
rect 19392 13948 19398 14000
rect 20286 13960 21220 13988
rect 21085 13923 21143 13929
rect 21085 13889 21097 13923
rect 21131 13889 21143 13923
rect 21192 13920 21220 13960
rect 21818 13948 21824 14000
rect 21876 13988 21882 14000
rect 23400 13997 23428 14028
rect 25685 14025 25697 14059
rect 25731 14056 25743 14059
rect 25774 14056 25780 14068
rect 25731 14028 25780 14056
rect 25731 14025 25743 14028
rect 25685 14019 25743 14025
rect 25774 14016 25780 14028
rect 25832 14016 25838 14068
rect 26326 14056 26332 14068
rect 26287 14028 26332 14056
rect 26326 14016 26332 14028
rect 26384 14016 26390 14068
rect 27246 14016 27252 14068
rect 27304 14056 27310 14068
rect 27801 14059 27859 14065
rect 27801 14056 27813 14059
rect 27304 14028 27813 14056
rect 27304 14016 27310 14028
rect 27801 14025 27813 14028
rect 27847 14025 27859 14059
rect 27801 14019 27859 14025
rect 28258 14016 28264 14068
rect 28316 14056 28322 14068
rect 36170 14056 36176 14068
rect 28316 14028 36176 14056
rect 28316 14016 28322 14028
rect 36170 14016 36176 14028
rect 36228 14016 36234 14068
rect 22465 13991 22523 13997
rect 22465 13988 22477 13991
rect 21876 13960 22477 13988
rect 21876 13948 21882 13960
rect 22465 13957 22477 13960
rect 22511 13957 22523 13991
rect 22465 13951 22523 13957
rect 23385 13991 23443 13997
rect 23385 13957 23397 13991
rect 23431 13957 23443 13991
rect 23385 13951 23443 13957
rect 24026 13948 24032 14000
rect 24084 13988 24090 14000
rect 24084 13960 24129 13988
rect 24084 13948 24090 13960
rect 24578 13948 24584 14000
rect 24636 13988 24642 14000
rect 24762 13988 24768 14000
rect 24636 13960 24768 13988
rect 24636 13948 24642 13960
rect 24762 13948 24768 13960
rect 24820 13988 24826 14000
rect 24949 13991 25007 13997
rect 24949 13988 24961 13991
rect 24820 13960 24961 13988
rect 24820 13948 24826 13960
rect 24949 13957 24961 13960
rect 24995 13957 25007 13991
rect 24949 13951 25007 13957
rect 22094 13920 22100 13932
rect 21192 13892 22100 13920
rect 21085 13883 21143 13889
rect 18785 13855 18843 13861
rect 18785 13852 18797 13855
rect 17972 13824 18797 13852
rect 9214 13784 9220 13796
rect 8772 13756 9220 13784
rect 9214 13744 9220 13756
rect 9272 13744 9278 13796
rect 9766 13744 9772 13796
rect 9824 13784 9830 13796
rect 11238 13784 11244 13796
rect 9824 13756 11244 13784
rect 9824 13744 9830 13756
rect 11238 13744 11244 13756
rect 11296 13784 11302 13796
rect 11296 13756 12664 13784
rect 11296 13744 11302 13756
rect 6178 13716 6184 13728
rect 5736 13688 6184 13716
rect 6178 13676 6184 13688
rect 6236 13716 6242 13728
rect 6730 13716 6736 13728
rect 6236 13688 6736 13716
rect 6236 13676 6242 13688
rect 6730 13676 6736 13688
rect 6788 13676 6794 13728
rect 6914 13676 6920 13728
rect 6972 13716 6978 13728
rect 7190 13716 7196 13728
rect 6972 13688 7196 13716
rect 6972 13676 6978 13688
rect 7190 13676 7196 13688
rect 7248 13676 7254 13728
rect 7742 13676 7748 13728
rect 7800 13716 7806 13728
rect 8202 13716 8208 13728
rect 7800 13688 8208 13716
rect 7800 13676 7806 13688
rect 8202 13676 8208 13688
rect 8260 13676 8266 13728
rect 8478 13676 8484 13728
rect 8536 13716 8542 13728
rect 12342 13716 12348 13728
rect 8536 13688 12348 13716
rect 8536 13676 8542 13688
rect 12342 13676 12348 13688
rect 12400 13676 12406 13728
rect 12636 13716 12664 13756
rect 16574 13744 16580 13796
rect 16632 13784 16638 13796
rect 17972 13784 18000 13824
rect 18785 13821 18797 13824
rect 18831 13821 18843 13855
rect 19061 13855 19119 13861
rect 19061 13852 19073 13855
rect 18785 13815 18843 13821
rect 18892 13824 19073 13852
rect 16632 13756 18000 13784
rect 16632 13744 16638 13756
rect 18414 13744 18420 13796
rect 18472 13784 18478 13796
rect 18892 13784 18920 13824
rect 19061 13821 19073 13824
rect 19107 13852 19119 13855
rect 20530 13852 20536 13864
rect 19107 13824 20536 13852
rect 19107 13821 19119 13824
rect 19061 13815 19119 13821
rect 20530 13812 20536 13824
rect 20588 13812 20594 13864
rect 21100 13852 21128 13883
rect 22094 13880 22100 13892
rect 22152 13880 22158 13932
rect 25590 13920 25596 13932
rect 25551 13892 25596 13920
rect 25590 13880 25596 13892
rect 25648 13880 25654 13932
rect 25866 13880 25872 13932
rect 25924 13920 25930 13932
rect 26237 13923 26295 13929
rect 26237 13920 26249 13923
rect 25924 13892 26249 13920
rect 25924 13880 25930 13892
rect 26237 13889 26249 13892
rect 26283 13889 26295 13923
rect 27154 13920 27160 13932
rect 27115 13892 27160 13920
rect 26237 13883 26295 13889
rect 27154 13880 27160 13892
rect 27212 13880 27218 13932
rect 27249 13923 27307 13929
rect 27249 13889 27261 13923
rect 27295 13920 27307 13923
rect 27338 13920 27344 13932
rect 27295 13892 27344 13920
rect 27295 13889 27307 13892
rect 27249 13883 27307 13889
rect 27338 13880 27344 13892
rect 27396 13880 27402 13932
rect 28721 13923 28779 13929
rect 28721 13889 28733 13923
rect 28767 13920 28779 13923
rect 29825 13923 29883 13929
rect 29825 13920 29837 13923
rect 28767 13892 29837 13920
rect 28767 13889 28779 13892
rect 28721 13883 28779 13889
rect 29825 13889 29837 13892
rect 29871 13889 29883 13923
rect 31478 13920 31484 13932
rect 31439 13892 31484 13920
rect 29825 13883 29883 13889
rect 31478 13880 31484 13892
rect 31536 13880 31542 13932
rect 38010 13920 38016 13932
rect 37971 13892 38016 13920
rect 38010 13880 38016 13892
rect 38068 13880 38074 13932
rect 22373 13855 22431 13861
rect 21100 13824 22094 13852
rect 20990 13784 20996 13796
rect 18472 13756 18920 13784
rect 20088 13756 20996 13784
rect 18472 13744 18478 13756
rect 12786 13719 12844 13725
rect 12786 13716 12798 13719
rect 12636 13688 12798 13716
rect 12786 13685 12798 13688
rect 12832 13685 12844 13719
rect 12786 13679 12844 13685
rect 14090 13676 14096 13728
rect 14148 13716 14154 13728
rect 14277 13719 14335 13725
rect 14277 13716 14289 13719
rect 14148 13688 14289 13716
rect 14148 13676 14154 13688
rect 14277 13685 14289 13688
rect 14323 13716 14335 13719
rect 14458 13716 14464 13728
rect 14323 13688 14464 13716
rect 14323 13685 14335 13688
rect 14277 13679 14335 13685
rect 14458 13676 14464 13688
rect 14516 13676 14522 13728
rect 17218 13676 17224 13728
rect 17276 13716 17282 13728
rect 20088 13716 20116 13756
rect 20990 13744 20996 13756
rect 21048 13784 21054 13796
rect 21910 13784 21916 13796
rect 21048 13756 21916 13784
rect 21048 13744 21054 13756
rect 21910 13744 21916 13756
rect 21968 13744 21974 13796
rect 22066 13784 22094 13824
rect 22373 13821 22385 13855
rect 22419 13852 22431 13855
rect 22419 13824 23336 13852
rect 22419 13821 22431 13824
rect 22373 13815 22431 13821
rect 22922 13784 22928 13796
rect 22066 13756 22928 13784
rect 22922 13744 22928 13756
rect 22980 13744 22986 13796
rect 23308 13784 23336 13824
rect 23382 13812 23388 13864
rect 23440 13852 23446 13864
rect 23937 13855 23995 13861
rect 23937 13852 23949 13855
rect 23440 13824 23949 13852
rect 23440 13812 23446 13824
rect 23937 13821 23949 13824
rect 23983 13821 23995 13855
rect 23937 13815 23995 13821
rect 28905 13855 28963 13861
rect 28905 13821 28917 13855
rect 28951 13852 28963 13855
rect 29730 13852 29736 13864
rect 28951 13824 29736 13852
rect 28951 13821 28963 13824
rect 28905 13815 28963 13821
rect 29730 13812 29736 13824
rect 29788 13812 29794 13864
rect 25958 13784 25964 13796
rect 23308 13756 25964 13784
rect 25958 13744 25964 13756
rect 26016 13744 26022 13796
rect 17276 13688 20116 13716
rect 17276 13676 17282 13688
rect 20346 13676 20352 13728
rect 20404 13716 20410 13728
rect 21450 13716 21456 13728
rect 20404 13688 21456 13716
rect 20404 13676 20410 13688
rect 21450 13676 21456 13688
rect 21508 13676 21514 13728
rect 27614 13676 27620 13728
rect 27672 13716 27678 13728
rect 28442 13716 28448 13728
rect 27672 13688 28448 13716
rect 27672 13676 27678 13688
rect 28442 13676 28448 13688
rect 28500 13716 28506 13728
rect 29089 13719 29147 13725
rect 29089 13716 29101 13719
rect 28500 13688 29101 13716
rect 28500 13676 28506 13688
rect 29089 13685 29101 13688
rect 29135 13685 29147 13719
rect 31294 13716 31300 13728
rect 31255 13688 31300 13716
rect 29089 13679 29147 13685
rect 31294 13676 31300 13688
rect 31352 13676 31358 13728
rect 38194 13716 38200 13728
rect 38155 13688 38200 13716
rect 38194 13676 38200 13688
rect 38252 13676 38258 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 5902 13472 5908 13524
rect 5960 13512 5966 13524
rect 8294 13512 8300 13524
rect 5960 13484 8300 13512
rect 5960 13472 5966 13484
rect 8294 13472 8300 13484
rect 8352 13472 8358 13524
rect 9122 13472 9128 13524
rect 9180 13512 9186 13524
rect 9180 13484 10732 13512
rect 9180 13472 9186 13484
rect 8573 13447 8631 13453
rect 8573 13413 8585 13447
rect 8619 13444 8631 13447
rect 8619 13416 9260 13444
rect 8619 13413 8631 13416
rect 8573 13407 8631 13413
rect 4614 13336 4620 13388
rect 4672 13376 4678 13388
rect 5258 13376 5264 13388
rect 4672 13348 5264 13376
rect 4672 13336 4678 13348
rect 5258 13336 5264 13348
rect 5316 13336 5322 13388
rect 6730 13336 6736 13388
rect 6788 13376 6794 13388
rect 6825 13379 6883 13385
rect 6825 13376 6837 13379
rect 6788 13348 6837 13376
rect 6788 13336 6794 13348
rect 6825 13345 6837 13348
rect 6871 13376 6883 13379
rect 7834 13376 7840 13388
rect 6871 13348 7840 13376
rect 6871 13345 6883 13348
rect 6825 13339 6883 13345
rect 7834 13336 7840 13348
rect 7892 13336 7898 13388
rect 8294 13336 8300 13388
rect 8352 13336 8358 13388
rect 9122 13376 9128 13388
rect 9083 13348 9128 13376
rect 9122 13336 9128 13348
rect 9180 13336 9186 13388
rect 9232 13376 9260 13416
rect 9766 13376 9772 13388
rect 9232 13348 9772 13376
rect 9766 13336 9772 13348
rect 9824 13336 9830 13388
rect 4706 13308 4712 13320
rect 4667 13280 4712 13308
rect 4706 13268 4712 13280
rect 4764 13268 4770 13320
rect 5169 13311 5227 13317
rect 5169 13277 5181 13311
rect 5215 13308 5227 13311
rect 5276 13308 5304 13336
rect 5810 13308 5816 13320
rect 5215 13280 5304 13308
rect 5771 13280 5816 13308
rect 5215 13277 5227 13280
rect 5169 13271 5227 13277
rect 5810 13268 5816 13280
rect 5868 13268 5874 13320
rect 5905 13311 5963 13317
rect 5905 13277 5917 13311
rect 5951 13308 5963 13311
rect 8312 13308 8340 13336
rect 5951 13280 6868 13308
rect 8312 13280 8432 13308
rect 5951 13277 5963 13280
rect 5905 13271 5963 13277
rect 5261 13243 5319 13249
rect 5261 13209 5273 13243
rect 5307 13209 5319 13243
rect 6840 13240 6868 13280
rect 7006 13240 7012 13252
rect 6840 13212 7012 13240
rect 5261 13203 5319 13209
rect 4525 13175 4583 13181
rect 4525 13141 4537 13175
rect 4571 13172 4583 13175
rect 4614 13172 4620 13184
rect 4571 13144 4620 13172
rect 4571 13141 4583 13144
rect 4525 13135 4583 13141
rect 4614 13132 4620 13144
rect 4672 13132 4678 13184
rect 4706 13132 4712 13184
rect 4764 13172 4770 13184
rect 4890 13172 4896 13184
rect 4764 13144 4896 13172
rect 4764 13132 4770 13144
rect 4890 13132 4896 13144
rect 4948 13132 4954 13184
rect 5276 13172 5304 13203
rect 7006 13200 7012 13212
rect 7064 13200 7070 13252
rect 7101 13243 7159 13249
rect 7101 13209 7113 13243
rect 7147 13240 7159 13243
rect 7190 13240 7196 13252
rect 7147 13212 7196 13240
rect 7147 13209 7159 13212
rect 7101 13203 7159 13209
rect 7190 13200 7196 13212
rect 7248 13200 7254 13252
rect 8404 13240 8432 13280
rect 7300 13212 7590 13240
rect 8404 13212 9260 13240
rect 7300 13172 7328 13212
rect 5276 13144 7328 13172
rect 7466 13132 7472 13184
rect 7524 13172 7530 13184
rect 8478 13172 8484 13184
rect 7524 13144 8484 13172
rect 7524 13132 7530 13144
rect 8478 13132 8484 13144
rect 8536 13132 8542 13184
rect 9232 13172 9260 13212
rect 9306 13200 9312 13252
rect 9364 13240 9370 13252
rect 9401 13243 9459 13249
rect 9401 13240 9413 13243
rect 9364 13212 9413 13240
rect 9364 13200 9370 13212
rect 9401 13209 9413 13212
rect 9447 13209 9459 13243
rect 10704 13240 10732 13484
rect 12526 13472 12532 13524
rect 12584 13512 12590 13524
rect 15194 13512 15200 13524
rect 12584 13484 15200 13512
rect 12584 13472 12590 13484
rect 15194 13472 15200 13484
rect 15252 13472 15258 13524
rect 17034 13472 17040 13524
rect 17092 13512 17098 13524
rect 17494 13512 17500 13524
rect 17092 13484 17500 13512
rect 17092 13472 17098 13484
rect 17494 13472 17500 13484
rect 17552 13472 17558 13524
rect 18230 13472 18236 13524
rect 18288 13512 18294 13524
rect 18325 13515 18383 13521
rect 18325 13512 18337 13515
rect 18288 13484 18337 13512
rect 18288 13472 18294 13484
rect 18325 13481 18337 13484
rect 18371 13512 18383 13515
rect 19702 13512 19708 13524
rect 18371 13484 19708 13512
rect 18371 13481 18383 13484
rect 18325 13475 18383 13481
rect 19702 13472 19708 13484
rect 19760 13472 19766 13524
rect 21818 13512 21824 13524
rect 21779 13484 21824 13512
rect 21818 13472 21824 13484
rect 21876 13472 21882 13524
rect 26694 13512 26700 13524
rect 22112 13484 26700 13512
rect 13630 13444 13636 13456
rect 13591 13416 13636 13444
rect 13630 13404 13636 13416
rect 13688 13404 13694 13456
rect 10873 13379 10931 13385
rect 10873 13345 10885 13379
rect 10919 13376 10931 13379
rect 12158 13376 12164 13388
rect 10919 13348 12164 13376
rect 10919 13345 10931 13348
rect 10873 13339 10931 13345
rect 12158 13336 12164 13348
rect 12216 13336 12222 13388
rect 12710 13336 12716 13388
rect 12768 13376 12774 13388
rect 13722 13376 13728 13388
rect 12768 13348 13728 13376
rect 12768 13336 12774 13348
rect 13722 13336 13728 13348
rect 13780 13336 13786 13388
rect 14550 13376 14556 13388
rect 14511 13348 14556 13376
rect 14550 13336 14556 13348
rect 14608 13376 14614 13388
rect 14918 13376 14924 13388
rect 14608 13348 14924 13376
rect 14608 13336 14614 13348
rect 14918 13336 14924 13348
rect 14976 13336 14982 13388
rect 21082 13376 21088 13388
rect 15948 13348 21088 13376
rect 11882 13308 11888 13320
rect 11843 13280 11888 13308
rect 11882 13268 11888 13280
rect 11940 13268 11946 13320
rect 13998 13268 14004 13320
rect 14056 13308 14062 13320
rect 14277 13311 14335 13317
rect 14277 13308 14289 13311
rect 14056 13280 14289 13308
rect 14056 13268 14062 13280
rect 14277 13277 14289 13280
rect 14323 13277 14335 13311
rect 14277 13271 14335 13277
rect 9401 13203 9459 13209
rect 9646 13212 9890 13240
rect 10704 13212 12650 13240
rect 9646 13172 9674 13212
rect 15010 13200 15016 13252
rect 15068 13200 15074 13252
rect 9232 13144 9674 13172
rect 14090 13132 14096 13184
rect 14148 13172 14154 13184
rect 15948 13172 15976 13348
rect 21082 13336 21088 13348
rect 21140 13376 21146 13388
rect 21177 13379 21235 13385
rect 21177 13376 21189 13379
rect 21140 13348 21189 13376
rect 21140 13336 21146 13348
rect 21177 13345 21189 13348
rect 21223 13345 21235 13379
rect 21177 13339 21235 13345
rect 16574 13308 16580 13320
rect 16535 13280 16580 13308
rect 16574 13268 16580 13280
rect 16632 13268 16638 13320
rect 19334 13268 19340 13320
rect 19392 13308 19398 13320
rect 19429 13311 19487 13317
rect 19429 13308 19441 13311
rect 19392 13280 19441 13308
rect 19392 13268 19398 13280
rect 19429 13277 19441 13280
rect 19475 13277 19487 13311
rect 19429 13271 19487 13277
rect 21634 13268 21640 13320
rect 21692 13308 21698 13320
rect 21729 13311 21787 13317
rect 21729 13308 21741 13311
rect 21692 13280 21741 13308
rect 21692 13268 21698 13280
rect 21729 13277 21741 13280
rect 21775 13277 21787 13311
rect 21729 13271 21787 13277
rect 16850 13240 16856 13252
rect 16811 13212 16856 13240
rect 16850 13200 16856 13212
rect 16908 13200 16914 13252
rect 17310 13200 17316 13252
rect 17368 13200 17374 13252
rect 19702 13240 19708 13252
rect 19663 13212 19708 13240
rect 19702 13200 19708 13212
rect 19760 13200 19766 13252
rect 21818 13240 21824 13252
rect 20930 13212 21824 13240
rect 21818 13200 21824 13212
rect 21876 13200 21882 13252
rect 14148 13144 15976 13172
rect 16025 13175 16083 13181
rect 14148 13132 14154 13144
rect 16025 13141 16037 13175
rect 16071 13172 16083 13175
rect 16298 13172 16304 13184
rect 16071 13144 16304 13172
rect 16071 13141 16083 13144
rect 16025 13135 16083 13141
rect 16298 13132 16304 13144
rect 16356 13172 16362 13184
rect 22112 13172 22140 13484
rect 26694 13472 26700 13484
rect 26752 13472 26758 13524
rect 27341 13515 27399 13521
rect 27341 13481 27353 13515
rect 27387 13512 27399 13515
rect 27614 13512 27620 13524
rect 27387 13484 27620 13512
rect 27387 13481 27399 13484
rect 27341 13475 27399 13481
rect 27614 13472 27620 13484
rect 27672 13472 27678 13524
rect 29730 13512 29736 13524
rect 29691 13484 29736 13512
rect 29730 13472 29736 13484
rect 29788 13472 29794 13524
rect 22830 13404 22836 13456
rect 22888 13444 22894 13456
rect 22888 13416 23520 13444
rect 22888 13404 22894 13416
rect 23201 13379 23259 13385
rect 23201 13345 23213 13379
rect 23247 13376 23259 13379
rect 23290 13376 23296 13388
rect 23247 13348 23296 13376
rect 23247 13345 23259 13348
rect 23201 13339 23259 13345
rect 23290 13336 23296 13348
rect 23348 13336 23354 13388
rect 23492 13385 23520 13416
rect 24394 13404 24400 13456
rect 24452 13444 24458 13456
rect 24452 13416 24992 13444
rect 24452 13404 24458 13416
rect 23477 13379 23535 13385
rect 23477 13345 23489 13379
rect 23523 13345 23535 13379
rect 24670 13376 24676 13388
rect 24631 13348 24676 13376
rect 23477 13339 23535 13345
rect 24670 13336 24676 13348
rect 24728 13336 24734 13388
rect 24964 13385 24992 13416
rect 27430 13404 27436 13456
rect 27488 13444 27494 13456
rect 27488 13416 28580 13444
rect 27488 13404 27494 13416
rect 28552 13385 28580 13416
rect 24949 13379 25007 13385
rect 24949 13345 24961 13379
rect 24995 13345 25007 13379
rect 24949 13339 25007 13345
rect 26881 13379 26939 13385
rect 26881 13345 26893 13379
rect 26927 13376 26939 13379
rect 27893 13379 27951 13385
rect 27893 13376 27905 13379
rect 26927 13348 27905 13376
rect 26927 13345 26939 13348
rect 26881 13339 26939 13345
rect 27893 13345 27905 13348
rect 27939 13345 27951 13379
rect 27893 13339 27951 13345
rect 28537 13379 28595 13385
rect 28537 13345 28549 13379
rect 28583 13376 28595 13379
rect 30834 13376 30840 13388
rect 28583 13348 30840 13376
rect 28583 13345 28595 13348
rect 28537 13339 28595 13345
rect 30834 13336 30840 13348
rect 30892 13336 30898 13388
rect 22373 13311 22431 13317
rect 22373 13277 22385 13311
rect 22419 13308 22431 13311
rect 22922 13308 22928 13320
rect 22419 13280 22928 13308
rect 22419 13277 22431 13280
rect 22373 13271 22431 13277
rect 22922 13268 22928 13280
rect 22980 13268 22986 13320
rect 26697 13311 26755 13317
rect 26697 13277 26709 13311
rect 26743 13308 26755 13311
rect 27614 13308 27620 13320
rect 26743 13280 27620 13308
rect 26743 13277 26755 13280
rect 26697 13271 26755 13277
rect 27614 13268 27620 13280
rect 27672 13268 27678 13320
rect 27801 13311 27859 13317
rect 27801 13277 27813 13311
rect 27847 13277 27859 13311
rect 27801 13271 27859 13277
rect 28721 13311 28779 13317
rect 28721 13277 28733 13311
rect 28767 13308 28779 13311
rect 29178 13308 29184 13320
rect 28767 13280 29184 13308
rect 28767 13277 28779 13280
rect 28721 13271 28779 13277
rect 23293 13243 23351 13249
rect 23293 13209 23305 13243
rect 23339 13209 23351 13243
rect 23293 13203 23351 13209
rect 16356 13144 22140 13172
rect 22465 13175 22523 13181
rect 16356 13132 16362 13144
rect 22465 13141 22477 13175
rect 22511 13172 22523 13175
rect 23308 13172 23336 13203
rect 24486 13200 24492 13252
rect 24544 13240 24550 13252
rect 24765 13243 24823 13249
rect 24765 13240 24777 13243
rect 24544 13212 24777 13240
rect 24544 13200 24550 13212
rect 24765 13209 24777 13212
rect 24811 13209 24823 13243
rect 24765 13203 24823 13209
rect 27816 13240 27844 13271
rect 29178 13268 29184 13280
rect 29236 13268 29242 13320
rect 29914 13308 29920 13320
rect 29875 13280 29920 13308
rect 29914 13268 29920 13280
rect 29972 13268 29978 13320
rect 29086 13240 29092 13252
rect 27816 13212 29092 13240
rect 22511 13144 23336 13172
rect 22511 13141 22523 13144
rect 22465 13135 22523 13141
rect 23934 13132 23940 13184
rect 23992 13172 23998 13184
rect 27816 13172 27844 13212
rect 29086 13200 29092 13212
rect 29144 13200 29150 13252
rect 23992 13144 27844 13172
rect 29181 13175 29239 13181
rect 23992 13132 23998 13144
rect 29181 13141 29193 13175
rect 29227 13172 29239 13175
rect 29362 13172 29368 13184
rect 29227 13144 29368 13172
rect 29227 13141 29239 13144
rect 29181 13135 29239 13141
rect 29362 13132 29368 13144
rect 29420 13132 29426 13184
rect 30650 13132 30656 13184
rect 30708 13172 30714 13184
rect 30745 13175 30803 13181
rect 30745 13172 30757 13175
rect 30708 13144 30757 13172
rect 30708 13132 30714 13144
rect 30745 13141 30757 13144
rect 30791 13141 30803 13175
rect 30745 13135 30803 13141
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 3970 12928 3976 12980
rect 4028 12968 4034 12980
rect 4065 12971 4123 12977
rect 4065 12968 4077 12971
rect 4028 12940 4077 12968
rect 4028 12928 4034 12940
rect 4065 12937 4077 12940
rect 4111 12937 4123 12971
rect 4065 12931 4123 12937
rect 5905 12971 5963 12977
rect 5905 12937 5917 12971
rect 5951 12968 5963 12971
rect 8754 12968 8760 12980
rect 5951 12940 8760 12968
rect 5951 12937 5963 12940
rect 5905 12931 5963 12937
rect 8754 12928 8760 12940
rect 8812 12928 8818 12980
rect 9030 12928 9036 12980
rect 9088 12968 9094 12980
rect 9306 12968 9312 12980
rect 9088 12940 9312 12968
rect 9088 12928 9094 12940
rect 9306 12928 9312 12940
rect 9364 12928 9370 12980
rect 11606 12968 11612 12980
rect 10244 12940 11612 12968
rect 3234 12860 3240 12912
rect 3292 12900 3298 12912
rect 3292 12872 6868 12900
rect 3292 12860 3298 12872
rect 6840 12844 6868 12872
rect 7374 12860 7380 12912
rect 7432 12900 7438 12912
rect 10244 12900 10272 12940
rect 11606 12928 11612 12940
rect 11664 12928 11670 12980
rect 11974 12928 11980 12980
rect 12032 12968 12038 12980
rect 13998 12968 14004 12980
rect 12032 12940 14004 12968
rect 12032 12928 12038 12940
rect 13998 12928 14004 12940
rect 14056 12928 14062 12980
rect 14734 12928 14740 12980
rect 14792 12968 14798 12980
rect 15010 12968 15016 12980
rect 14792 12940 15016 12968
rect 14792 12928 14798 12940
rect 15010 12928 15016 12940
rect 15068 12928 15074 12980
rect 15378 12928 15384 12980
rect 15436 12968 15442 12980
rect 16206 12968 16212 12980
rect 15436 12940 16068 12968
rect 16167 12940 16212 12968
rect 15436 12928 15442 12940
rect 7432 12872 8510 12900
rect 10152 12872 10272 12900
rect 11348 12872 12834 12900
rect 7432 12860 7438 12872
rect 1581 12835 1639 12841
rect 1581 12801 1593 12835
rect 1627 12801 1639 12835
rect 1581 12795 1639 12801
rect 1596 12764 1624 12795
rect 1854 12792 1860 12844
rect 1912 12832 1918 12844
rect 3973 12835 4031 12841
rect 3973 12832 3985 12835
rect 1912 12804 3985 12832
rect 1912 12792 1918 12804
rect 3973 12801 3985 12804
rect 4019 12801 4031 12835
rect 3973 12795 4031 12801
rect 5074 12792 5080 12844
rect 5132 12832 5138 12844
rect 5169 12835 5227 12841
rect 5169 12832 5181 12835
rect 5132 12804 5181 12832
rect 5132 12792 5138 12804
rect 5169 12801 5181 12804
rect 5215 12801 5227 12835
rect 5169 12795 5227 12801
rect 5813 12835 5871 12841
rect 5813 12801 5825 12835
rect 5859 12832 5871 12835
rect 5902 12832 5908 12844
rect 5859 12804 5908 12832
rect 5859 12801 5871 12804
rect 5813 12795 5871 12801
rect 5902 12792 5908 12804
rect 5960 12832 5966 12844
rect 6178 12832 6184 12844
rect 5960 12804 6184 12832
rect 5960 12792 5966 12804
rect 6178 12792 6184 12804
rect 6236 12792 6242 12844
rect 6822 12792 6828 12844
rect 6880 12832 6886 12844
rect 7101 12835 7159 12841
rect 7101 12832 7113 12835
rect 6880 12804 7113 12832
rect 6880 12792 6886 12804
rect 7101 12801 7113 12804
rect 7147 12801 7159 12835
rect 7101 12795 7159 12801
rect 7190 12792 7196 12844
rect 7248 12832 7254 12844
rect 7742 12832 7748 12844
rect 7248 12804 7604 12832
rect 7703 12804 7748 12832
rect 7248 12792 7254 12804
rect 5261 12767 5319 12773
rect 1596 12736 2774 12764
rect 2746 12696 2774 12736
rect 5261 12733 5273 12767
rect 5307 12764 5319 12767
rect 7466 12764 7472 12776
rect 5307 12736 7472 12764
rect 5307 12733 5319 12736
rect 5261 12727 5319 12733
rect 7466 12724 7472 12736
rect 7524 12724 7530 12776
rect 7576 12764 7604 12804
rect 7742 12792 7748 12804
rect 7800 12792 7806 12844
rect 10152 12841 10180 12872
rect 10137 12835 10195 12841
rect 10137 12801 10149 12835
rect 10183 12801 10195 12835
rect 10137 12795 10195 12801
rect 7650 12764 7656 12776
rect 7576 12736 7656 12764
rect 7650 12724 7656 12736
rect 7708 12724 7714 12776
rect 8021 12767 8079 12773
rect 8021 12733 8033 12767
rect 8067 12764 8079 12767
rect 9766 12764 9772 12776
rect 8067 12736 9772 12764
rect 8067 12733 8079 12736
rect 8021 12727 8079 12733
rect 9766 12724 9772 12736
rect 9824 12724 9830 12776
rect 10318 12724 10324 12776
rect 10376 12764 10382 12776
rect 10376 12736 10421 12764
rect 10376 12724 10382 12736
rect 6914 12696 6920 12708
rect 2746 12668 6920 12696
rect 6914 12656 6920 12668
rect 6972 12656 6978 12708
rect 7374 12696 7380 12708
rect 7116 12668 7380 12696
rect 1762 12628 1768 12640
rect 1723 12600 1768 12628
rect 1762 12588 1768 12600
rect 1820 12588 1826 12640
rect 3602 12588 3608 12640
rect 3660 12628 3666 12640
rect 3970 12628 3976 12640
rect 3660 12600 3976 12628
rect 3660 12588 3666 12600
rect 3970 12588 3976 12600
rect 4028 12588 4034 12640
rect 4706 12588 4712 12640
rect 4764 12628 4770 12640
rect 7116 12628 7144 12668
rect 7374 12656 7380 12668
rect 7432 12656 7438 12708
rect 9030 12656 9036 12708
rect 9088 12696 9094 12708
rect 9214 12696 9220 12708
rect 9088 12668 9220 12696
rect 9088 12656 9094 12668
rect 9214 12656 9220 12668
rect 9272 12656 9278 12708
rect 11348 12696 11376 12872
rect 13814 12860 13820 12912
rect 13872 12900 13878 12912
rect 16040 12900 16068 12940
rect 16206 12928 16212 12940
rect 16264 12928 16270 12980
rect 19518 12968 19524 12980
rect 17052 12940 19524 12968
rect 17052 12900 17080 12940
rect 19518 12928 19524 12940
rect 19576 12968 19582 12980
rect 19978 12968 19984 12980
rect 19576 12940 19984 12968
rect 19576 12928 19582 12940
rect 19978 12928 19984 12940
rect 20036 12928 20042 12980
rect 22465 12971 22523 12977
rect 22465 12968 22477 12971
rect 20088 12940 22477 12968
rect 13872 12872 15226 12900
rect 16040 12872 17080 12900
rect 17129 12903 17187 12909
rect 13872 12860 13878 12872
rect 17129 12869 17141 12903
rect 17175 12900 17187 12903
rect 17218 12900 17224 12912
rect 17175 12872 17224 12900
rect 17175 12869 17187 12872
rect 17129 12863 17187 12869
rect 17218 12860 17224 12872
rect 17276 12860 17282 12912
rect 20088 12900 20116 12940
rect 22465 12937 22477 12940
rect 22511 12937 22523 12971
rect 22465 12931 22523 12937
rect 22646 12928 22652 12980
rect 22704 12968 22710 12980
rect 23109 12971 23167 12977
rect 23109 12968 23121 12971
rect 22704 12940 23121 12968
rect 22704 12928 22710 12940
rect 23109 12937 23121 12940
rect 23155 12937 23167 12971
rect 26234 12968 26240 12980
rect 23109 12931 23167 12937
rect 24044 12940 26240 12968
rect 23842 12900 23848 12912
rect 18354 12872 20116 12900
rect 20930 12872 23848 12900
rect 23842 12860 23848 12872
rect 23900 12860 23906 12912
rect 11974 12792 11980 12844
rect 12032 12832 12038 12844
rect 12069 12835 12127 12841
rect 12069 12832 12081 12835
rect 12032 12804 12081 12832
rect 12032 12792 12038 12804
rect 12069 12801 12081 12804
rect 12115 12801 12127 12835
rect 12069 12795 12127 12801
rect 13998 12792 14004 12844
rect 14056 12832 14062 12844
rect 14461 12835 14519 12841
rect 14461 12832 14473 12835
rect 14056 12804 14473 12832
rect 14056 12792 14062 12804
rect 14461 12801 14473 12804
rect 14507 12801 14519 12835
rect 14461 12795 14519 12801
rect 19334 12792 19340 12844
rect 19392 12832 19398 12844
rect 19429 12835 19487 12841
rect 19429 12832 19441 12835
rect 19392 12804 19441 12832
rect 19392 12792 19398 12804
rect 19429 12801 19441 12804
rect 19475 12801 19487 12835
rect 19429 12795 19487 12801
rect 22002 12792 22008 12844
rect 22060 12832 22066 12844
rect 22373 12835 22431 12841
rect 22373 12832 22385 12835
rect 22060 12804 22385 12832
rect 22060 12792 22066 12804
rect 22373 12801 22385 12804
rect 22419 12801 22431 12835
rect 22373 12795 22431 12801
rect 22462 12792 22468 12844
rect 22520 12832 22526 12844
rect 23017 12835 23075 12841
rect 23017 12832 23029 12835
rect 22520 12804 23029 12832
rect 22520 12792 22526 12804
rect 23017 12801 23029 12804
rect 23063 12832 23075 12835
rect 24044 12832 24072 12940
rect 26234 12928 26240 12940
rect 26292 12928 26298 12980
rect 26329 12971 26387 12977
rect 26329 12937 26341 12971
rect 26375 12968 26387 12971
rect 26418 12968 26424 12980
rect 26375 12940 26424 12968
rect 26375 12937 26387 12940
rect 26329 12931 26387 12937
rect 26418 12928 26424 12940
rect 26476 12968 26482 12980
rect 26694 12968 26700 12980
rect 26476 12940 26700 12968
rect 26476 12928 26482 12940
rect 26694 12928 26700 12940
rect 26752 12928 26758 12980
rect 29178 12968 29184 12980
rect 29139 12940 29184 12968
rect 29178 12928 29184 12940
rect 29236 12928 29242 12980
rect 24302 12900 24308 12912
rect 24263 12872 24308 12900
rect 24302 12860 24308 12872
rect 24360 12860 24366 12912
rect 25682 12832 25688 12844
rect 23063 12804 24072 12832
rect 25643 12804 25688 12832
rect 23063 12801 23075 12804
rect 23017 12795 23075 12801
rect 25682 12792 25688 12804
rect 25740 12792 25746 12844
rect 29089 12835 29147 12841
rect 29089 12832 29101 12835
rect 27448 12804 29101 12832
rect 11698 12724 11704 12776
rect 11756 12764 11762 12776
rect 11992 12764 12020 12792
rect 11756 12736 12020 12764
rect 12345 12767 12403 12773
rect 11756 12724 11762 12736
rect 12345 12733 12357 12767
rect 12391 12764 12403 12767
rect 14090 12764 14096 12776
rect 12391 12736 14096 12764
rect 12391 12733 12403 12736
rect 12345 12727 12403 12733
rect 14090 12724 14096 12736
rect 14148 12724 14154 12776
rect 14737 12767 14795 12773
rect 14737 12733 14749 12767
rect 14783 12764 14795 12767
rect 15378 12764 15384 12776
rect 14783 12736 15384 12764
rect 14783 12733 14795 12736
rect 14737 12727 14795 12733
rect 15378 12724 15384 12736
rect 15436 12724 15442 12776
rect 15746 12724 15752 12776
rect 15804 12764 15810 12776
rect 16298 12764 16304 12776
rect 15804 12736 16304 12764
rect 15804 12724 15810 12736
rect 16298 12724 16304 12736
rect 16356 12724 16362 12776
rect 16574 12724 16580 12776
rect 16632 12764 16638 12776
rect 16853 12767 16911 12773
rect 16853 12764 16865 12767
rect 16632 12736 16865 12764
rect 16632 12724 16638 12736
rect 16853 12733 16865 12736
rect 16899 12733 16911 12767
rect 16853 12727 16911 12733
rect 18601 12767 18659 12773
rect 18601 12733 18613 12767
rect 18647 12764 18659 12767
rect 19705 12767 19763 12773
rect 19705 12764 19717 12767
rect 18647 12736 19717 12764
rect 18647 12733 18659 12736
rect 18601 12727 18659 12733
rect 19705 12733 19717 12736
rect 19751 12764 19763 12767
rect 20346 12764 20352 12776
rect 19751 12736 20352 12764
rect 19751 12733 19763 12736
rect 19705 12727 19763 12733
rect 20346 12724 20352 12736
rect 20404 12724 20410 12776
rect 20714 12724 20720 12776
rect 20772 12764 20778 12776
rect 21453 12767 21511 12773
rect 21453 12764 21465 12767
rect 20772 12736 21465 12764
rect 20772 12724 20778 12736
rect 21453 12733 21465 12736
rect 21499 12764 21511 12767
rect 23934 12764 23940 12776
rect 21499 12736 23940 12764
rect 21499 12733 21511 12736
rect 21453 12727 21511 12733
rect 22388 12708 22416 12736
rect 23934 12724 23940 12736
rect 23992 12724 23998 12776
rect 24213 12767 24271 12773
rect 24213 12733 24225 12767
rect 24259 12764 24271 12767
rect 24670 12764 24676 12776
rect 24259 12736 24676 12764
rect 24259 12733 24271 12736
rect 24213 12727 24271 12733
rect 24670 12724 24676 12736
rect 24728 12724 24734 12776
rect 25869 12767 25927 12773
rect 25869 12733 25881 12767
rect 25915 12764 25927 12767
rect 26418 12764 26424 12776
rect 25915 12736 26424 12764
rect 25915 12733 25927 12736
rect 25869 12727 25927 12733
rect 26418 12724 26424 12736
rect 26476 12724 26482 12776
rect 9416 12668 11376 12696
rect 4764 12600 7144 12628
rect 7193 12631 7251 12637
rect 4764 12588 4770 12600
rect 7193 12597 7205 12631
rect 7239 12628 7251 12631
rect 8202 12628 8208 12640
rect 7239 12600 8208 12628
rect 7239 12597 7251 12600
rect 7193 12591 7251 12597
rect 8202 12588 8208 12600
rect 8260 12588 8266 12640
rect 8570 12588 8576 12640
rect 8628 12628 8634 12640
rect 9416 12628 9444 12668
rect 11422 12656 11428 12708
rect 11480 12696 11486 12708
rect 11480 12668 11928 12696
rect 11480 12656 11486 12668
rect 8628 12600 9444 12628
rect 9493 12631 9551 12637
rect 8628 12588 8634 12600
rect 9493 12597 9505 12631
rect 9539 12628 9551 12631
rect 9674 12628 9680 12640
rect 9539 12600 9680 12628
rect 9539 12597 9551 12600
rect 9493 12591 9551 12597
rect 9674 12588 9680 12600
rect 9732 12588 9738 12640
rect 11900 12628 11928 12668
rect 18524 12668 19564 12696
rect 13817 12631 13875 12637
rect 13817 12628 13829 12631
rect 11900 12600 13829 12628
rect 13817 12597 13829 12600
rect 13863 12597 13875 12631
rect 13817 12591 13875 12597
rect 14182 12588 14188 12640
rect 14240 12628 14246 12640
rect 14458 12628 14464 12640
rect 14240 12600 14464 12628
rect 14240 12588 14246 12600
rect 14458 12588 14464 12600
rect 14516 12588 14522 12640
rect 17494 12588 17500 12640
rect 17552 12628 17558 12640
rect 18524 12628 18552 12668
rect 17552 12600 18552 12628
rect 19536 12628 19564 12668
rect 21266 12656 21272 12708
rect 21324 12696 21330 12708
rect 21726 12696 21732 12708
rect 21324 12668 21732 12696
rect 21324 12656 21330 12668
rect 21726 12656 21732 12668
rect 21784 12696 21790 12708
rect 21784 12668 22094 12696
rect 21784 12656 21790 12668
rect 21634 12628 21640 12640
rect 19536 12600 21640 12628
rect 17552 12588 17558 12600
rect 21634 12588 21640 12600
rect 21692 12588 21698 12640
rect 22066 12628 22094 12668
rect 22370 12656 22376 12708
rect 22428 12656 22434 12708
rect 22830 12656 22836 12708
rect 22888 12696 22894 12708
rect 24765 12699 24823 12705
rect 24765 12696 24777 12699
rect 22888 12668 24777 12696
rect 22888 12656 22894 12668
rect 24765 12665 24777 12668
rect 24811 12665 24823 12699
rect 24765 12659 24823 12665
rect 27448 12628 27476 12804
rect 29089 12801 29101 12804
rect 29135 12832 29147 12835
rect 30466 12832 30472 12844
rect 29135 12804 30472 12832
rect 29135 12801 29147 12804
rect 29089 12795 29147 12801
rect 30466 12792 30472 12804
rect 30524 12792 30530 12844
rect 30650 12832 30656 12844
rect 30611 12804 30656 12832
rect 30650 12792 30656 12804
rect 30708 12792 30714 12844
rect 30837 12835 30895 12841
rect 30837 12801 30849 12835
rect 30883 12832 30895 12835
rect 31294 12832 31300 12844
rect 30883 12804 31300 12832
rect 30883 12801 30895 12804
rect 30837 12795 30895 12801
rect 31294 12792 31300 12804
rect 31352 12792 31358 12844
rect 34422 12792 34428 12844
rect 34480 12832 34486 12844
rect 38013 12835 38071 12841
rect 38013 12832 38025 12835
rect 34480 12804 38025 12832
rect 34480 12792 34486 12804
rect 38013 12801 38025 12804
rect 38059 12801 38071 12835
rect 38013 12795 38071 12801
rect 27982 12764 27988 12776
rect 27943 12736 27988 12764
rect 27982 12724 27988 12736
rect 28040 12724 28046 12776
rect 28166 12764 28172 12776
rect 28127 12736 28172 12764
rect 28166 12724 28172 12736
rect 28224 12724 28230 12776
rect 29362 12656 29368 12708
rect 29420 12696 29426 12708
rect 31021 12699 31079 12705
rect 31021 12696 31033 12699
rect 29420 12668 31033 12696
rect 29420 12656 29426 12668
rect 31021 12665 31033 12668
rect 31067 12665 31079 12699
rect 31021 12659 31079 12665
rect 22066 12600 27476 12628
rect 28629 12631 28687 12637
rect 28629 12597 28641 12631
rect 28675 12628 28687 12631
rect 28994 12628 29000 12640
rect 28675 12600 29000 12628
rect 28675 12597 28687 12600
rect 28629 12591 28687 12597
rect 28994 12588 29000 12600
rect 29052 12588 29058 12640
rect 38194 12628 38200 12640
rect 38155 12600 38200 12628
rect 38194 12588 38200 12600
rect 38252 12588 38258 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 5442 12384 5448 12436
rect 5500 12424 5506 12436
rect 9214 12424 9220 12436
rect 5500 12396 9220 12424
rect 5500 12384 5506 12396
rect 9214 12384 9220 12396
rect 9272 12384 9278 12436
rect 9858 12424 9864 12436
rect 9819 12396 9864 12424
rect 9858 12384 9864 12396
rect 9916 12384 9922 12436
rect 10042 12384 10048 12436
rect 10100 12424 10106 12436
rect 10670 12427 10728 12433
rect 10670 12424 10682 12427
rect 10100 12396 10682 12424
rect 10100 12384 10106 12396
rect 10670 12393 10682 12396
rect 10716 12393 10728 12427
rect 10670 12387 10728 12393
rect 11422 12384 11428 12436
rect 11480 12424 11486 12436
rect 13262 12424 13268 12436
rect 11480 12396 13268 12424
rect 11480 12384 11486 12396
rect 13262 12384 13268 12396
rect 13320 12384 13326 12436
rect 13633 12427 13691 12433
rect 13633 12393 13645 12427
rect 13679 12424 13691 12427
rect 13814 12424 13820 12436
rect 13679 12396 13820 12424
rect 13679 12393 13691 12396
rect 13633 12387 13691 12393
rect 13814 12384 13820 12396
rect 13872 12384 13878 12436
rect 15746 12384 15752 12436
rect 15804 12424 15810 12436
rect 18506 12424 18512 12436
rect 15804 12396 17264 12424
rect 18467 12396 18512 12424
rect 15804 12384 15810 12396
rect 2958 12316 2964 12368
rect 3016 12356 3022 12368
rect 5902 12356 5908 12368
rect 3016 12328 5908 12356
rect 3016 12316 3022 12328
rect 5902 12316 5908 12328
rect 5960 12316 5966 12368
rect 10410 12356 10416 12368
rect 9784 12328 10416 12356
rect 6730 12288 6736 12300
rect 6691 12260 6736 12288
rect 6730 12248 6736 12260
rect 6788 12248 6794 12300
rect 7009 12291 7067 12297
rect 7009 12257 7021 12291
rect 7055 12288 7067 12291
rect 9674 12288 9680 12300
rect 7055 12260 9680 12288
rect 7055 12257 7067 12260
rect 7009 12251 7067 12257
rect 9674 12248 9680 12260
rect 9732 12248 9738 12300
rect 9122 12220 9128 12232
rect 9083 12192 9128 12220
rect 9122 12180 9128 12192
rect 9180 12180 9186 12232
rect 9784 12229 9812 12328
rect 10410 12316 10416 12328
rect 10468 12316 10474 12368
rect 11238 12248 11244 12300
rect 11296 12288 11302 12300
rect 11296 12260 12020 12288
rect 11296 12248 11302 12260
rect 9769 12223 9827 12229
rect 9769 12189 9781 12223
rect 9815 12189 9827 12223
rect 10410 12220 10416 12232
rect 10371 12192 10416 12220
rect 9769 12183 9827 12189
rect 10410 12180 10416 12192
rect 10468 12180 10474 12232
rect 7098 12112 7104 12164
rect 7156 12152 7162 12164
rect 7156 12124 7498 12152
rect 8312 12124 10916 12152
rect 7156 12112 7162 12124
rect 2590 12044 2596 12096
rect 2648 12084 2654 12096
rect 8312 12084 8340 12124
rect 8478 12084 8484 12096
rect 2648 12056 8340 12084
rect 8439 12056 8484 12084
rect 2648 12044 2654 12056
rect 8478 12044 8484 12056
rect 8536 12044 8542 12096
rect 9217 12087 9275 12093
rect 9217 12053 9229 12087
rect 9263 12084 9275 12087
rect 10778 12084 10784 12096
rect 9263 12056 10784 12084
rect 9263 12053 9275 12056
rect 9217 12047 9275 12053
rect 10778 12044 10784 12056
rect 10836 12044 10842 12096
rect 10888 12084 10916 12124
rect 10962 12112 10968 12164
rect 11020 12152 11026 12164
rect 11992 12152 12020 12260
rect 12250 12248 12256 12300
rect 12308 12288 12314 12300
rect 12437 12291 12495 12297
rect 12437 12288 12449 12291
rect 12308 12260 12449 12288
rect 12308 12248 12314 12260
rect 12437 12257 12449 12260
rect 12483 12257 12495 12291
rect 12437 12251 12495 12257
rect 12710 12248 12716 12300
rect 12768 12288 12774 12300
rect 14921 12291 14979 12297
rect 14921 12288 14933 12291
rect 12768 12260 14933 12288
rect 12768 12248 12774 12260
rect 14921 12257 14933 12260
rect 14967 12288 14979 12291
rect 15562 12288 15568 12300
rect 14967 12260 15568 12288
rect 14967 12257 14979 12260
rect 14921 12251 14979 12257
rect 15562 12248 15568 12260
rect 15620 12248 15626 12300
rect 15933 12291 15991 12297
rect 15933 12257 15945 12291
rect 15979 12288 15991 12291
rect 16574 12288 16580 12300
rect 15979 12260 16580 12288
rect 15979 12257 15991 12260
rect 15933 12251 15991 12257
rect 16574 12248 16580 12260
rect 16632 12248 16638 12300
rect 17236 12288 17264 12396
rect 18506 12384 18512 12396
rect 18564 12384 18570 12436
rect 20898 12424 20904 12436
rect 20088 12396 20904 12424
rect 18230 12316 18236 12368
rect 18288 12356 18294 12368
rect 20088 12356 20116 12396
rect 20898 12384 20904 12396
rect 20956 12424 20962 12436
rect 21726 12424 21732 12436
rect 20956 12396 21732 12424
rect 20956 12384 20962 12396
rect 21726 12384 21732 12396
rect 21784 12384 21790 12436
rect 22094 12384 22100 12436
rect 22152 12424 22158 12436
rect 23198 12424 23204 12436
rect 22152 12396 23204 12424
rect 22152 12384 22158 12396
rect 23198 12384 23204 12396
rect 23256 12384 23262 12436
rect 24578 12424 24584 12436
rect 23308 12396 24584 12424
rect 18288 12328 20116 12356
rect 18288 12316 18294 12328
rect 21450 12316 21456 12368
rect 21508 12356 21514 12368
rect 23308 12356 23336 12396
rect 24578 12384 24584 12396
rect 24636 12384 24642 12436
rect 26418 12424 26424 12436
rect 26379 12396 26424 12424
rect 26418 12384 26424 12396
rect 26476 12384 26482 12436
rect 28166 12384 28172 12436
rect 28224 12424 28230 12436
rect 28445 12427 28503 12433
rect 28445 12424 28457 12427
rect 28224 12396 28457 12424
rect 28224 12384 28230 12396
rect 28445 12393 28457 12396
rect 28491 12393 28503 12427
rect 28445 12387 28503 12393
rect 33778 12384 33784 12436
rect 33836 12424 33842 12436
rect 34514 12424 34520 12436
rect 33836 12396 34520 12424
rect 33836 12384 33842 12396
rect 34514 12384 34520 12396
rect 34572 12384 34578 12436
rect 24949 12359 25007 12365
rect 24949 12356 24961 12359
rect 21508 12328 23336 12356
rect 23768 12328 24961 12356
rect 21508 12316 21514 12328
rect 17957 12291 18015 12297
rect 17957 12288 17969 12291
rect 17236 12260 17969 12288
rect 17957 12257 17969 12260
rect 18003 12257 18015 12291
rect 17957 12251 18015 12257
rect 19426 12248 19432 12300
rect 19484 12288 19490 12300
rect 19981 12291 20039 12297
rect 19981 12288 19993 12291
rect 19484 12260 19993 12288
rect 19484 12248 19490 12260
rect 19981 12257 19993 12260
rect 20027 12257 20039 12291
rect 19981 12251 20039 12257
rect 20257 12291 20315 12297
rect 20257 12257 20269 12291
rect 20303 12288 20315 12291
rect 21542 12288 21548 12300
rect 20303 12260 21548 12288
rect 20303 12257 20315 12260
rect 20257 12251 20315 12257
rect 21542 12248 21548 12260
rect 21600 12248 21606 12300
rect 21910 12248 21916 12300
rect 21968 12288 21974 12300
rect 22005 12291 22063 12297
rect 22005 12288 22017 12291
rect 21968 12260 22017 12288
rect 21968 12248 21974 12260
rect 22005 12257 22017 12260
rect 22051 12257 22063 12291
rect 22005 12251 22063 12257
rect 22094 12248 22100 12300
rect 22152 12288 22158 12300
rect 22925 12291 22983 12297
rect 22925 12288 22937 12291
rect 22152 12260 22937 12288
rect 22152 12248 22158 12260
rect 22925 12257 22937 12260
rect 22971 12257 22983 12291
rect 22925 12251 22983 12257
rect 23382 12248 23388 12300
rect 23440 12288 23446 12300
rect 23477 12291 23535 12297
rect 23477 12288 23489 12291
rect 23440 12260 23489 12288
rect 23440 12248 23446 12260
rect 23477 12257 23489 12260
rect 23523 12257 23535 12291
rect 23477 12251 23535 12257
rect 12802 12180 12808 12232
rect 12860 12220 12866 12232
rect 12897 12223 12955 12229
rect 12897 12220 12909 12223
rect 12860 12192 12909 12220
rect 12860 12180 12866 12192
rect 12897 12189 12909 12192
rect 12943 12189 12955 12223
rect 12897 12183 12955 12189
rect 13541 12223 13599 12229
rect 13541 12189 13553 12223
rect 13587 12220 13599 12223
rect 13722 12220 13728 12232
rect 13587 12192 13728 12220
rect 13587 12189 13599 12192
rect 13541 12183 13599 12189
rect 13722 12180 13728 12192
rect 13780 12180 13786 12232
rect 14747 12223 14805 12229
rect 14747 12189 14759 12223
rect 14793 12220 14805 12223
rect 15470 12220 15476 12232
rect 14793 12192 15476 12220
rect 14793 12189 14805 12192
rect 14747 12183 14805 12189
rect 15470 12180 15476 12192
rect 15528 12180 15534 12232
rect 18414 12220 18420 12232
rect 18375 12192 18420 12220
rect 18414 12180 18420 12192
rect 18472 12180 18478 12232
rect 21634 12180 21640 12232
rect 21692 12220 21698 12232
rect 21692 12192 22324 12220
rect 21692 12180 21698 12192
rect 14826 12152 14832 12164
rect 11020 12124 11178 12152
rect 11992 12124 14832 12152
rect 11020 12112 11026 12124
rect 14826 12112 14832 12124
rect 14884 12112 14890 12164
rect 16209 12155 16267 12161
rect 16209 12121 16221 12155
rect 16255 12152 16267 12155
rect 16482 12152 16488 12164
rect 16255 12124 16488 12152
rect 16255 12121 16267 12124
rect 16209 12115 16267 12121
rect 16482 12112 16488 12124
rect 16540 12112 16546 12164
rect 16666 12112 16672 12164
rect 16724 12112 16730 12164
rect 19978 12152 19984 12164
rect 19260 12124 19984 12152
rect 12710 12084 12716 12096
rect 10888 12056 12716 12084
rect 12710 12044 12716 12056
rect 12768 12044 12774 12096
rect 12989 12087 13047 12093
rect 12989 12053 13001 12087
rect 13035 12084 13047 12087
rect 19260 12084 19288 12124
rect 19978 12112 19984 12124
rect 20036 12112 20042 12164
rect 21482 12124 22094 12152
rect 22066 12096 22094 12124
rect 13035 12056 19288 12084
rect 13035 12053 13047 12056
rect 12989 12047 13047 12053
rect 19334 12044 19340 12096
rect 19392 12084 19398 12096
rect 19518 12084 19524 12096
rect 19392 12056 19524 12084
rect 19392 12044 19398 12056
rect 19518 12044 19524 12056
rect 19576 12044 19582 12096
rect 22066 12056 22100 12096
rect 22094 12044 22100 12056
rect 22152 12044 22158 12096
rect 22296 12084 22324 12192
rect 22370 12112 22376 12164
rect 22428 12152 22434 12164
rect 23017 12155 23075 12161
rect 23017 12152 23029 12155
rect 22428 12124 23029 12152
rect 22428 12112 22434 12124
rect 23017 12121 23029 12124
rect 23063 12121 23075 12155
rect 23017 12115 23075 12121
rect 23290 12112 23296 12164
rect 23348 12152 23354 12164
rect 23768 12152 23796 12328
rect 24949 12325 24961 12328
rect 24995 12325 25007 12359
rect 24949 12319 25007 12325
rect 23348 12124 23796 12152
rect 23860 12260 25728 12288
rect 23348 12112 23354 12124
rect 23566 12084 23572 12096
rect 22296 12056 23572 12084
rect 23566 12044 23572 12056
rect 23624 12084 23630 12096
rect 23860 12084 23888 12260
rect 24581 12223 24639 12229
rect 24581 12189 24593 12223
rect 24627 12189 24639 12223
rect 24762 12220 24768 12232
rect 24723 12192 24768 12220
rect 24581 12183 24639 12189
rect 24596 12152 24624 12183
rect 24762 12180 24768 12192
rect 24820 12180 24826 12232
rect 25700 12229 25728 12260
rect 25685 12223 25743 12229
rect 25685 12189 25697 12223
rect 25731 12189 25743 12223
rect 26326 12220 26332 12232
rect 26287 12192 26332 12220
rect 25685 12183 25743 12189
rect 26326 12180 26332 12192
rect 26384 12180 26390 12232
rect 28350 12220 28356 12232
rect 28311 12192 28356 12220
rect 28350 12180 28356 12192
rect 28408 12180 28414 12232
rect 30101 12223 30159 12229
rect 30101 12189 30113 12223
rect 30147 12220 30159 12223
rect 30466 12220 30472 12232
rect 30147 12192 30472 12220
rect 30147 12189 30159 12192
rect 30101 12183 30159 12189
rect 30466 12180 30472 12192
rect 30524 12180 30530 12232
rect 25130 12152 25136 12164
rect 24596 12124 25136 12152
rect 25130 12112 25136 12124
rect 25188 12112 25194 12164
rect 28258 12152 28264 12164
rect 25240 12124 28264 12152
rect 23624 12056 23888 12084
rect 23624 12044 23630 12056
rect 24486 12044 24492 12096
rect 24544 12084 24550 12096
rect 25240 12084 25268 12124
rect 28258 12112 28264 12124
rect 28316 12112 28322 12164
rect 24544 12056 25268 12084
rect 24544 12044 24550 12056
rect 25314 12044 25320 12096
rect 25372 12084 25378 12096
rect 25777 12087 25835 12093
rect 25777 12084 25789 12087
rect 25372 12056 25789 12084
rect 25372 12044 25378 12056
rect 25777 12053 25789 12056
rect 25823 12053 25835 12087
rect 25777 12047 25835 12053
rect 29454 12044 29460 12096
rect 29512 12084 29518 12096
rect 29917 12087 29975 12093
rect 29917 12084 29929 12087
rect 29512 12056 29929 12084
rect 29512 12044 29518 12056
rect 29917 12053 29929 12056
rect 29963 12053 29975 12087
rect 29917 12047 29975 12053
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 10410 11880 10416 11892
rect 7944 11852 10416 11880
rect 7944 11753 7972 11852
rect 10410 11840 10416 11852
rect 10468 11840 10474 11892
rect 10778 11840 10784 11892
rect 10836 11880 10842 11892
rect 10836 11852 14412 11880
rect 10836 11840 10842 11852
rect 8202 11772 8208 11824
rect 8260 11812 8266 11824
rect 11514 11812 11520 11824
rect 8260 11784 8694 11812
rect 9876 11784 11520 11812
rect 8260 11772 8266 11784
rect 7929 11747 7987 11753
rect 7929 11713 7941 11747
rect 7975 11713 7987 11747
rect 7929 11707 7987 11713
rect 8205 11679 8263 11685
rect 8205 11645 8217 11679
rect 8251 11676 8263 11679
rect 9876 11676 9904 11784
rect 11514 11772 11520 11784
rect 11572 11772 11578 11824
rect 11882 11772 11888 11824
rect 11940 11812 11946 11824
rect 11977 11815 12035 11821
rect 11977 11812 11989 11815
rect 11940 11784 11989 11812
rect 11940 11772 11946 11784
rect 11977 11781 11989 11784
rect 12023 11781 12035 11815
rect 11977 11775 12035 11781
rect 12434 11772 12440 11824
rect 12492 11772 12498 11824
rect 14277 11815 14335 11821
rect 14277 11812 14289 11815
rect 13372 11784 14289 11812
rect 9953 11747 10011 11753
rect 9953 11713 9965 11747
rect 9999 11744 10011 11747
rect 10318 11744 10324 11756
rect 9999 11716 10324 11744
rect 9999 11713 10011 11716
rect 9953 11707 10011 11713
rect 10318 11704 10324 11716
rect 10376 11704 10382 11756
rect 10686 11704 10692 11756
rect 10744 11744 10750 11756
rect 10965 11747 11023 11753
rect 10965 11744 10977 11747
rect 10744 11716 10977 11744
rect 10744 11704 10750 11716
rect 10965 11713 10977 11716
rect 11011 11713 11023 11747
rect 10965 11707 11023 11713
rect 11054 11704 11060 11756
rect 11112 11744 11118 11756
rect 11701 11747 11759 11753
rect 11701 11744 11713 11747
rect 11112 11716 11713 11744
rect 11112 11704 11118 11716
rect 11701 11713 11713 11716
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 8251 11648 9904 11676
rect 8251 11645 8263 11648
rect 8205 11639 8263 11645
rect 10410 11636 10416 11688
rect 10468 11676 10474 11688
rect 11072 11676 11100 11704
rect 10468 11648 11100 11676
rect 10468 11636 10474 11648
rect 11146 11636 11152 11688
rect 11204 11676 11210 11688
rect 13372 11676 13400 11784
rect 14277 11781 14289 11784
rect 14323 11781 14335 11815
rect 14384 11812 14412 11852
rect 14550 11840 14556 11892
rect 14608 11880 14614 11892
rect 15746 11880 15752 11892
rect 14608 11852 15752 11880
rect 14608 11840 14614 11852
rect 15746 11840 15752 11852
rect 15804 11840 15810 11892
rect 16482 11840 16488 11892
rect 16540 11880 16546 11892
rect 18230 11880 18236 11892
rect 16540 11852 18236 11880
rect 16540 11840 16546 11852
rect 18230 11840 18236 11852
rect 18288 11840 18294 11892
rect 18877 11883 18935 11889
rect 18877 11849 18889 11883
rect 18923 11880 18935 11883
rect 19334 11880 19340 11892
rect 18923 11852 19340 11880
rect 18923 11849 18935 11852
rect 18877 11843 18935 11849
rect 19334 11840 19340 11852
rect 19392 11840 19398 11892
rect 22370 11880 22376 11892
rect 19444 11852 22094 11880
rect 22331 11852 22376 11880
rect 14384 11784 14766 11812
rect 14277 11775 14335 11781
rect 17402 11772 17408 11824
rect 17460 11812 17466 11824
rect 17460 11784 17505 11812
rect 17460 11772 17466 11784
rect 17862 11772 17868 11824
rect 17920 11772 17926 11824
rect 18966 11772 18972 11824
rect 19024 11812 19030 11824
rect 19444 11812 19472 11852
rect 21174 11812 21180 11824
rect 19024 11784 19472 11812
rect 20930 11784 21180 11812
rect 19024 11772 19030 11784
rect 21174 11772 21180 11784
rect 21232 11772 21238 11824
rect 22066 11812 22094 11852
rect 22370 11840 22376 11852
rect 22428 11840 22434 11892
rect 24762 11880 24768 11892
rect 23124 11852 24624 11880
rect 24723 11852 24768 11880
rect 23124 11812 23152 11852
rect 23290 11812 23296 11824
rect 22066 11784 23152 11812
rect 23251 11784 23296 11812
rect 23290 11772 23296 11784
rect 23348 11772 23354 11824
rect 23382 11772 23388 11824
rect 23440 11812 23446 11824
rect 24596 11812 24624 11852
rect 24762 11840 24768 11852
rect 24820 11840 24826 11892
rect 26326 11880 26332 11892
rect 25332 11852 26332 11880
rect 25332 11812 25360 11852
rect 26326 11840 26332 11852
rect 26384 11840 26390 11892
rect 30466 11880 30472 11892
rect 30427 11852 30472 11880
rect 30466 11840 30472 11852
rect 30524 11840 30530 11892
rect 30834 11840 30840 11892
rect 30892 11880 30898 11892
rect 32401 11883 32459 11889
rect 32401 11880 32413 11883
rect 30892 11852 32413 11880
rect 30892 11840 30898 11852
rect 32401 11849 32413 11852
rect 32447 11849 32459 11883
rect 32401 11843 32459 11849
rect 25498 11812 25504 11824
rect 23440 11784 24532 11812
rect 24596 11784 25360 11812
rect 25459 11784 25504 11812
rect 23440 11772 23446 11784
rect 16574 11704 16580 11756
rect 16632 11744 16638 11756
rect 17129 11747 17187 11753
rect 17129 11744 17141 11747
rect 16632 11716 17141 11744
rect 16632 11704 16638 11716
rect 17129 11713 17141 11716
rect 17175 11713 17187 11747
rect 19426 11744 19432 11756
rect 19387 11716 19432 11744
rect 17129 11707 17187 11713
rect 19426 11704 19432 11716
rect 19484 11704 19490 11756
rect 21082 11744 21088 11756
rect 20995 11716 21088 11744
rect 13998 11676 14004 11688
rect 11204 11648 13400 11676
rect 13911 11648 14004 11676
rect 11204 11636 11210 11648
rect 13998 11636 14004 11648
rect 14056 11676 14062 11688
rect 16666 11676 16672 11688
rect 14056 11648 16672 11676
rect 14056 11636 14062 11648
rect 16666 11636 16672 11648
rect 16724 11636 16730 11688
rect 19705 11679 19763 11685
rect 19705 11645 19717 11679
rect 19751 11676 19763 11679
rect 21008 11676 21036 11716
rect 21082 11704 21088 11716
rect 21140 11744 21146 11756
rect 22281 11747 22339 11753
rect 21140 11716 22094 11744
rect 21140 11704 21146 11716
rect 19751 11648 21036 11676
rect 21453 11679 21511 11685
rect 19751 11645 19763 11648
rect 19705 11639 19763 11645
rect 21453 11645 21465 11679
rect 21499 11645 21511 11679
rect 21453 11639 21511 11645
rect 9214 11568 9220 11620
rect 9272 11608 9278 11620
rect 9858 11608 9864 11620
rect 9272 11580 9864 11608
rect 9272 11568 9278 11580
rect 9858 11568 9864 11580
rect 9916 11568 9922 11620
rect 18874 11568 18880 11620
rect 18932 11608 18938 11620
rect 18932 11580 19564 11608
rect 18932 11568 18938 11580
rect 5626 11500 5632 11552
rect 5684 11540 5690 11552
rect 10962 11540 10968 11552
rect 5684 11512 10968 11540
rect 5684 11500 5690 11512
rect 10962 11500 10968 11512
rect 11020 11500 11026 11552
rect 11057 11543 11115 11549
rect 11057 11509 11069 11543
rect 11103 11540 11115 11543
rect 11238 11540 11244 11552
rect 11103 11512 11244 11540
rect 11103 11509 11115 11512
rect 11057 11503 11115 11509
rect 11238 11500 11244 11512
rect 11296 11500 11302 11552
rect 13354 11500 13360 11552
rect 13412 11540 13418 11552
rect 13449 11543 13507 11549
rect 13449 11540 13461 11543
rect 13412 11512 13461 11540
rect 13412 11500 13418 11512
rect 13449 11509 13461 11512
rect 13495 11509 13507 11543
rect 13449 11503 13507 11509
rect 15749 11543 15807 11549
rect 15749 11509 15761 11543
rect 15795 11540 15807 11543
rect 17126 11540 17132 11552
rect 15795 11512 17132 11540
rect 15795 11509 15807 11512
rect 15749 11503 15807 11509
rect 17126 11500 17132 11512
rect 17184 11540 17190 11552
rect 18966 11540 18972 11552
rect 17184 11512 18972 11540
rect 17184 11500 17190 11512
rect 18966 11500 18972 11512
rect 19024 11500 19030 11552
rect 19536 11540 19564 11580
rect 21468 11540 21496 11639
rect 19536 11512 21496 11540
rect 22066 11540 22094 11716
rect 22281 11713 22293 11747
rect 22327 11713 22339 11747
rect 24504 11744 24532 11784
rect 25498 11772 25504 11784
rect 25556 11772 25562 11824
rect 26786 11772 26792 11824
rect 26844 11812 26850 11824
rect 27249 11815 27307 11821
rect 27249 11812 27261 11815
rect 26844 11784 27261 11812
rect 26844 11772 26850 11784
rect 27249 11781 27261 11784
rect 27295 11781 27307 11815
rect 27249 11775 27307 11781
rect 27341 11815 27399 11821
rect 27341 11781 27353 11815
rect 27387 11812 27399 11815
rect 27890 11812 27896 11824
rect 27387 11784 27896 11812
rect 27387 11781 27399 11784
rect 27341 11775 27399 11781
rect 27890 11772 27896 11784
rect 27948 11772 27954 11824
rect 29362 11812 29368 11824
rect 29323 11784 29368 11812
rect 29362 11772 29368 11784
rect 29420 11772 29426 11824
rect 29454 11772 29460 11824
rect 29512 11812 29518 11824
rect 29512 11784 29557 11812
rect 29512 11772 29518 11784
rect 24673 11747 24731 11753
rect 24673 11744 24685 11747
rect 24504 11716 24685 11744
rect 22281 11707 22339 11713
rect 24673 11713 24685 11716
rect 24719 11713 24731 11747
rect 30650 11744 30656 11756
rect 30611 11716 30656 11744
rect 24673 11707 24731 11713
rect 22296 11620 22324 11707
rect 30650 11704 30656 11716
rect 30708 11704 30714 11756
rect 32309 11747 32367 11753
rect 32309 11713 32321 11747
rect 32355 11744 32367 11747
rect 34054 11744 34060 11756
rect 32355 11716 34060 11744
rect 32355 11713 32367 11716
rect 32309 11707 32367 11713
rect 34054 11704 34060 11716
rect 34112 11704 34118 11756
rect 23201 11679 23259 11685
rect 23201 11645 23213 11679
rect 23247 11645 23259 11679
rect 23201 11639 23259 11645
rect 22278 11568 22284 11620
rect 22336 11568 22342 11620
rect 23216 11608 23244 11639
rect 23658 11636 23664 11688
rect 23716 11676 23722 11688
rect 24210 11676 24216 11688
rect 23716 11648 24216 11676
rect 23716 11636 23722 11648
rect 24210 11636 24216 11648
rect 24268 11676 24274 11688
rect 25409 11679 25467 11685
rect 24268 11648 25360 11676
rect 24268 11636 24274 11648
rect 24670 11608 24676 11620
rect 23216 11580 24676 11608
rect 24670 11568 24676 11580
rect 24728 11568 24734 11620
rect 25332 11608 25360 11648
rect 25409 11645 25421 11679
rect 25455 11676 25467 11679
rect 26234 11676 26240 11688
rect 25455 11648 26240 11676
rect 25455 11645 25467 11648
rect 25409 11639 25467 11645
rect 26234 11636 26240 11648
rect 26292 11636 26298 11688
rect 26329 11679 26387 11685
rect 26329 11645 26341 11679
rect 26375 11645 26387 11679
rect 27614 11676 27620 11688
rect 27575 11648 27620 11676
rect 26329 11639 26387 11645
rect 26344 11608 26372 11639
rect 27614 11636 27620 11648
rect 27672 11676 27678 11688
rect 29641 11679 29699 11685
rect 29641 11676 29653 11679
rect 27672 11648 29653 11676
rect 27672 11636 27678 11648
rect 29641 11645 29653 11648
rect 29687 11645 29699 11679
rect 29641 11639 29699 11645
rect 25332 11580 26372 11608
rect 28350 11540 28356 11552
rect 22066 11512 28356 11540
rect 28350 11500 28356 11512
rect 28408 11540 28414 11552
rect 29914 11540 29920 11552
rect 28408 11512 29920 11540
rect 28408 11500 28414 11512
rect 29914 11500 29920 11512
rect 29972 11500 29978 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 2516 11308 2774 11336
rect 1762 11132 1768 11144
rect 1723 11104 1768 11132
rect 1762 11092 1768 11104
rect 1820 11092 1826 11144
rect 2516 11141 2544 11308
rect 2746 11268 2774 11308
rect 5718 11296 5724 11348
rect 5776 11336 5782 11348
rect 5776 11308 8432 11336
rect 5776 11296 5782 11308
rect 6454 11268 6460 11280
rect 2746 11240 6460 11268
rect 6454 11228 6460 11240
rect 6512 11228 6518 11280
rect 8404 11268 8432 11308
rect 8478 11296 8484 11348
rect 8536 11336 8542 11348
rect 11146 11336 11152 11348
rect 8536 11308 11152 11336
rect 8536 11296 8542 11308
rect 11146 11296 11152 11308
rect 11204 11296 11210 11348
rect 11964 11339 12022 11345
rect 11964 11305 11976 11339
rect 12010 11336 12022 11339
rect 12010 11308 13952 11336
rect 12010 11305 12022 11308
rect 11964 11299 12022 11305
rect 8662 11268 8668 11280
rect 8404 11240 8668 11268
rect 8662 11228 8668 11240
rect 8720 11268 8726 11280
rect 9490 11268 9496 11280
rect 8720 11240 9496 11268
rect 8720 11228 8726 11240
rect 9490 11228 9496 11240
rect 9548 11228 9554 11280
rect 12986 11228 12992 11280
rect 13044 11268 13050 11280
rect 13354 11268 13360 11280
rect 13044 11240 13360 11268
rect 13044 11228 13050 11240
rect 13354 11228 13360 11240
rect 13412 11228 13418 11280
rect 13924 11268 13952 11308
rect 22094 11296 22100 11348
rect 22152 11336 22158 11348
rect 23198 11336 23204 11348
rect 22152 11308 23060 11336
rect 23159 11308 23204 11336
rect 22152 11296 22158 11308
rect 14090 11268 14096 11280
rect 13924 11240 14096 11268
rect 14090 11228 14096 11240
rect 14148 11228 14154 11280
rect 18874 11228 18880 11280
rect 18932 11268 18938 11280
rect 22278 11268 22284 11280
rect 18932 11240 22284 11268
rect 18932 11228 18938 11240
rect 22278 11228 22284 11240
rect 22336 11228 22342 11280
rect 23032 11268 23060 11308
rect 23198 11296 23204 11308
rect 23256 11296 23262 11348
rect 23842 11336 23848 11348
rect 23803 11308 23848 11336
rect 23842 11296 23848 11308
rect 23900 11296 23906 11348
rect 27890 11336 27896 11348
rect 27851 11308 27896 11336
rect 27890 11296 27896 11308
rect 27948 11296 27954 11348
rect 23566 11268 23572 11280
rect 23032 11240 23572 11268
rect 23566 11228 23572 11240
rect 23624 11228 23630 11280
rect 25130 11228 25136 11280
rect 25188 11268 25194 11280
rect 27798 11268 27804 11280
rect 25188 11240 27804 11268
rect 25188 11228 25194 11240
rect 27798 11228 27804 11240
rect 27856 11228 27862 11280
rect 38194 11268 38200 11280
rect 38155 11240 38200 11268
rect 38194 11228 38200 11240
rect 38252 11228 38258 11280
rect 6730 11160 6736 11212
rect 6788 11200 6794 11212
rect 6825 11203 6883 11209
rect 6825 11200 6837 11203
rect 6788 11172 6837 11200
rect 6788 11160 6794 11172
rect 6825 11169 6837 11172
rect 6871 11169 6883 11203
rect 6825 11163 6883 11169
rect 7101 11203 7159 11209
rect 7101 11169 7113 11203
rect 7147 11200 7159 11203
rect 8573 11203 8631 11209
rect 7147 11172 8524 11200
rect 7147 11169 7159 11172
rect 7101 11163 7159 11169
rect 2501 11135 2559 11141
rect 2501 11101 2513 11135
rect 2547 11101 2559 11135
rect 8496 11132 8524 11172
rect 8573 11169 8585 11203
rect 8619 11200 8631 11203
rect 9769 11203 9827 11209
rect 8619 11172 9352 11200
rect 8619 11169 8631 11172
rect 8573 11163 8631 11169
rect 8496 11104 8984 11132
rect 2501 11095 2559 11101
rect 8956 11076 8984 11104
rect 5994 11064 6000 11076
rect 1596 11036 6000 11064
rect 1596 11005 1624 11036
rect 5994 11024 6000 11036
rect 6052 11024 6058 11076
rect 6546 11024 6552 11076
rect 6604 11064 6610 11076
rect 6604 11036 7052 11064
rect 6604 11024 6610 11036
rect 1581 10999 1639 11005
rect 1581 10965 1593 10999
rect 1627 10965 1639 10999
rect 2314 10996 2320 11008
rect 2275 10968 2320 10996
rect 1581 10959 1639 10965
rect 2314 10956 2320 10968
rect 2372 10956 2378 11008
rect 7024 10996 7052 11036
rect 7208 11036 7590 11064
rect 7208 10996 7236 11036
rect 8938 11024 8944 11076
rect 8996 11064 9002 11076
rect 9324 11064 9352 11172
rect 9769 11169 9781 11203
rect 9815 11200 9827 11203
rect 10778 11200 10784 11212
rect 9815 11172 10784 11200
rect 9815 11169 9827 11172
rect 9769 11163 9827 11169
rect 10778 11160 10784 11172
rect 10836 11160 10842 11212
rect 11698 11200 11704 11212
rect 11659 11172 11704 11200
rect 11698 11160 11704 11172
rect 11756 11160 11762 11212
rect 12526 11160 12532 11212
rect 12584 11200 12590 11212
rect 13725 11203 13783 11209
rect 13725 11200 13737 11203
rect 12584 11172 13737 11200
rect 12584 11160 12590 11172
rect 13725 11169 13737 11172
rect 13771 11169 13783 11203
rect 13725 11163 13783 11169
rect 14277 11203 14335 11209
rect 14277 11169 14289 11203
rect 14323 11200 14335 11203
rect 16574 11200 16580 11212
rect 14323 11172 16580 11200
rect 14323 11169 14335 11172
rect 14277 11163 14335 11169
rect 16574 11160 16580 11172
rect 16632 11160 16638 11212
rect 16666 11160 16672 11212
rect 16724 11200 16730 11212
rect 16761 11203 16819 11209
rect 16761 11200 16773 11203
rect 16724 11172 16773 11200
rect 16724 11160 16730 11172
rect 16761 11169 16773 11172
rect 16807 11169 16819 11203
rect 16761 11163 16819 11169
rect 17037 11203 17095 11209
rect 17037 11169 17049 11203
rect 17083 11200 17095 11203
rect 18046 11200 18052 11212
rect 17083 11172 18052 11200
rect 17083 11169 17095 11172
rect 17037 11163 17095 11169
rect 18046 11160 18052 11172
rect 18104 11200 18110 11212
rect 18230 11200 18236 11212
rect 18104 11172 18236 11200
rect 18104 11160 18110 11172
rect 18230 11160 18236 11172
rect 18288 11160 18294 11212
rect 18506 11200 18512 11212
rect 18467 11172 18512 11200
rect 18506 11160 18512 11172
rect 18564 11200 18570 11212
rect 18782 11200 18788 11212
rect 18564 11172 18788 11200
rect 18564 11160 18570 11172
rect 18782 11160 18788 11172
rect 18840 11160 18846 11212
rect 19242 11160 19248 11212
rect 19300 11200 19306 11212
rect 19426 11200 19432 11212
rect 19300 11172 19432 11200
rect 19300 11160 19306 11172
rect 19426 11160 19432 11172
rect 19484 11200 19490 11212
rect 20165 11203 20223 11209
rect 20165 11200 20177 11203
rect 19484 11172 20177 11200
rect 19484 11160 19490 11172
rect 20165 11169 20177 11172
rect 20211 11169 20223 11203
rect 20165 11163 20223 11169
rect 21542 11160 21548 11212
rect 21600 11200 21606 11212
rect 26234 11200 26240 11212
rect 21600 11172 26096 11200
rect 26195 11172 26240 11200
rect 21600 11160 21606 11172
rect 9490 11132 9496 11144
rect 9451 11104 9496 11132
rect 9490 11092 9496 11104
rect 9548 11092 9554 11144
rect 10870 11092 10876 11144
rect 10928 11092 10934 11144
rect 18598 11092 18604 11144
rect 18656 11132 18662 11144
rect 23014 11132 23020 11144
rect 18656 11104 23020 11132
rect 18656 11092 18662 11104
rect 23014 11092 23020 11104
rect 23072 11132 23078 11144
rect 23109 11135 23167 11141
rect 23109 11132 23121 11135
rect 23072 11104 23121 11132
rect 23072 11092 23078 11104
rect 23109 11101 23121 11104
rect 23155 11101 23167 11135
rect 23109 11095 23167 11101
rect 23753 11135 23811 11141
rect 23753 11101 23765 11135
rect 23799 11132 23811 11135
rect 24210 11132 24216 11144
rect 23799 11104 24216 11132
rect 23799 11101 23811 11104
rect 23753 11095 23811 11101
rect 9674 11064 9680 11076
rect 8996 11036 9260 11064
rect 9324 11036 9680 11064
rect 8996 11024 9002 11036
rect 7024 10968 7236 10996
rect 7374 10956 7380 11008
rect 7432 10996 7438 11008
rect 8110 10996 8116 11008
rect 7432 10968 8116 10996
rect 7432 10956 7438 10968
rect 8110 10956 8116 10968
rect 8168 10956 8174 11008
rect 9232 10996 9260 11036
rect 9674 11024 9680 11036
rect 9732 11024 9738 11076
rect 11974 11024 11980 11076
rect 12032 11064 12038 11076
rect 12032 11036 12466 11064
rect 12032 11024 12038 11036
rect 13354 11024 13360 11076
rect 13412 11064 13418 11076
rect 13998 11064 14004 11076
rect 13412 11036 14004 11064
rect 13412 11024 13418 11036
rect 13998 11024 14004 11036
rect 14056 11024 14062 11076
rect 14550 11064 14556 11076
rect 14511 11036 14556 11064
rect 14550 11024 14556 11036
rect 14608 11024 14614 11076
rect 14826 11024 14832 11076
rect 14884 11064 14890 11076
rect 16298 11064 16304 11076
rect 14884 11036 15042 11064
rect 16211 11036 16304 11064
rect 14884 11024 14890 11036
rect 16298 11024 16304 11036
rect 16356 11064 16362 11076
rect 17034 11064 17040 11076
rect 16356 11036 17040 11064
rect 16356 11024 16362 11036
rect 17034 11024 17040 11036
rect 17092 11024 17098 11076
rect 18322 11064 18328 11076
rect 18262 11036 18328 11064
rect 18322 11024 18328 11036
rect 18380 11024 18386 11076
rect 19426 11064 19432 11076
rect 18432 11036 18644 11064
rect 19387 11036 19432 11064
rect 11241 10999 11299 11005
rect 11241 10996 11253 10999
rect 9232 10968 11253 10996
rect 11241 10965 11253 10968
rect 11287 10965 11299 10999
rect 11241 10959 11299 10965
rect 11514 10956 11520 11008
rect 11572 10996 11578 11008
rect 18432 10996 18460 11036
rect 11572 10968 18460 10996
rect 18616 10996 18644 11036
rect 19426 11024 19432 11036
rect 19484 11024 19490 11076
rect 22002 11024 22008 11076
rect 22060 11064 22066 11076
rect 23768 11064 23796 11095
rect 24210 11092 24216 11104
rect 24268 11092 24274 11144
rect 26068 11132 26096 11172
rect 26234 11160 26240 11172
rect 26292 11160 26298 11212
rect 28442 11200 28448 11212
rect 28403 11172 28448 11200
rect 28442 11160 28448 11172
rect 28500 11160 28506 11212
rect 30650 11200 30656 11212
rect 28552 11172 30656 11200
rect 27801 11135 27859 11141
rect 27801 11132 27813 11135
rect 26068 11104 27813 11132
rect 27801 11101 27813 11104
rect 27847 11132 27859 11135
rect 28552 11132 28580 11172
rect 30650 11160 30656 11172
rect 30708 11160 30714 11212
rect 27847 11104 28580 11132
rect 28629 11135 28687 11141
rect 27847 11101 27859 11104
rect 27801 11095 27859 11101
rect 28629 11101 28641 11135
rect 28675 11132 28687 11135
rect 29270 11132 29276 11144
rect 28675 11104 29276 11132
rect 28675 11101 28687 11104
rect 28629 11095 28687 11101
rect 29270 11092 29276 11104
rect 29328 11092 29334 11144
rect 29914 11132 29920 11144
rect 29875 11104 29920 11132
rect 29914 11092 29920 11104
rect 29972 11092 29978 11144
rect 37366 11132 37372 11144
rect 37327 11104 37372 11132
rect 37366 11092 37372 11104
rect 37424 11092 37430 11144
rect 38013 11135 38071 11141
rect 38013 11101 38025 11135
rect 38059 11101 38071 11135
rect 38013 11095 38071 11101
rect 25130 11064 25136 11076
rect 22060 11036 23796 11064
rect 25091 11036 25136 11064
rect 22060 11024 22066 11036
rect 25130 11024 25136 11036
rect 25188 11024 25194 11076
rect 25225 11067 25283 11073
rect 25225 11033 25237 11067
rect 25271 11064 25283 11067
rect 25314 11064 25320 11076
rect 25271 11036 25320 11064
rect 25271 11033 25283 11036
rect 25225 11027 25283 11033
rect 25314 11024 25320 11036
rect 25372 11024 25378 11076
rect 25406 11024 25412 11076
rect 25464 11064 25470 11076
rect 25777 11067 25835 11073
rect 25777 11064 25789 11067
rect 25464 11036 25789 11064
rect 25464 11024 25470 11036
rect 25777 11033 25789 11036
rect 25823 11064 25835 11067
rect 25866 11064 25872 11076
rect 25823 11036 25872 11064
rect 25823 11033 25835 11036
rect 25777 11027 25835 11033
rect 25866 11024 25872 11036
rect 25924 11024 25930 11076
rect 29086 11064 29092 11076
rect 29047 11036 29092 11064
rect 29086 11024 29092 11036
rect 29144 11024 29150 11076
rect 36906 11024 36912 11076
rect 36964 11064 36970 11076
rect 38028 11064 38056 11095
rect 36964 11036 38056 11064
rect 36964 11024 36970 11036
rect 28994 10996 29000 11008
rect 18616 10968 29000 10996
rect 11572 10956 11578 10968
rect 28994 10956 29000 10968
rect 29052 10956 29058 11008
rect 29454 10956 29460 11008
rect 29512 10996 29518 11008
rect 29733 10999 29791 11005
rect 29733 10996 29745 10999
rect 29512 10968 29745 10996
rect 29512 10956 29518 10968
rect 29733 10965 29745 10968
rect 29779 10965 29791 10999
rect 37458 10996 37464 11008
rect 37419 10968 37464 10996
rect 29733 10959 29791 10965
rect 37458 10956 37464 10968
rect 37516 10956 37522 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 1581 10795 1639 10801
rect 1581 10761 1593 10795
rect 1627 10792 1639 10795
rect 1946 10792 1952 10804
rect 1627 10764 1952 10792
rect 1627 10761 1639 10764
rect 1581 10755 1639 10761
rect 1946 10752 1952 10764
rect 2004 10752 2010 10804
rect 3789 10795 3847 10801
rect 3789 10761 3801 10795
rect 3835 10792 3847 10795
rect 4798 10792 4804 10804
rect 3835 10764 4804 10792
rect 3835 10761 3847 10764
rect 3789 10755 3847 10761
rect 4798 10752 4804 10764
rect 4856 10752 4862 10804
rect 7374 10752 7380 10804
rect 7432 10752 7438 10804
rect 7926 10752 7932 10804
rect 7984 10792 7990 10804
rect 9033 10795 9091 10801
rect 9033 10792 9045 10795
rect 7984 10764 9045 10792
rect 7984 10752 7990 10764
rect 9033 10761 9045 10764
rect 9079 10761 9091 10795
rect 9033 10755 9091 10761
rect 10870 10752 10876 10804
rect 10928 10792 10934 10804
rect 12161 10795 12219 10801
rect 12161 10792 12173 10795
rect 10928 10764 12173 10792
rect 10928 10752 10934 10764
rect 12161 10761 12173 10764
rect 12207 10761 12219 10795
rect 12161 10755 12219 10761
rect 12342 10752 12348 10804
rect 12400 10792 12406 10804
rect 12618 10792 12624 10804
rect 12400 10764 12624 10792
rect 12400 10752 12406 10764
rect 12618 10752 12624 10764
rect 12676 10752 12682 10804
rect 12805 10795 12863 10801
rect 12805 10761 12817 10795
rect 12851 10792 12863 10795
rect 15105 10795 15163 10801
rect 12851 10764 13492 10792
rect 12851 10761 12863 10764
rect 12805 10755 12863 10761
rect 7392 10724 7420 10752
rect 4816 10696 7420 10724
rect 4816 10668 4844 10696
rect 7466 10684 7472 10736
rect 7524 10724 7530 10736
rect 10318 10724 10324 10736
rect 7524 10696 8050 10724
rect 9646 10696 10324 10724
rect 7524 10684 7530 10696
rect 1762 10656 1768 10668
rect 1723 10628 1768 10656
rect 1762 10616 1768 10628
rect 1820 10616 1826 10668
rect 2593 10659 2651 10665
rect 2593 10625 2605 10659
rect 2639 10656 2651 10659
rect 2774 10656 2780 10668
rect 2639 10628 2780 10656
rect 2639 10625 2651 10628
rect 2593 10619 2651 10625
rect 2774 10616 2780 10628
rect 2832 10616 2838 10668
rect 3697 10659 3755 10665
rect 3697 10625 3709 10659
rect 3743 10625 3755 10659
rect 3697 10619 3755 10625
rect 1946 10548 1952 10600
rect 2004 10588 2010 10600
rect 3712 10588 3740 10619
rect 4798 10616 4804 10668
rect 4856 10616 4862 10668
rect 2004 10560 3740 10588
rect 2004 10548 2010 10560
rect 6822 10548 6828 10600
rect 6880 10588 6886 10600
rect 7285 10591 7343 10597
rect 7285 10588 7297 10591
rect 6880 10560 7297 10588
rect 6880 10548 6886 10560
rect 7285 10557 7297 10560
rect 7331 10557 7343 10591
rect 7285 10551 7343 10557
rect 7561 10591 7619 10597
rect 7561 10557 7573 10591
rect 7607 10588 7619 10591
rect 9646 10588 9674 10696
rect 10318 10684 10324 10696
rect 10376 10684 10382 10736
rect 10502 10684 10508 10736
rect 10560 10724 10566 10736
rect 10686 10724 10692 10736
rect 10560 10696 10692 10724
rect 10560 10684 10566 10696
rect 10686 10684 10692 10696
rect 10744 10724 10750 10736
rect 13464 10724 13492 10764
rect 15105 10761 15117 10795
rect 15151 10792 15163 10795
rect 15194 10792 15200 10804
rect 15151 10764 15200 10792
rect 15151 10761 15163 10764
rect 15105 10755 15163 10761
rect 15194 10752 15200 10764
rect 15252 10792 15258 10804
rect 16022 10792 16028 10804
rect 15252 10764 16028 10792
rect 15252 10752 15258 10764
rect 16022 10752 16028 10764
rect 16080 10752 16086 10804
rect 17144 10764 18552 10792
rect 10744 10696 12112 10724
rect 13464 10696 14122 10724
rect 10744 10684 10750 10696
rect 10137 10659 10195 10665
rect 10137 10625 10149 10659
rect 10183 10625 10195 10659
rect 10137 10619 10195 10625
rect 7607 10560 9674 10588
rect 10152 10588 10180 10619
rect 10226 10616 10232 10668
rect 10284 10656 10290 10668
rect 10778 10656 10784 10668
rect 10284 10628 10784 10656
rect 10284 10616 10290 10628
rect 10778 10616 10784 10628
rect 10836 10616 10842 10668
rect 10873 10659 10931 10665
rect 10873 10625 10885 10659
rect 10919 10656 10931 10659
rect 11974 10656 11980 10668
rect 10919 10628 11980 10656
rect 10919 10625 10931 10628
rect 10873 10619 10931 10625
rect 11974 10616 11980 10628
rect 12032 10616 12038 10668
rect 12084 10665 12112 10696
rect 15286 10684 15292 10736
rect 15344 10724 15350 10736
rect 17144 10724 17172 10764
rect 15344 10696 17172 10724
rect 15344 10684 15350 10696
rect 17954 10684 17960 10736
rect 18012 10684 18018 10736
rect 18524 10724 18552 10764
rect 18598 10752 18604 10804
rect 18656 10792 18662 10804
rect 19334 10792 19340 10804
rect 18656 10764 19340 10792
rect 18656 10752 18662 10764
rect 19334 10752 19340 10764
rect 19392 10752 19398 10804
rect 20254 10792 20260 10804
rect 19904 10764 20260 10792
rect 19904 10724 19932 10764
rect 20254 10752 20260 10764
rect 20312 10752 20318 10804
rect 20438 10752 20444 10804
rect 20496 10792 20502 10804
rect 20496 10764 22094 10792
rect 20496 10752 20502 10764
rect 18524 10696 19932 10724
rect 12069 10659 12127 10665
rect 12069 10625 12081 10659
rect 12115 10625 12127 10659
rect 12069 10619 12127 10625
rect 12526 10616 12532 10668
rect 12584 10656 12590 10668
rect 12713 10659 12771 10665
rect 12713 10656 12725 10659
rect 12584 10628 12725 10656
rect 12584 10616 12590 10628
rect 12713 10625 12725 10628
rect 12759 10656 12771 10659
rect 13354 10656 13360 10668
rect 12759 10628 13216 10656
rect 13315 10628 13360 10656
rect 12759 10625 12771 10628
rect 12713 10619 12771 10625
rect 11422 10588 11428 10600
rect 10152 10560 11428 10588
rect 7607 10557 7619 10560
rect 7561 10551 7619 10557
rect 11422 10548 11428 10560
rect 11480 10588 11486 10600
rect 11698 10588 11704 10600
rect 11480 10560 11704 10588
rect 11480 10548 11486 10560
rect 11698 10548 11704 10560
rect 11756 10548 11762 10600
rect 13188 10588 13216 10628
rect 13354 10616 13360 10628
rect 13412 10616 13418 10668
rect 15838 10616 15844 10668
rect 15896 10656 15902 10668
rect 16114 10656 16120 10668
rect 15896 10628 16120 10656
rect 15896 10616 15902 10628
rect 16114 10616 16120 10628
rect 16172 10616 16178 10668
rect 13633 10591 13691 10597
rect 13188 10560 13492 10588
rect 8570 10480 8576 10532
rect 8628 10520 8634 10532
rect 10229 10523 10287 10529
rect 8628 10492 9996 10520
rect 8628 10480 8634 10492
rect 2685 10455 2743 10461
rect 2685 10421 2697 10455
rect 2731 10452 2743 10455
rect 9858 10452 9864 10464
rect 2731 10424 9864 10452
rect 2731 10421 2743 10424
rect 2685 10415 2743 10421
rect 9858 10412 9864 10424
rect 9916 10412 9922 10464
rect 9968 10452 9996 10492
rect 10229 10489 10241 10523
rect 10275 10520 10287 10523
rect 10275 10492 12296 10520
rect 10275 10489 10287 10492
rect 10229 10483 10287 10489
rect 10318 10452 10324 10464
rect 9968 10424 10324 10452
rect 10318 10412 10324 10424
rect 10376 10412 10382 10464
rect 12268 10452 12296 10492
rect 12710 10452 12716 10464
rect 12268 10424 12716 10452
rect 12710 10412 12716 10424
rect 12768 10412 12774 10464
rect 13464 10452 13492 10560
rect 13633 10557 13645 10591
rect 13679 10588 13691 10591
rect 16942 10588 16948 10600
rect 13679 10560 15884 10588
rect 16903 10560 16948 10588
rect 13679 10557 13691 10560
rect 13633 10551 13691 10557
rect 13722 10452 13728 10464
rect 13464 10424 13728 10452
rect 13722 10412 13728 10424
rect 13780 10412 13786 10464
rect 15856 10452 15884 10560
rect 16942 10548 16948 10560
rect 17000 10548 17006 10600
rect 17221 10591 17279 10597
rect 17221 10557 17233 10591
rect 17267 10588 17279 10591
rect 17862 10588 17868 10600
rect 17267 10560 17868 10588
rect 17267 10557 17279 10560
rect 17221 10551 17279 10557
rect 17862 10548 17868 10560
rect 17920 10548 17926 10600
rect 18524 10588 18552 10696
rect 19978 10684 19984 10736
rect 20036 10684 20042 10736
rect 19242 10656 19248 10668
rect 19203 10628 19248 10656
rect 19242 10616 19248 10628
rect 19300 10616 19306 10668
rect 18693 10591 18751 10597
rect 18693 10588 18705 10591
rect 18524 10560 18705 10588
rect 18693 10557 18705 10560
rect 18739 10557 18751 10591
rect 18693 10551 18751 10557
rect 18782 10548 18788 10600
rect 18840 10588 18846 10600
rect 19521 10591 19579 10597
rect 19521 10588 19533 10591
rect 18840 10560 19533 10588
rect 18840 10548 18846 10560
rect 19521 10557 19533 10560
rect 19567 10557 19579 10591
rect 19521 10551 19579 10557
rect 19610 10548 19616 10600
rect 19668 10588 19674 10600
rect 21818 10588 21824 10600
rect 19668 10560 21824 10588
rect 19668 10548 19674 10560
rect 21818 10548 21824 10560
rect 21876 10548 21882 10600
rect 18230 10480 18236 10532
rect 18288 10520 18294 10532
rect 22066 10520 22094 10764
rect 25498 10752 25504 10804
rect 25556 10792 25562 10804
rect 25593 10795 25651 10801
rect 25593 10792 25605 10795
rect 25556 10764 25605 10792
rect 25556 10752 25562 10764
rect 25593 10761 25605 10764
rect 25639 10761 25651 10795
rect 29270 10792 29276 10804
rect 29231 10764 29276 10792
rect 25593 10755 25651 10761
rect 29270 10752 29276 10764
rect 29328 10752 29334 10804
rect 35161 10795 35219 10801
rect 35161 10761 35173 10795
rect 35207 10792 35219 10795
rect 36906 10792 36912 10804
rect 35207 10764 36912 10792
rect 35207 10761 35219 10764
rect 35161 10755 35219 10761
rect 36906 10752 36912 10764
rect 36964 10752 36970 10804
rect 23750 10724 23756 10736
rect 23711 10696 23756 10724
rect 23750 10684 23756 10696
rect 23808 10684 23814 10736
rect 25958 10684 25964 10736
rect 26016 10724 26022 10736
rect 31754 10724 31760 10736
rect 26016 10696 31760 10724
rect 26016 10684 26022 10696
rect 31754 10684 31760 10696
rect 31812 10684 31818 10736
rect 22554 10656 22560 10668
rect 22515 10628 22560 10656
rect 22554 10616 22560 10628
rect 22612 10616 22618 10668
rect 25501 10659 25559 10665
rect 25501 10625 25513 10659
rect 25547 10625 25559 10659
rect 29454 10656 29460 10668
rect 29415 10628 29460 10656
rect 25501 10619 25559 10625
rect 23474 10548 23480 10600
rect 23532 10588 23538 10600
rect 23661 10591 23719 10597
rect 23661 10588 23673 10591
rect 23532 10560 23673 10588
rect 23532 10548 23538 10560
rect 23661 10557 23673 10560
rect 23707 10588 23719 10591
rect 23842 10588 23848 10600
rect 23707 10560 23848 10588
rect 23707 10557 23719 10560
rect 23661 10551 23719 10557
rect 23842 10548 23848 10560
rect 23900 10548 23906 10600
rect 23937 10591 23995 10597
rect 23937 10557 23949 10591
rect 23983 10557 23995 10591
rect 23937 10551 23995 10557
rect 23952 10520 23980 10551
rect 24946 10520 24952 10532
rect 18288 10492 18828 10520
rect 22066 10492 24952 10520
rect 18288 10480 18294 10492
rect 16114 10452 16120 10464
rect 15856 10424 16120 10452
rect 16114 10412 16120 10424
rect 16172 10452 16178 10464
rect 17678 10452 17684 10464
rect 16172 10424 17684 10452
rect 16172 10412 16178 10424
rect 17678 10412 17684 10424
rect 17736 10412 17742 10464
rect 18800 10452 18828 10492
rect 24946 10480 24952 10492
rect 25004 10480 25010 10532
rect 20993 10455 21051 10461
rect 20993 10452 21005 10455
rect 18800 10424 21005 10452
rect 20993 10421 21005 10424
rect 21039 10421 21051 10455
rect 20993 10415 21051 10421
rect 21910 10412 21916 10464
rect 21968 10452 21974 10464
rect 22649 10455 22707 10461
rect 22649 10452 22661 10455
rect 21968 10424 22661 10452
rect 21968 10412 21974 10424
rect 22649 10421 22661 10424
rect 22695 10421 22707 10455
rect 22649 10415 22707 10421
rect 22830 10412 22836 10464
rect 22888 10452 22894 10464
rect 25516 10452 25544 10619
rect 29454 10616 29460 10628
rect 29512 10616 29518 10668
rect 34514 10656 34520 10668
rect 34475 10628 34520 10656
rect 34514 10616 34520 10628
rect 34572 10616 34578 10668
rect 35345 10659 35403 10665
rect 35345 10625 35357 10659
rect 35391 10625 35403 10659
rect 38010 10656 38016 10668
rect 37971 10628 38016 10656
rect 35345 10619 35403 10625
rect 33134 10548 33140 10600
rect 33192 10588 33198 10600
rect 35360 10588 35388 10619
rect 38010 10616 38016 10628
rect 38068 10616 38074 10668
rect 33192 10560 35388 10588
rect 33192 10548 33198 10560
rect 22888 10424 25544 10452
rect 34333 10455 34391 10461
rect 22888 10412 22894 10424
rect 34333 10421 34345 10455
rect 34379 10452 34391 10455
rect 35526 10452 35532 10464
rect 34379 10424 35532 10452
rect 34379 10421 34391 10424
rect 34333 10415 34391 10421
rect 35526 10412 35532 10424
rect 35584 10412 35590 10464
rect 38194 10452 38200 10464
rect 38155 10424 38200 10452
rect 38194 10412 38200 10424
rect 38252 10412 38258 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 3973 10251 4031 10257
rect 3973 10217 3985 10251
rect 4019 10248 4031 10251
rect 8573 10251 8631 10257
rect 4019 10220 8248 10248
rect 4019 10217 4031 10220
rect 3973 10211 4031 10217
rect 2685 10183 2743 10189
rect 2685 10149 2697 10183
rect 2731 10180 2743 10183
rect 6454 10180 6460 10192
rect 2731 10152 6460 10180
rect 2731 10149 2743 10152
rect 2685 10143 2743 10149
rect 6454 10140 6460 10152
rect 6512 10140 6518 10192
rect 8220 10180 8248 10220
rect 8573 10217 8585 10251
rect 8619 10248 8631 10251
rect 9030 10248 9036 10260
rect 8619 10220 9036 10248
rect 8619 10217 8631 10220
rect 8573 10211 8631 10217
rect 9030 10208 9036 10220
rect 9088 10208 9094 10260
rect 9692 10220 11008 10248
rect 9692 10180 9720 10220
rect 8220 10152 9720 10180
rect 10980 10180 11008 10220
rect 11330 10208 11336 10260
rect 11388 10248 11394 10260
rect 11425 10251 11483 10257
rect 11425 10248 11437 10251
rect 11388 10220 11437 10248
rect 11388 10208 11394 10220
rect 11425 10217 11437 10220
rect 11471 10217 11483 10251
rect 11425 10211 11483 10217
rect 11698 10208 11704 10260
rect 11756 10248 11762 10260
rect 16022 10248 16028 10260
rect 11756 10220 16028 10248
rect 11756 10208 11762 10220
rect 16022 10208 16028 10220
rect 16080 10208 16086 10260
rect 18601 10251 18659 10257
rect 16132 10220 17356 10248
rect 11514 10180 11520 10192
rect 10980 10152 11520 10180
rect 11514 10140 11520 10152
rect 11572 10140 11578 10192
rect 13630 10180 13636 10192
rect 13591 10152 13636 10180
rect 13630 10140 13636 10152
rect 13688 10140 13694 10192
rect 13722 10140 13728 10192
rect 13780 10180 13786 10192
rect 16132 10180 16160 10220
rect 17328 10192 17356 10220
rect 18601 10217 18613 10251
rect 18647 10248 18659 10251
rect 23109 10251 23167 10257
rect 18647 10220 21680 10248
rect 18647 10217 18659 10220
rect 18601 10211 18659 10217
rect 13780 10152 16160 10180
rect 13780 10140 13786 10152
rect 17310 10140 17316 10192
rect 17368 10180 17374 10192
rect 17368 10152 18184 10180
rect 17368 10140 17374 10152
rect 3329 10115 3387 10121
rect 3329 10081 3341 10115
rect 3375 10112 3387 10115
rect 5534 10112 5540 10124
rect 3375 10084 5540 10112
rect 3375 10081 3387 10084
rect 3329 10075 3387 10081
rect 5534 10072 5540 10084
rect 5592 10072 5598 10124
rect 7101 10115 7159 10121
rect 7101 10081 7113 10115
rect 7147 10112 7159 10115
rect 15102 10112 15108 10124
rect 7147 10084 13584 10112
rect 7147 10081 7159 10084
rect 7101 10075 7159 10081
rect 1949 10047 2007 10053
rect 1949 10013 1961 10047
rect 1995 10044 2007 10047
rect 2593 10047 2651 10053
rect 2593 10044 2605 10047
rect 1995 10016 2605 10044
rect 1995 10013 2007 10016
rect 1949 10007 2007 10013
rect 2593 10013 2605 10016
rect 2639 10044 2651 10047
rect 2774 10044 2780 10056
rect 2639 10016 2780 10044
rect 2639 10013 2651 10016
rect 2593 10007 2651 10013
rect 2774 10004 2780 10016
rect 2832 10044 2838 10056
rect 3237 10047 3295 10053
rect 3237 10044 3249 10047
rect 2832 10016 3249 10044
rect 2832 10004 2838 10016
rect 3237 10013 3249 10016
rect 3283 10044 3295 10047
rect 4157 10047 4215 10053
rect 3283 10016 3924 10044
rect 3283 10013 3295 10016
rect 3237 10007 3295 10013
rect 3896 9988 3924 10016
rect 4157 10013 4169 10047
rect 4203 10044 4215 10047
rect 4798 10044 4804 10056
rect 4203 10016 4804 10044
rect 4203 10013 4215 10016
rect 4157 10007 4215 10013
rect 4798 10004 4804 10016
rect 4856 10004 4862 10056
rect 4982 10004 4988 10056
rect 5040 10044 5046 10056
rect 5442 10044 5448 10056
rect 5040 10016 5448 10044
rect 5040 10004 5046 10016
rect 5442 10004 5448 10016
rect 5500 10004 5506 10056
rect 5810 10004 5816 10056
rect 5868 10044 5874 10056
rect 6546 10044 6552 10056
rect 5868 10016 6552 10044
rect 5868 10004 5874 10016
rect 6546 10004 6552 10016
rect 6604 10004 6610 10056
rect 6822 10044 6828 10056
rect 6783 10016 6828 10044
rect 6822 10004 6828 10016
rect 6880 10004 6886 10056
rect 8570 10004 8576 10056
rect 8628 10044 8634 10056
rect 9490 10044 9496 10056
rect 8628 10016 9496 10044
rect 8628 10004 8634 10016
rect 9490 10004 9496 10016
rect 9548 10044 9554 10056
rect 9677 10047 9735 10053
rect 9677 10044 9689 10047
rect 9548 10016 9689 10044
rect 9548 10004 9554 10016
rect 9677 10013 9689 10016
rect 9723 10013 9735 10047
rect 11882 10044 11888 10056
rect 11843 10016 11888 10044
rect 9677 10007 9735 10013
rect 11882 10004 11888 10016
rect 11940 10004 11946 10056
rect 2041 9979 2099 9985
rect 2041 9945 2053 9979
rect 2087 9976 2099 9979
rect 2087 9948 2774 9976
rect 2087 9945 2099 9948
rect 2041 9939 2099 9945
rect 2746 9908 2774 9948
rect 3878 9936 3884 9988
rect 3936 9976 3942 9988
rect 5718 9976 5724 9988
rect 3936 9948 5724 9976
rect 3936 9936 3942 9948
rect 5718 9936 5724 9948
rect 5776 9976 5782 9988
rect 6086 9976 6092 9988
rect 5776 9948 6092 9976
rect 5776 9936 5782 9948
rect 6086 9936 6092 9948
rect 6144 9936 6150 9988
rect 7006 9936 7012 9988
rect 7064 9976 7070 9988
rect 9950 9976 9956 9988
rect 7064 9948 7590 9976
rect 9911 9948 9956 9976
rect 7064 9936 7070 9948
rect 9950 9936 9956 9948
rect 10008 9936 10014 9988
rect 10226 9936 10232 9988
rect 10284 9976 10290 9988
rect 12161 9979 12219 9985
rect 10284 9948 10442 9976
rect 10284 9936 10290 9948
rect 12161 9945 12173 9979
rect 12207 9976 12219 9979
rect 12207 9948 12434 9976
rect 12207 9945 12219 9948
rect 12161 9939 12219 9945
rect 4982 9908 4988 9920
rect 2746 9880 4988 9908
rect 4982 9868 4988 9880
rect 5040 9868 5046 9920
rect 5350 9868 5356 9920
rect 5408 9908 5414 9920
rect 9766 9908 9772 9920
rect 5408 9880 9772 9908
rect 5408 9868 5414 9880
rect 9766 9868 9772 9880
rect 9824 9868 9830 9920
rect 12406 9908 12434 9948
rect 12618 9936 12624 9988
rect 12676 9936 12682 9988
rect 13556 9976 13584 10084
rect 14936 10084 15108 10112
rect 14936 10053 14964 10084
rect 15102 10072 15108 10084
rect 15160 10112 15166 10124
rect 16298 10112 16304 10124
rect 15160 10084 16304 10112
rect 15160 10072 15166 10084
rect 16298 10072 16304 10084
rect 16356 10072 16362 10124
rect 16850 10072 16856 10124
rect 16908 10112 16914 10124
rect 16908 10084 17540 10112
rect 16908 10072 16914 10084
rect 14921 10047 14979 10053
rect 14921 10013 14933 10047
rect 14967 10013 14979 10047
rect 14921 10007 14979 10013
rect 15470 10004 15476 10056
rect 15528 10044 15534 10056
rect 16025 10047 16083 10053
rect 16025 10044 16037 10047
rect 15528 10016 16037 10044
rect 15528 10004 15534 10016
rect 16025 10013 16037 10016
rect 16071 10013 16083 10047
rect 17512 10044 17540 10084
rect 17862 10072 17868 10124
rect 17920 10112 17926 10124
rect 18049 10115 18107 10121
rect 18049 10112 18061 10115
rect 17920 10084 18061 10112
rect 17920 10072 17926 10084
rect 18049 10081 18061 10084
rect 18095 10081 18107 10115
rect 18156 10112 18184 10152
rect 18230 10140 18236 10192
rect 18288 10180 18294 10192
rect 19610 10180 19616 10192
rect 18288 10152 19616 10180
rect 18288 10140 18294 10152
rect 19610 10140 19616 10152
rect 19668 10140 19674 10192
rect 21652 10180 21680 10220
rect 23109 10217 23121 10251
rect 23155 10248 23167 10251
rect 23290 10248 23296 10260
rect 23155 10220 23296 10248
rect 23155 10217 23167 10220
rect 23109 10211 23167 10217
rect 23290 10208 23296 10220
rect 23348 10208 23354 10260
rect 37829 10251 37887 10257
rect 37829 10217 37841 10251
rect 37875 10248 37887 10251
rect 38010 10248 38016 10260
rect 37875 10220 38016 10248
rect 37875 10217 37887 10220
rect 37829 10211 37887 10217
rect 38010 10208 38016 10220
rect 38068 10208 38074 10260
rect 24026 10180 24032 10192
rect 21652 10152 24032 10180
rect 24026 10140 24032 10152
rect 24084 10140 24090 10192
rect 18156 10084 18644 10112
rect 18049 10075 18107 10081
rect 18509 10047 18567 10053
rect 18509 10044 18521 10047
rect 17512 10016 18521 10044
rect 16025 10007 16083 10013
rect 18509 10013 18521 10016
rect 18555 10013 18567 10047
rect 18509 10007 18567 10013
rect 15194 9976 15200 9988
rect 13556 9948 15200 9976
rect 15194 9936 15200 9948
rect 15252 9936 15258 9988
rect 16301 9979 16359 9985
rect 16301 9945 16313 9979
rect 16347 9945 16359 9979
rect 17586 9976 17592 9988
rect 17526 9948 17592 9976
rect 16301 9939 16359 9945
rect 13906 9908 13912 9920
rect 12406 9880 13912 9908
rect 13906 9868 13912 9880
rect 13964 9868 13970 9920
rect 15013 9911 15071 9917
rect 15013 9877 15025 9911
rect 15059 9908 15071 9911
rect 15286 9908 15292 9920
rect 15059 9880 15292 9908
rect 15059 9877 15071 9880
rect 15013 9871 15071 9877
rect 15286 9868 15292 9880
rect 15344 9868 15350 9920
rect 16316 9908 16344 9939
rect 17586 9936 17592 9948
rect 17644 9936 17650 9988
rect 18616 9976 18644 10084
rect 18966 10072 18972 10124
rect 19024 10112 19030 10124
rect 20162 10112 20168 10124
rect 19024 10084 20168 10112
rect 19024 10072 19030 10084
rect 20162 10072 20168 10084
rect 20220 10072 20226 10124
rect 20530 10072 20536 10124
rect 20588 10112 20594 10124
rect 21545 10115 21603 10121
rect 21545 10112 21557 10115
rect 20588 10084 21557 10112
rect 20588 10072 20594 10084
rect 21545 10081 21557 10084
rect 21591 10081 21603 10115
rect 21545 10075 21603 10081
rect 21818 10072 21824 10124
rect 21876 10112 21882 10124
rect 24670 10112 24676 10124
rect 21876 10084 22094 10112
rect 24631 10084 24676 10112
rect 21876 10072 21882 10084
rect 19334 10004 19340 10056
rect 19392 10044 19398 10056
rect 19797 10047 19855 10053
rect 19797 10044 19809 10047
rect 19392 10016 19809 10044
rect 19392 10004 19398 10016
rect 19797 10013 19809 10016
rect 19843 10013 19855 10047
rect 22066 10044 22094 10084
rect 24670 10072 24676 10084
rect 24728 10072 24734 10124
rect 23017 10047 23075 10053
rect 23017 10044 23029 10047
rect 22066 10016 23029 10044
rect 19797 10007 19855 10013
rect 23017 10013 23029 10016
rect 23063 10013 23075 10047
rect 23017 10007 23075 10013
rect 37458 10004 37464 10056
rect 37516 10044 37522 10056
rect 38013 10047 38071 10053
rect 38013 10044 38025 10047
rect 37516 10016 38025 10044
rect 37516 10004 37522 10016
rect 38013 10013 38025 10016
rect 38059 10013 38071 10047
rect 38013 10007 38071 10013
rect 19978 9976 19984 9988
rect 18616 9948 19984 9976
rect 19978 9936 19984 9948
rect 20036 9936 20042 9988
rect 20073 9979 20131 9985
rect 20073 9945 20085 9979
rect 20119 9976 20131 9979
rect 20162 9976 20168 9988
rect 20119 9948 20168 9976
rect 20119 9945 20131 9948
rect 20073 9939 20131 9945
rect 20162 9936 20168 9948
rect 20220 9936 20226 9988
rect 22738 9976 22744 9988
rect 21298 9948 22744 9976
rect 22738 9936 22744 9948
rect 22796 9936 22802 9988
rect 24762 9936 24768 9988
rect 24820 9976 24826 9988
rect 25685 9979 25743 9985
rect 24820 9948 24865 9976
rect 24820 9936 24826 9948
rect 25685 9945 25697 9979
rect 25731 9976 25743 9979
rect 25958 9976 25964 9988
rect 25731 9948 25964 9976
rect 25731 9945 25743 9948
rect 25685 9939 25743 9945
rect 25958 9936 25964 9948
rect 26016 9936 26022 9988
rect 18966 9908 18972 9920
rect 16316 9880 18972 9908
rect 18966 9868 18972 9880
rect 19024 9868 19030 9920
rect 20180 9908 20208 9936
rect 27154 9908 27160 9920
rect 20180 9880 27160 9908
rect 27154 9868 27160 9880
rect 27212 9868 27218 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 4522 9664 4528 9716
rect 4580 9704 4586 9716
rect 4580 9676 4625 9704
rect 4580 9664 4586 9676
rect 4798 9664 4804 9716
rect 4856 9704 4862 9716
rect 4856 9676 5488 9704
rect 4856 9664 4862 9676
rect 2222 9596 2228 9648
rect 2280 9636 2286 9648
rect 5460 9636 5488 9676
rect 5534 9664 5540 9716
rect 5592 9704 5598 9716
rect 9030 9704 9036 9716
rect 5592 9676 9036 9704
rect 5592 9664 5598 9676
rect 9030 9664 9036 9676
rect 9088 9664 9094 9716
rect 9582 9664 9588 9716
rect 9640 9704 9646 9716
rect 12526 9704 12532 9716
rect 9640 9676 12532 9704
rect 9640 9664 9646 9676
rect 12526 9664 12532 9676
rect 12584 9664 12590 9716
rect 13630 9704 13636 9716
rect 13004 9676 13636 9704
rect 2280 9608 4831 9636
rect 5460 9608 8510 9636
rect 2280 9596 2286 9608
rect 1673 9571 1731 9577
rect 1673 9537 1685 9571
rect 1719 9568 1731 9571
rect 2130 9568 2136 9580
rect 1719 9540 2136 9568
rect 1719 9537 1731 9540
rect 1673 9531 1731 9537
rect 2130 9528 2136 9540
rect 2188 9568 2194 9580
rect 2317 9571 2375 9577
rect 2317 9568 2329 9571
rect 2188 9540 2329 9568
rect 2188 9528 2194 9540
rect 2317 9537 2329 9540
rect 2363 9568 2375 9571
rect 2590 9568 2596 9580
rect 2363 9540 2596 9568
rect 2363 9537 2375 9540
rect 2317 9531 2375 9537
rect 2590 9528 2596 9540
rect 2648 9528 2654 9580
rect 3234 9568 3240 9580
rect 3195 9540 3240 9568
rect 3234 9528 3240 9540
rect 3292 9528 3298 9580
rect 3878 9568 3884 9580
rect 3839 9540 3884 9568
rect 3878 9528 3884 9540
rect 3936 9528 3942 9580
rect 4246 9528 4252 9580
rect 4304 9568 4310 9580
rect 4701 9571 4759 9577
rect 4304 9566 4660 9568
rect 4701 9566 4713 9571
rect 4304 9540 4713 9566
rect 4304 9528 4310 9540
rect 4632 9538 4713 9540
rect 4701 9537 4713 9538
rect 4747 9537 4759 9571
rect 4803 9568 4831 9608
rect 9490 9596 9496 9648
rect 9548 9636 9554 9648
rect 10965 9639 11023 9645
rect 10965 9636 10977 9639
rect 9548 9608 10977 9636
rect 9548 9596 9554 9608
rect 10965 9605 10977 9608
rect 11011 9605 11023 9639
rect 13004 9636 13032 9676
rect 13630 9664 13636 9676
rect 13688 9664 13694 9716
rect 15378 9664 15384 9716
rect 15436 9704 15442 9716
rect 22554 9704 22560 9716
rect 15436 9676 22560 9704
rect 15436 9664 15442 9676
rect 22554 9664 22560 9676
rect 22612 9664 22618 9716
rect 10965 9599 11023 9605
rect 11348 9608 13032 9636
rect 5353 9571 5411 9577
rect 5353 9568 5365 9571
rect 4803 9540 5365 9568
rect 4701 9531 4759 9537
rect 5353 9537 5365 9540
rect 5399 9537 5411 9571
rect 5353 9531 5411 9537
rect 10134 9528 10140 9580
rect 10192 9568 10198 9580
rect 10229 9571 10287 9577
rect 10229 9568 10241 9571
rect 10192 9540 10241 9568
rect 10192 9528 10198 9540
rect 10229 9537 10241 9540
rect 10275 9537 10287 9571
rect 10229 9531 10287 9537
rect 2409 9503 2467 9509
rect 2409 9469 2421 9503
rect 2455 9500 2467 9503
rect 3786 9500 3792 9512
rect 2455 9472 3792 9500
rect 2455 9469 2467 9472
rect 2409 9463 2467 9469
rect 3786 9460 3792 9472
rect 3844 9460 3850 9512
rect 4154 9460 4160 9512
rect 4212 9500 4218 9512
rect 5445 9503 5503 9509
rect 5445 9500 5457 9503
rect 4212 9472 5457 9500
rect 4212 9460 4218 9472
rect 5445 9469 5457 9472
rect 5491 9469 5503 9503
rect 5445 9463 5503 9469
rect 6822 9460 6828 9512
rect 6880 9500 6886 9512
rect 7745 9503 7803 9509
rect 7745 9500 7757 9503
rect 6880 9472 7757 9500
rect 6880 9460 6886 9472
rect 7745 9469 7757 9472
rect 7791 9469 7803 9503
rect 7745 9463 7803 9469
rect 8021 9503 8079 9509
rect 8021 9469 8033 9503
rect 8067 9500 8079 9503
rect 11348 9500 11376 9608
rect 13078 9596 13084 9648
rect 13136 9596 13142 9648
rect 14366 9596 14372 9648
rect 14424 9636 14430 9648
rect 14734 9636 14740 9648
rect 14424 9608 14740 9636
rect 14424 9596 14430 9608
rect 14734 9596 14740 9608
rect 14792 9596 14798 9648
rect 15470 9636 15476 9648
rect 15431 9608 15476 9636
rect 15470 9596 15476 9608
rect 15528 9596 15534 9648
rect 17770 9636 17776 9648
rect 15856 9608 17776 9636
rect 11701 9571 11759 9577
rect 11701 9537 11713 9571
rect 11747 9568 11759 9571
rect 12250 9568 12256 9580
rect 11747 9540 12256 9568
rect 11747 9537 11759 9540
rect 11701 9531 11759 9537
rect 12250 9528 12256 9540
rect 12308 9528 12314 9580
rect 14642 9568 14648 9580
rect 14603 9540 14648 9568
rect 14642 9528 14648 9540
rect 14700 9528 14706 9580
rect 15010 9528 15016 9580
rect 15068 9568 15074 9580
rect 15856 9568 15884 9608
rect 17770 9596 17776 9608
rect 17828 9596 17834 9648
rect 19150 9636 19156 9648
rect 18722 9608 19156 9636
rect 19150 9596 19156 9608
rect 19208 9596 19214 9648
rect 23658 9596 23664 9648
rect 23716 9636 23722 9648
rect 23753 9639 23811 9645
rect 23753 9636 23765 9639
rect 23716 9608 23765 9636
rect 23716 9596 23722 9608
rect 23753 9605 23765 9608
rect 23799 9605 23811 9639
rect 23753 9599 23811 9605
rect 30193 9639 30251 9645
rect 30193 9605 30205 9639
rect 30239 9636 30251 9639
rect 33134 9636 33140 9648
rect 30239 9608 33140 9636
rect 30239 9605 30251 9608
rect 30193 9599 30251 9605
rect 33134 9596 33140 9608
rect 33192 9596 33198 9648
rect 16022 9568 16028 9580
rect 15068 9540 15884 9568
rect 15983 9540 16028 9568
rect 15068 9528 15074 9540
rect 16022 9528 16028 9540
rect 16080 9528 16086 9580
rect 16942 9528 16948 9580
rect 17000 9568 17006 9580
rect 17221 9571 17279 9577
rect 17221 9568 17233 9571
rect 17000 9540 17233 9568
rect 17000 9528 17006 9540
rect 17221 9537 17233 9540
rect 17267 9537 17279 9571
rect 30101 9571 30159 9577
rect 20838 9540 22094 9568
rect 17221 9531 17279 9537
rect 8067 9472 11376 9500
rect 8067 9469 8079 9472
rect 8021 9463 8079 9469
rect 11882 9460 11888 9512
rect 11940 9500 11946 9512
rect 12342 9500 12348 9512
rect 11940 9472 12348 9500
rect 11940 9460 11946 9472
rect 12342 9460 12348 9472
rect 12400 9460 12406 9512
rect 12621 9503 12679 9509
rect 12621 9469 12633 9503
rect 12667 9500 12679 9503
rect 16206 9500 16212 9512
rect 12667 9472 16212 9500
rect 12667 9469 12679 9472
rect 12621 9463 12679 9469
rect 16206 9460 16212 9472
rect 16264 9460 16270 9512
rect 17497 9503 17555 9509
rect 17497 9469 17509 9503
rect 17543 9500 17555 9503
rect 18506 9500 18512 9512
rect 17543 9472 18512 9500
rect 17543 9469 17555 9472
rect 17497 9463 17555 9469
rect 18506 9460 18512 9472
rect 18564 9460 18570 9512
rect 18966 9500 18972 9512
rect 18927 9472 18972 9500
rect 18966 9460 18972 9472
rect 19024 9460 19030 9512
rect 19334 9460 19340 9512
rect 19392 9500 19398 9512
rect 19429 9503 19487 9509
rect 19429 9500 19441 9503
rect 19392 9472 19441 9500
rect 19392 9460 19398 9472
rect 19429 9469 19441 9472
rect 19475 9469 19487 9503
rect 19429 9463 19487 9469
rect 19705 9503 19763 9509
rect 19705 9469 19717 9503
rect 19751 9500 19763 9503
rect 20714 9500 20720 9512
rect 19751 9472 20720 9500
rect 19751 9469 19763 9472
rect 19705 9463 19763 9469
rect 20714 9460 20720 9472
rect 20772 9460 20778 9512
rect 21082 9460 21088 9512
rect 21140 9500 21146 9512
rect 21177 9503 21235 9509
rect 21177 9500 21189 9503
rect 21140 9472 21189 9500
rect 21140 9460 21146 9472
rect 21177 9469 21189 9472
rect 21223 9469 21235 9503
rect 21177 9463 21235 9469
rect 3326 9432 3332 9444
rect 3287 9404 3332 9432
rect 3326 9392 3332 9404
rect 3384 9392 3390 9444
rect 3973 9435 4031 9441
rect 3973 9401 3985 9435
rect 4019 9432 4031 9435
rect 5626 9432 5632 9444
rect 4019 9404 5632 9432
rect 4019 9401 4031 9404
rect 3973 9395 4031 9401
rect 5626 9392 5632 9404
rect 5684 9392 5690 9444
rect 15102 9432 15108 9444
rect 13740 9404 15108 9432
rect 1765 9367 1823 9373
rect 1765 9333 1777 9367
rect 1811 9364 1823 9367
rect 5810 9364 5816 9376
rect 1811 9336 5816 9364
rect 1811 9333 1823 9336
rect 1765 9327 1823 9333
rect 5810 9324 5816 9336
rect 5868 9324 5874 9376
rect 6914 9324 6920 9376
rect 6972 9364 6978 9376
rect 9306 9364 9312 9376
rect 6972 9336 9312 9364
rect 6972 9324 6978 9336
rect 9306 9324 9312 9336
rect 9364 9364 9370 9376
rect 9493 9367 9551 9373
rect 9493 9364 9505 9367
rect 9364 9336 9505 9364
rect 9364 9324 9370 9336
rect 9493 9333 9505 9336
rect 9539 9333 9551 9367
rect 9493 9327 9551 9333
rect 11793 9367 11851 9373
rect 11793 9333 11805 9367
rect 11839 9364 11851 9367
rect 13740 9364 13768 9404
rect 15102 9392 15108 9404
rect 15160 9392 15166 9444
rect 22066 9432 22094 9540
rect 30101 9537 30113 9571
rect 30147 9568 30159 9571
rect 30374 9568 30380 9580
rect 30147 9540 30380 9568
rect 30147 9537 30159 9540
rect 30101 9531 30159 9537
rect 30374 9528 30380 9540
rect 30432 9528 30438 9580
rect 30834 9528 30840 9580
rect 30892 9568 30898 9580
rect 30929 9571 30987 9577
rect 30929 9568 30941 9571
rect 30892 9540 30941 9568
rect 30892 9528 30898 9540
rect 30929 9537 30941 9540
rect 30975 9537 30987 9571
rect 30929 9531 30987 9537
rect 31573 9571 31631 9577
rect 31573 9537 31585 9571
rect 31619 9537 31631 9571
rect 31573 9531 31631 9537
rect 23661 9503 23719 9509
rect 23661 9469 23673 9503
rect 23707 9500 23719 9503
rect 23934 9500 23940 9512
rect 23707 9472 23940 9500
rect 23707 9469 23719 9472
rect 23661 9463 23719 9469
rect 23934 9460 23940 9472
rect 23992 9460 23998 9512
rect 24026 9460 24032 9512
rect 24084 9500 24090 9512
rect 24084 9472 24129 9500
rect 24084 9460 24090 9472
rect 29270 9460 29276 9512
rect 29328 9500 29334 9512
rect 29365 9503 29423 9509
rect 29365 9500 29377 9503
rect 29328 9472 29377 9500
rect 29328 9460 29334 9472
rect 29365 9469 29377 9472
rect 29411 9469 29423 9503
rect 31588 9500 31616 9531
rect 29365 9463 29423 9469
rect 30760 9472 31616 9500
rect 25774 9432 25780 9444
rect 22066 9404 25780 9432
rect 25774 9392 25780 9404
rect 25832 9392 25838 9444
rect 30760 9441 30788 9472
rect 30745 9435 30803 9441
rect 30745 9401 30757 9435
rect 30791 9401 30803 9435
rect 30745 9395 30803 9401
rect 14090 9364 14096 9376
rect 11839 9336 13768 9364
rect 14051 9336 14096 9364
rect 11839 9333 11851 9336
rect 11793 9327 11851 9333
rect 14090 9324 14096 9336
rect 14148 9324 14154 9376
rect 15010 9324 15016 9376
rect 15068 9364 15074 9376
rect 16117 9367 16175 9373
rect 16117 9364 16129 9367
rect 15068 9336 16129 9364
rect 15068 9324 15074 9336
rect 16117 9333 16129 9336
rect 16163 9333 16175 9367
rect 16117 9327 16175 9333
rect 19242 9324 19248 9376
rect 19300 9364 19306 9376
rect 20898 9364 20904 9376
rect 19300 9336 20904 9364
rect 19300 9324 19306 9336
rect 20898 9324 20904 9336
rect 20956 9324 20962 9376
rect 29454 9324 29460 9376
rect 29512 9364 29518 9376
rect 31389 9367 31447 9373
rect 31389 9364 31401 9367
rect 29512 9336 31401 9364
rect 29512 9324 29518 9336
rect 31389 9333 31401 9336
rect 31435 9333 31447 9367
rect 31389 9327 31447 9333
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 2314 9120 2320 9172
rect 2372 9160 2378 9172
rect 2372 9132 4384 9160
rect 2372 9120 2378 9132
rect 2590 9052 2596 9104
rect 2648 9092 2654 9104
rect 4157 9095 4215 9101
rect 4157 9092 4169 9095
rect 2648 9064 4169 9092
rect 2648 9052 2654 9064
rect 4157 9061 4169 9064
rect 4203 9061 4215 9095
rect 4157 9055 4215 9061
rect 1596 8996 3740 9024
rect 1596 8965 1624 8996
rect 1581 8959 1639 8965
rect 1581 8925 1593 8959
rect 1627 8925 1639 8959
rect 1581 8919 1639 8925
rect 2317 8959 2375 8965
rect 2317 8925 2329 8959
rect 2363 8956 2375 8959
rect 2958 8956 2964 8968
rect 2363 8928 2964 8956
rect 2363 8925 2375 8928
rect 2317 8919 2375 8925
rect 2958 8916 2964 8928
rect 3016 8916 3022 8968
rect 3234 8956 3240 8968
rect 3195 8928 3240 8956
rect 3234 8916 3240 8928
rect 3292 8916 3298 8968
rect 2409 8891 2467 8897
rect 2409 8857 2421 8891
rect 2455 8888 2467 8891
rect 3712 8888 3740 8996
rect 4356 8965 4384 9132
rect 4522 9120 4528 9172
rect 4580 9160 4586 9172
rect 6914 9160 6920 9172
rect 4580 9132 6920 9160
rect 4580 9120 4586 9132
rect 6914 9120 6920 9132
rect 6972 9120 6978 9172
rect 7088 9163 7146 9169
rect 7088 9129 7100 9163
rect 7134 9160 7146 9163
rect 7834 9160 7840 9172
rect 7134 9132 7840 9160
rect 7134 9129 7146 9132
rect 7088 9123 7146 9129
rect 7834 9120 7840 9132
rect 7892 9120 7898 9172
rect 8404 9132 10456 9160
rect 8404 9104 8432 9132
rect 8386 9052 8392 9104
rect 8444 9052 8450 9104
rect 8846 9052 8852 9104
rect 8904 9092 8910 9104
rect 10428 9092 10456 9132
rect 10594 9120 10600 9172
rect 10652 9160 10658 9172
rect 10873 9163 10931 9169
rect 10873 9160 10885 9163
rect 10652 9132 10885 9160
rect 10652 9120 10658 9132
rect 10873 9129 10885 9132
rect 10919 9129 10931 9163
rect 14090 9160 14096 9172
rect 10873 9123 10931 9129
rect 10980 9132 14096 9160
rect 10980 9092 11008 9132
rect 14090 9120 14096 9132
rect 14148 9120 14154 9172
rect 14274 9120 14280 9172
rect 14332 9160 14338 9172
rect 14332 9132 15700 9160
rect 14332 9120 14338 9132
rect 8904 9064 9260 9092
rect 10428 9064 11008 9092
rect 13081 9095 13139 9101
rect 8904 9052 8910 9064
rect 9125 9027 9183 9033
rect 9125 9024 9137 9027
rect 4724 8996 5120 9024
rect 4341 8959 4399 8965
rect 4341 8925 4353 8959
rect 4387 8925 4399 8959
rect 4341 8919 4399 8925
rect 4614 8888 4620 8900
rect 2455 8860 3648 8888
rect 3712 8860 4620 8888
rect 2455 8857 2467 8860
rect 2409 8851 2467 8857
rect 1762 8820 1768 8832
rect 1723 8792 1768 8820
rect 1762 8780 1768 8792
rect 1820 8780 1826 8832
rect 2866 8780 2872 8832
rect 2924 8820 2930 8832
rect 3053 8823 3111 8829
rect 3053 8820 3065 8823
rect 2924 8792 3065 8820
rect 2924 8780 2930 8792
rect 3053 8789 3065 8792
rect 3099 8789 3111 8823
rect 3620 8820 3648 8860
rect 4614 8848 4620 8860
rect 4672 8848 4678 8900
rect 4724 8820 4752 8996
rect 4985 8959 5043 8965
rect 4985 8925 4997 8959
rect 5031 8925 5043 8959
rect 4985 8919 5043 8925
rect 3620 8792 4752 8820
rect 3053 8783 3111 8789
rect 4798 8780 4804 8832
rect 4856 8820 4862 8832
rect 5000 8820 5028 8919
rect 5092 8888 5120 8996
rect 6840 8996 9137 9024
rect 6840 8968 6868 8996
rect 9125 8993 9137 8996
rect 9171 8993 9183 9027
rect 9232 9024 9260 9064
rect 13081 9061 13093 9095
rect 13127 9092 13139 9095
rect 13906 9092 13912 9104
rect 13127 9064 13912 9092
rect 13127 9061 13139 9064
rect 13081 9055 13139 9061
rect 13906 9052 13912 9064
rect 13964 9052 13970 9104
rect 15672 9092 15700 9132
rect 16482 9120 16488 9172
rect 16540 9160 16546 9172
rect 21358 9160 21364 9172
rect 16540 9132 21364 9160
rect 16540 9120 16546 9132
rect 21358 9120 21364 9132
rect 21416 9120 21422 9172
rect 22738 9120 22744 9172
rect 22796 9160 22802 9172
rect 23017 9163 23075 9169
rect 23017 9160 23029 9163
rect 22796 9132 23029 9160
rect 22796 9120 22802 9132
rect 23017 9129 23029 9132
rect 23063 9129 23075 9163
rect 23658 9160 23664 9172
rect 23619 9132 23664 9160
rect 23017 9123 23075 9129
rect 23658 9120 23664 9132
rect 23716 9120 23722 9172
rect 15672 9064 19748 9092
rect 9398 9024 9404 9036
rect 9232 8996 9404 9024
rect 9125 8987 9183 8993
rect 9398 8984 9404 8996
rect 9456 8984 9462 9036
rect 9490 8984 9496 9036
rect 9548 9024 9554 9036
rect 11238 9024 11244 9036
rect 9548 8996 11244 9024
rect 9548 8984 9554 8996
rect 11238 8984 11244 8996
rect 11296 8984 11302 9036
rect 11333 9027 11391 9033
rect 11333 8993 11345 9027
rect 11379 9024 11391 9027
rect 12342 9024 12348 9036
rect 11379 8996 12348 9024
rect 11379 8993 11391 8996
rect 11333 8987 11391 8993
rect 12342 8984 12348 8996
rect 12400 9024 12406 9036
rect 12894 9024 12900 9036
rect 12400 8996 12900 9024
rect 12400 8984 12406 8996
rect 12894 8984 12900 8996
rect 12952 9024 12958 9036
rect 14369 9027 14427 9033
rect 14369 9024 14381 9027
rect 12952 8996 14381 9024
rect 12952 8984 12958 8996
rect 14369 8993 14381 8996
rect 14415 9024 14427 9027
rect 15378 9024 15384 9036
rect 14415 8996 15384 9024
rect 14415 8993 14427 8996
rect 14369 8987 14427 8993
rect 15378 8984 15384 8996
rect 15436 8984 15442 9036
rect 16850 8984 16856 9036
rect 16908 9024 16914 9036
rect 18693 9027 18751 9033
rect 18693 9024 18705 9027
rect 16908 8996 18705 9024
rect 16908 8984 16914 8996
rect 18693 8993 18705 8996
rect 18739 9024 18751 9027
rect 19334 9024 19340 9036
rect 18739 8996 19340 9024
rect 18739 8993 18751 8996
rect 18693 8987 18751 8993
rect 19334 8984 19340 8996
rect 19392 9024 19398 9036
rect 19613 9027 19671 9033
rect 19613 9024 19625 9027
rect 19392 8996 19625 9024
rect 19392 8984 19398 8996
rect 19613 8993 19625 8996
rect 19659 8993 19671 9027
rect 19720 9024 19748 9064
rect 20898 9052 20904 9104
rect 20956 9092 20962 9104
rect 25682 9092 25688 9104
rect 20956 9064 25688 9092
rect 20956 9052 20962 9064
rect 25682 9052 25688 9064
rect 25740 9052 25746 9104
rect 20254 9024 20260 9036
rect 19720 8996 20260 9024
rect 19613 8987 19671 8993
rect 20254 8984 20260 8996
rect 20312 8984 20318 9036
rect 20346 8984 20352 9036
rect 20404 9024 20410 9036
rect 29917 9027 29975 9033
rect 20404 8996 29868 9024
rect 20404 8984 20410 8996
rect 5166 8916 5172 8968
rect 5224 8956 5230 8968
rect 6822 8956 6828 8968
rect 5224 8928 6408 8956
rect 6783 8928 6828 8956
rect 5224 8916 5230 8928
rect 5258 8888 5264 8900
rect 5092 8860 5264 8888
rect 5258 8848 5264 8860
rect 5316 8848 5322 8900
rect 5445 8891 5503 8897
rect 5445 8857 5457 8891
rect 5491 8857 5503 8891
rect 6270 8888 6276 8900
rect 6231 8860 6276 8888
rect 5445 8851 5503 8857
rect 5166 8820 5172 8832
rect 4856 8792 4901 8820
rect 5000 8792 5172 8820
rect 4856 8780 4862 8792
rect 5166 8780 5172 8792
rect 5224 8780 5230 8832
rect 5460 8820 5488 8851
rect 6270 8848 6276 8860
rect 6328 8848 6334 8900
rect 6380 8888 6408 8928
rect 6822 8916 6828 8928
rect 6880 8916 6886 8968
rect 8478 8916 8484 8968
rect 8536 8956 8542 8968
rect 8846 8956 8852 8968
rect 8536 8928 8852 8956
rect 8536 8916 8542 8928
rect 8846 8916 8852 8928
rect 8904 8916 8910 8968
rect 12710 8916 12716 8968
rect 12768 8916 12774 8968
rect 16574 8956 16580 8968
rect 16535 8928 16580 8956
rect 16574 8916 16580 8928
rect 16632 8916 16638 8968
rect 19242 8916 19248 8968
rect 19300 8956 19306 8968
rect 21637 8959 21695 8965
rect 19300 8928 19656 8956
rect 19300 8916 19306 8928
rect 9306 8888 9312 8900
rect 6380 8860 7590 8888
rect 8404 8860 9312 8888
rect 7190 8820 7196 8832
rect 5460 8792 7196 8820
rect 7190 8780 7196 8792
rect 7248 8780 7254 8832
rect 7742 8780 7748 8832
rect 7800 8820 7806 8832
rect 8404 8820 8432 8860
rect 9306 8848 9312 8860
rect 9364 8848 9370 8900
rect 9398 8848 9404 8900
rect 9456 8888 9462 8900
rect 11609 8891 11667 8897
rect 9456 8860 9890 8888
rect 9456 8848 9462 8860
rect 11609 8857 11621 8891
rect 11655 8857 11667 8891
rect 11609 8851 11667 8857
rect 7800 8792 8432 8820
rect 8573 8823 8631 8829
rect 7800 8780 7806 8792
rect 8573 8789 8585 8823
rect 8619 8820 8631 8823
rect 9582 8820 9588 8832
rect 8619 8792 9588 8820
rect 8619 8789 8631 8792
rect 8573 8783 8631 8789
rect 9582 8780 9588 8792
rect 9640 8780 9646 8832
rect 9766 8780 9772 8832
rect 9824 8820 9830 8832
rect 10870 8820 10876 8832
rect 9824 8792 10876 8820
rect 9824 8780 9830 8792
rect 10870 8780 10876 8792
rect 10928 8780 10934 8832
rect 11624 8820 11652 8851
rect 14182 8848 14188 8900
rect 14240 8888 14246 8900
rect 14645 8891 14703 8897
rect 14645 8888 14657 8891
rect 14240 8860 14657 8888
rect 14240 8848 14246 8860
rect 14645 8857 14657 8860
rect 14691 8857 14703 8891
rect 14645 8851 14703 8857
rect 15102 8848 15108 8900
rect 15160 8848 15166 8900
rect 17954 8888 17960 8900
rect 17915 8860 17960 8888
rect 17954 8848 17960 8860
rect 18012 8888 18018 8900
rect 19426 8888 19432 8900
rect 18012 8860 19432 8888
rect 18012 8848 18018 8860
rect 19426 8848 19432 8860
rect 19484 8848 19490 8900
rect 19628 8888 19656 8928
rect 21637 8925 21649 8959
rect 21683 8956 21695 8959
rect 21726 8956 21732 8968
rect 21683 8928 21732 8956
rect 21683 8925 21695 8928
rect 21637 8919 21695 8925
rect 21726 8916 21732 8928
rect 21784 8916 21790 8968
rect 22925 8959 22983 8965
rect 22925 8925 22937 8959
rect 22971 8956 22983 8959
rect 23014 8956 23020 8968
rect 22971 8928 23020 8956
rect 22971 8925 22983 8928
rect 22925 8919 22983 8925
rect 19889 8891 19947 8897
rect 19889 8888 19901 8891
rect 19628 8860 19901 8888
rect 19889 8857 19901 8860
rect 19935 8857 19947 8891
rect 21174 8888 21180 8900
rect 21114 8860 21180 8888
rect 19889 8851 19947 8857
rect 21174 8848 21180 8860
rect 21232 8848 21238 8900
rect 12986 8820 12992 8832
rect 11624 8792 12992 8820
rect 12986 8780 12992 8792
rect 13044 8780 13050 8832
rect 13170 8780 13176 8832
rect 13228 8820 13234 8832
rect 16117 8823 16175 8829
rect 16117 8820 16129 8823
rect 13228 8792 16129 8820
rect 13228 8780 13234 8792
rect 16117 8789 16129 8792
rect 16163 8789 16175 8823
rect 16666 8820 16672 8832
rect 16627 8792 16672 8820
rect 16117 8783 16175 8789
rect 16666 8780 16672 8792
rect 16724 8780 16730 8832
rect 19444 8820 19472 8848
rect 20622 8820 20628 8832
rect 19444 8792 20628 8820
rect 20622 8780 20628 8792
rect 20680 8780 20686 8832
rect 20714 8780 20720 8832
rect 20772 8820 20778 8832
rect 21818 8820 21824 8832
rect 20772 8792 21824 8820
rect 20772 8780 20778 8792
rect 21818 8780 21824 8792
rect 21876 8780 21882 8832
rect 22940 8820 22968 8919
rect 23014 8916 23020 8928
rect 23072 8916 23078 8968
rect 23474 8916 23480 8968
rect 23532 8956 23538 8968
rect 23569 8959 23627 8965
rect 23569 8956 23581 8959
rect 23532 8928 23581 8956
rect 23532 8916 23538 8928
rect 23569 8925 23581 8928
rect 23615 8925 23627 8959
rect 23569 8919 23627 8925
rect 28629 8959 28687 8965
rect 28629 8925 28641 8959
rect 28675 8956 28687 8959
rect 29086 8956 29092 8968
rect 28675 8928 29092 8956
rect 28675 8925 28687 8928
rect 28629 8919 28687 8925
rect 29086 8916 29092 8928
rect 29144 8916 29150 8968
rect 29733 8959 29791 8965
rect 29733 8925 29745 8959
rect 29779 8925 29791 8959
rect 29840 8956 29868 8996
rect 29917 8993 29929 9027
rect 29963 9024 29975 9027
rect 30929 9027 30987 9033
rect 30929 9024 30941 9027
rect 29963 8996 30941 9024
rect 29963 8993 29975 8996
rect 29917 8987 29975 8993
rect 30929 8993 30941 8996
rect 30975 8993 30987 9027
rect 30929 8987 30987 8993
rect 30834 8956 30840 8968
rect 29840 8928 30840 8956
rect 29733 8919 29791 8925
rect 24946 8888 24952 8900
rect 24907 8860 24952 8888
rect 24946 8848 24952 8860
rect 25004 8848 25010 8900
rect 25038 8848 25044 8900
rect 25096 8888 25102 8900
rect 25958 8888 25964 8900
rect 25096 8860 25141 8888
rect 25700 8860 25964 8888
rect 25096 8848 25102 8860
rect 25700 8832 25728 8860
rect 25958 8848 25964 8860
rect 26016 8848 26022 8900
rect 26694 8848 26700 8900
rect 26752 8888 26758 8900
rect 29748 8888 29776 8919
rect 30834 8916 30840 8928
rect 30892 8916 30898 8968
rect 38286 8956 38292 8968
rect 38247 8928 38292 8956
rect 38286 8916 38292 8928
rect 38344 8916 38350 8968
rect 26752 8860 29776 8888
rect 26752 8848 26758 8860
rect 25590 8820 25596 8832
rect 22940 8792 25596 8820
rect 25590 8780 25596 8792
rect 25648 8780 25654 8832
rect 25682 8780 25688 8832
rect 25740 8780 25746 8832
rect 28721 8823 28779 8829
rect 28721 8789 28733 8823
rect 28767 8820 28779 8823
rect 30190 8820 30196 8832
rect 28767 8792 30196 8820
rect 28767 8789 28779 8792
rect 28721 8783 28779 8789
rect 30190 8780 30196 8792
rect 30248 8780 30254 8832
rect 30374 8820 30380 8832
rect 30335 8792 30380 8820
rect 30374 8780 30380 8792
rect 30432 8780 30438 8832
rect 38102 8820 38108 8832
rect 38063 8792 38108 8820
rect 38102 8780 38108 8792
rect 38160 8780 38166 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 1581 8619 1639 8625
rect 1581 8585 1593 8619
rect 1627 8616 1639 8619
rect 1854 8616 1860 8628
rect 1627 8588 1860 8616
rect 1627 8585 1639 8588
rect 1581 8579 1639 8585
rect 1854 8576 1860 8588
rect 1912 8576 1918 8628
rect 2222 8616 2228 8628
rect 2183 8588 2228 8616
rect 2222 8576 2228 8588
rect 2280 8576 2286 8628
rect 6822 8616 6828 8628
rect 4264 8588 6828 8616
rect 1394 8440 1400 8492
rect 1452 8480 1458 8492
rect 1765 8483 1823 8489
rect 1765 8480 1777 8483
rect 1452 8452 1777 8480
rect 1452 8440 1458 8452
rect 1765 8449 1777 8452
rect 1811 8449 1823 8483
rect 1765 8443 1823 8449
rect 1854 8440 1860 8492
rect 1912 8480 1918 8492
rect 2409 8483 2467 8489
rect 2409 8480 2421 8483
rect 1912 8452 2421 8480
rect 1912 8440 1918 8452
rect 2409 8449 2421 8452
rect 2455 8449 2467 8483
rect 3050 8480 3056 8492
rect 3011 8452 3056 8480
rect 2409 8443 2467 8449
rect 3050 8440 3056 8452
rect 3108 8440 3114 8492
rect 3789 8483 3847 8489
rect 3789 8449 3801 8483
rect 3835 8480 3847 8483
rect 3878 8480 3884 8492
rect 3835 8452 3884 8480
rect 3835 8449 3847 8452
rect 3789 8443 3847 8449
rect 3878 8440 3884 8452
rect 3936 8440 3942 8492
rect 4264 8489 4292 8588
rect 6822 8576 6828 8588
rect 6880 8616 6886 8628
rect 10134 8616 10140 8628
rect 6880 8588 7972 8616
rect 6880 8576 6886 8588
rect 4522 8548 4528 8560
rect 4483 8520 4528 8548
rect 4522 8508 4528 8520
rect 4580 8508 4586 8560
rect 5534 8508 5540 8560
rect 5592 8508 5598 8560
rect 6638 8548 6644 8560
rect 6599 8520 6644 8548
rect 6638 8508 6644 8520
rect 6696 8508 6702 8560
rect 7944 8557 7972 8588
rect 9048 8588 10140 8616
rect 7929 8551 7987 8557
rect 7929 8517 7941 8551
rect 7975 8517 7987 8551
rect 9048 8548 9076 8588
rect 10134 8576 10140 8588
rect 10192 8576 10198 8628
rect 13354 8576 13360 8628
rect 13412 8616 13418 8628
rect 14642 8616 14648 8628
rect 13412 8588 14648 8616
rect 13412 8576 13418 8588
rect 14642 8576 14648 8588
rect 14700 8616 14706 8628
rect 17954 8616 17960 8628
rect 14700 8588 17960 8616
rect 14700 8576 14706 8588
rect 7929 8511 7987 8517
rect 8588 8520 9076 8548
rect 4249 8483 4307 8489
rect 4249 8449 4261 8483
rect 4295 8449 4307 8483
rect 4249 8443 4307 8449
rect 6549 8483 6607 8489
rect 6549 8449 6561 8483
rect 6595 8449 6607 8483
rect 7190 8480 7196 8492
rect 7103 8452 7196 8480
rect 6549 8443 6607 8449
rect 6564 8412 6592 8443
rect 7190 8440 7196 8452
rect 7248 8480 7254 8492
rect 8588 8480 8616 8520
rect 9306 8508 9312 8560
rect 9364 8508 9370 8560
rect 12342 8548 12348 8560
rect 12303 8520 12348 8548
rect 12342 8508 12348 8520
rect 12400 8508 12406 8560
rect 13170 8508 13176 8560
rect 13228 8548 13234 8560
rect 13228 8520 13273 8548
rect 13228 8508 13234 8520
rect 13630 8508 13636 8560
rect 13688 8508 13694 8560
rect 14921 8551 14979 8557
rect 14921 8517 14933 8551
rect 14967 8548 14979 8551
rect 15102 8548 15108 8560
rect 14967 8520 15108 8548
rect 14967 8517 14979 8520
rect 14921 8511 14979 8517
rect 15102 8508 15108 8520
rect 15160 8508 15166 8560
rect 15396 8557 15424 8588
rect 17954 8576 17960 8588
rect 18012 8576 18018 8628
rect 18984 8588 21128 8616
rect 15381 8551 15439 8557
rect 15381 8517 15393 8551
rect 15427 8517 15439 8551
rect 17126 8548 17132 8560
rect 17087 8520 17132 8548
rect 15381 8511 15439 8517
rect 17126 8508 17132 8520
rect 17184 8508 17190 8560
rect 18984 8548 19012 8588
rect 19334 8548 19340 8560
rect 18354 8520 19012 8548
rect 19076 8520 19340 8548
rect 7248 8452 8616 8480
rect 7248 8440 7254 8452
rect 10226 8440 10232 8492
rect 10284 8480 10290 8492
rect 10502 8480 10508 8492
rect 10284 8452 10508 8480
rect 10284 8440 10290 8452
rect 10502 8440 10508 8452
rect 10560 8480 10566 8492
rect 10962 8480 10968 8492
rect 10560 8452 10968 8480
rect 10560 8440 10566 8452
rect 10962 8440 10968 8452
rect 11020 8440 11026 8492
rect 12250 8480 12256 8492
rect 12211 8452 12256 8480
rect 12250 8440 12256 8452
rect 12308 8440 12314 8492
rect 12894 8480 12900 8492
rect 12855 8452 12900 8480
rect 12894 8440 12900 8452
rect 12952 8440 12958 8492
rect 16850 8480 16856 8492
rect 16811 8452 16856 8480
rect 16850 8440 16856 8452
rect 16908 8440 16914 8492
rect 19076 8489 19104 8520
rect 19334 8508 19340 8520
rect 19392 8508 19398 8560
rect 20990 8548 20996 8560
rect 20562 8520 20996 8548
rect 20990 8508 20996 8520
rect 21048 8508 21054 8560
rect 19061 8483 19119 8489
rect 19061 8449 19073 8483
rect 19107 8449 19119 8483
rect 21100 8480 21128 8588
rect 21174 8576 21180 8628
rect 21232 8616 21238 8628
rect 22925 8619 22983 8625
rect 22925 8616 22937 8619
rect 21232 8588 22937 8616
rect 21232 8576 21238 8588
rect 22925 8585 22937 8588
rect 22971 8585 22983 8619
rect 22925 8579 22983 8585
rect 23566 8576 23572 8628
rect 23624 8616 23630 8628
rect 23753 8619 23811 8625
rect 23753 8616 23765 8619
rect 23624 8588 23765 8616
rect 23624 8576 23630 8588
rect 23753 8585 23765 8588
rect 23799 8585 23811 8619
rect 23753 8579 23811 8585
rect 24026 8576 24032 8628
rect 24084 8616 24090 8628
rect 24397 8619 24455 8625
rect 24397 8616 24409 8619
rect 24084 8588 24409 8616
rect 24084 8576 24090 8588
rect 24397 8585 24409 8588
rect 24443 8585 24455 8619
rect 25038 8616 25044 8628
rect 24999 8588 25044 8616
rect 24397 8579 24455 8585
rect 25038 8576 25044 8588
rect 25096 8576 25102 8628
rect 25961 8619 26019 8625
rect 25961 8585 25973 8619
rect 26007 8616 26019 8619
rect 26602 8616 26608 8628
rect 26007 8588 26608 8616
rect 26007 8585 26019 8588
rect 25961 8579 26019 8585
rect 26602 8576 26608 8588
rect 26660 8576 26666 8628
rect 29917 8619 29975 8625
rect 29917 8585 29929 8619
rect 29963 8616 29975 8619
rect 30374 8616 30380 8628
rect 29963 8588 30380 8616
rect 29963 8585 29975 8588
rect 29917 8579 29975 8585
rect 30374 8576 30380 8588
rect 30432 8576 30438 8628
rect 24118 8508 24124 8560
rect 24176 8548 24182 8560
rect 24176 8520 24992 8548
rect 24176 8508 24182 8520
rect 21100 8452 21220 8480
rect 19061 8443 19119 8449
rect 2884 8384 6592 8412
rect 2884 8353 2912 8384
rect 7098 8372 7104 8424
rect 7156 8412 7162 8424
rect 7558 8412 7564 8424
rect 7156 8384 7564 8412
rect 7156 8372 7162 8384
rect 7558 8372 7564 8384
rect 7616 8372 7622 8424
rect 8570 8412 8576 8424
rect 8531 8384 8576 8412
rect 8570 8372 8576 8384
rect 8628 8372 8634 8424
rect 8846 8412 8852 8424
rect 8807 8384 8852 8412
rect 8846 8372 8852 8384
rect 8904 8372 8910 8424
rect 8938 8372 8944 8424
rect 8996 8412 9002 8424
rect 10321 8415 10379 8421
rect 10321 8412 10333 8415
rect 8996 8384 10333 8412
rect 8996 8372 9002 8384
rect 10321 8381 10333 8384
rect 10367 8381 10379 8415
rect 10321 8375 10379 8381
rect 11057 8415 11115 8421
rect 11057 8381 11069 8415
rect 11103 8412 11115 8415
rect 12434 8412 12440 8424
rect 11103 8384 12440 8412
rect 11103 8381 11115 8384
rect 11057 8375 11115 8381
rect 12434 8372 12440 8384
rect 12492 8372 12498 8424
rect 16114 8412 16120 8424
rect 16075 8384 16120 8412
rect 16114 8372 16120 8384
rect 16172 8372 16178 8424
rect 19337 8415 19395 8421
rect 19337 8381 19349 8415
rect 19383 8412 19395 8415
rect 20070 8412 20076 8424
rect 19383 8384 20076 8412
rect 19383 8381 19395 8384
rect 19337 8375 19395 8381
rect 20070 8372 20076 8384
rect 20128 8372 20134 8424
rect 21085 8415 21143 8421
rect 21085 8381 21097 8415
rect 21131 8381 21143 8415
rect 21192 8412 21220 8452
rect 21358 8440 21364 8492
rect 21416 8480 21422 8492
rect 22833 8483 22891 8489
rect 22833 8480 22845 8483
rect 21416 8452 22845 8480
rect 21416 8440 21422 8452
rect 22833 8449 22845 8452
rect 22879 8449 22891 8483
rect 23658 8480 23664 8492
rect 23571 8452 23664 8480
rect 22833 8443 22891 8449
rect 23658 8440 23664 8452
rect 23716 8480 23722 8492
rect 24210 8480 24216 8492
rect 23716 8452 24216 8480
rect 23716 8440 23722 8452
rect 24210 8440 24216 8452
rect 24268 8440 24274 8492
rect 24964 8489 24992 8520
rect 24305 8483 24363 8489
rect 24305 8449 24317 8483
rect 24351 8449 24363 8483
rect 24305 8443 24363 8449
rect 24949 8483 25007 8489
rect 24949 8449 24961 8483
rect 24995 8449 25007 8483
rect 24949 8443 25007 8449
rect 25869 8483 25927 8489
rect 25869 8449 25881 8483
rect 25915 8480 25927 8483
rect 25958 8480 25964 8492
rect 25915 8452 25964 8480
rect 25915 8449 25927 8452
rect 25869 8443 25927 8449
rect 23382 8412 23388 8424
rect 21192 8384 23388 8412
rect 21085 8375 21143 8381
rect 2869 8347 2927 8353
rect 2869 8313 2881 8347
rect 2915 8313 2927 8347
rect 2869 8307 2927 8313
rect 5997 8347 6055 8353
rect 5997 8313 6009 8347
rect 6043 8344 6055 8347
rect 8478 8344 8484 8356
rect 6043 8316 8484 8344
rect 6043 8313 6055 8316
rect 5997 8307 6055 8313
rect 8478 8304 8484 8316
rect 8536 8304 8542 8356
rect 10134 8304 10140 8356
rect 10192 8344 10198 8356
rect 12894 8344 12900 8356
rect 10192 8316 12900 8344
rect 10192 8304 10198 8316
rect 12894 8304 12900 8316
rect 12952 8304 12958 8356
rect 18601 8347 18659 8353
rect 18601 8313 18613 8347
rect 18647 8344 18659 8347
rect 18647 8316 19196 8344
rect 18647 8313 18659 8316
rect 18601 8307 18659 8313
rect 3605 8279 3663 8285
rect 3605 8245 3617 8279
rect 3651 8276 3663 8279
rect 3970 8276 3976 8288
rect 3651 8248 3976 8276
rect 3651 8245 3663 8248
rect 3605 8239 3663 8245
rect 3970 8236 3976 8248
rect 4028 8236 4034 8288
rect 6822 8236 6828 8288
rect 6880 8276 6886 8288
rect 8018 8276 8024 8288
rect 6880 8248 8024 8276
rect 6880 8236 6886 8248
rect 8018 8236 8024 8248
rect 8076 8276 8082 8288
rect 8938 8276 8944 8288
rect 8076 8248 8944 8276
rect 8076 8236 8082 8248
rect 8938 8236 8944 8248
rect 8996 8236 9002 8288
rect 10042 8236 10048 8288
rect 10100 8276 10106 8288
rect 10594 8276 10600 8288
rect 10100 8248 10600 8276
rect 10100 8236 10106 8248
rect 10594 8236 10600 8248
rect 10652 8236 10658 8288
rect 14550 8236 14556 8288
rect 14608 8276 14614 8288
rect 15838 8276 15844 8288
rect 14608 8248 15844 8276
rect 14608 8236 14614 8248
rect 15838 8236 15844 8248
rect 15896 8236 15902 8288
rect 19168 8276 19196 8316
rect 20438 8304 20444 8356
rect 20496 8344 20502 8356
rect 21100 8344 21128 8375
rect 23382 8372 23388 8384
rect 23440 8372 23446 8424
rect 21266 8344 21272 8356
rect 20496 8316 21036 8344
rect 21100 8316 21272 8344
rect 20496 8304 20502 8316
rect 20346 8276 20352 8288
rect 19168 8248 20352 8276
rect 20346 8236 20352 8248
rect 20404 8236 20410 8288
rect 21008 8276 21036 8316
rect 21266 8304 21272 8316
rect 21324 8304 21330 8356
rect 24320 8344 24348 8443
rect 25958 8440 25964 8452
rect 26016 8440 26022 8492
rect 27338 8480 27344 8492
rect 27299 8452 27344 8480
rect 27338 8440 27344 8452
rect 27396 8440 27402 8492
rect 28442 8480 28448 8492
rect 28403 8452 28448 8480
rect 28442 8440 28448 8452
rect 28500 8440 28506 8492
rect 29270 8480 29276 8492
rect 29231 8452 29276 8480
rect 29270 8440 29276 8452
rect 29328 8440 29334 8492
rect 29454 8480 29460 8492
rect 29415 8452 29460 8480
rect 29454 8440 29460 8452
rect 29512 8440 29518 8492
rect 30377 8483 30435 8489
rect 30377 8449 30389 8483
rect 30423 8480 30435 8483
rect 38102 8480 38108 8492
rect 30423 8452 38108 8480
rect 30423 8449 30435 8452
rect 30377 8443 30435 8449
rect 38102 8440 38108 8452
rect 38160 8440 38166 8492
rect 21376 8316 24348 8344
rect 27157 8347 27215 8353
rect 21376 8276 21404 8316
rect 27157 8313 27169 8347
rect 27203 8344 27215 8347
rect 27706 8344 27712 8356
rect 27203 8316 27712 8344
rect 27203 8313 27215 8316
rect 27157 8307 27215 8313
rect 27706 8304 27712 8316
rect 27764 8304 27770 8356
rect 28626 8344 28632 8356
rect 28587 8316 28632 8344
rect 28626 8304 28632 8316
rect 28684 8304 28690 8356
rect 30466 8344 30472 8356
rect 30427 8316 30472 8344
rect 30466 8304 30472 8316
rect 30524 8304 30530 8356
rect 21008 8248 21404 8276
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 1946 8072 1952 8084
rect 1907 8044 1952 8072
rect 1946 8032 1952 8044
rect 2004 8032 2010 8084
rect 5445 8075 5503 8081
rect 5445 8041 5457 8075
rect 5491 8072 5503 8075
rect 5534 8072 5540 8084
rect 5491 8044 5540 8072
rect 5491 8041 5503 8044
rect 5445 8035 5503 8041
rect 5534 8032 5540 8044
rect 5592 8032 5598 8084
rect 7374 8032 7380 8084
rect 7432 8072 7438 8084
rect 14908 8075 14966 8081
rect 7432 8044 12434 8072
rect 7432 8032 7438 8044
rect 4062 8004 4068 8016
rect 4023 7976 4068 8004
rect 4062 7964 4068 7976
rect 4120 7964 4126 8016
rect 5902 7964 5908 8016
rect 5960 8004 5966 8016
rect 8481 8007 8539 8013
rect 5960 7976 6868 8004
rect 5960 7964 5966 7976
rect 3602 7936 3608 7948
rect 3252 7908 3608 7936
rect 1578 7828 1584 7880
rect 1636 7868 1642 7880
rect 3252 7877 3280 7908
rect 3602 7896 3608 7908
rect 3660 7936 3666 7948
rect 3660 7908 5120 7936
rect 3660 7896 3666 7908
rect 5092 7880 5120 7908
rect 6270 7896 6276 7948
rect 6328 7936 6334 7948
rect 6730 7936 6736 7948
rect 6328 7908 6736 7936
rect 6328 7896 6334 7908
rect 6730 7896 6736 7908
rect 6788 7896 6794 7948
rect 6840 7936 6868 7976
rect 8481 7973 8493 8007
rect 8527 8004 8539 8007
rect 8662 8004 8668 8016
rect 8527 7976 8668 8004
rect 8527 7973 8539 7976
rect 8481 7967 8539 7973
rect 8662 7964 8668 7976
rect 8720 7964 8726 8016
rect 10594 7964 10600 8016
rect 10652 8004 10658 8016
rect 10873 8007 10931 8013
rect 10873 8004 10885 8007
rect 10652 7976 10885 8004
rect 10652 7964 10658 7976
rect 10873 7973 10885 7976
rect 10919 7973 10931 8007
rect 12406 8004 12434 8044
rect 14908 8041 14920 8075
rect 14954 8072 14966 8075
rect 16758 8072 16764 8084
rect 14954 8044 16764 8072
rect 14954 8041 14966 8044
rect 14908 8035 14966 8041
rect 16758 8032 16764 8044
rect 16816 8032 16822 8084
rect 18877 8075 18935 8081
rect 18877 8041 18889 8075
rect 18923 8072 18935 8075
rect 19058 8072 19064 8084
rect 18923 8044 19064 8072
rect 18923 8041 18935 8044
rect 18877 8035 18935 8041
rect 19058 8032 19064 8044
rect 19116 8032 19122 8084
rect 20990 8032 20996 8084
rect 21048 8072 21054 8084
rect 23293 8075 23351 8081
rect 23293 8072 23305 8075
rect 21048 8044 23305 8072
rect 21048 8032 21054 8044
rect 23293 8041 23305 8044
rect 23339 8041 23351 8075
rect 23293 8035 23351 8041
rect 23750 8032 23756 8084
rect 23808 8072 23814 8084
rect 24673 8075 24731 8081
rect 23808 8044 24624 8072
rect 23808 8032 23814 8044
rect 14550 8004 14556 8016
rect 12406 7976 14556 8004
rect 10873 7967 10931 7973
rect 14550 7964 14556 7976
rect 14608 7964 14614 8016
rect 16393 8007 16451 8013
rect 16393 7973 16405 8007
rect 16439 8004 16451 8007
rect 18690 8004 18696 8016
rect 16439 7976 17264 8004
rect 16439 7973 16451 7976
rect 16393 7967 16451 7973
rect 6840 7908 8248 7936
rect 2133 7871 2191 7877
rect 2133 7868 2145 7871
rect 1636 7840 2145 7868
rect 1636 7828 1642 7840
rect 2133 7837 2145 7840
rect 2179 7837 2191 7871
rect 2133 7831 2191 7837
rect 2593 7871 2651 7877
rect 2593 7837 2605 7871
rect 2639 7837 2651 7871
rect 2593 7831 2651 7837
rect 3237 7871 3295 7877
rect 3237 7837 3249 7871
rect 3283 7837 3295 7871
rect 3970 7868 3976 7880
rect 3931 7840 3976 7868
rect 3237 7831 3295 7837
rect 2608 7800 2636 7831
rect 3970 7828 3976 7840
rect 4028 7828 4034 7880
rect 4709 7871 4767 7877
rect 4709 7837 4721 7871
rect 4755 7837 4767 7871
rect 4709 7831 4767 7837
rect 4614 7800 4620 7812
rect 2608 7772 4620 7800
rect 4614 7760 4620 7772
rect 4672 7800 4678 7812
rect 4724 7800 4752 7831
rect 5074 7828 5080 7880
rect 5132 7868 5138 7880
rect 5353 7871 5411 7877
rect 5353 7868 5365 7871
rect 5132 7840 5365 7868
rect 5132 7828 5138 7840
rect 5353 7837 5365 7840
rect 5399 7837 5411 7871
rect 5353 7831 5411 7837
rect 5997 7871 6055 7877
rect 5997 7837 6009 7871
rect 6043 7868 6055 7871
rect 6546 7868 6552 7880
rect 6043 7840 6552 7868
rect 6043 7837 6055 7840
rect 5997 7831 6055 7837
rect 6546 7828 6552 7840
rect 6604 7828 6610 7880
rect 8220 7868 8248 7908
rect 8570 7896 8576 7948
rect 8628 7936 8634 7948
rect 9125 7939 9183 7945
rect 9125 7936 9137 7939
rect 8628 7908 9137 7936
rect 8628 7896 8634 7908
rect 9125 7905 9137 7908
rect 9171 7905 9183 7939
rect 9125 7899 9183 7905
rect 9401 7939 9459 7945
rect 9401 7905 9413 7939
rect 9447 7936 9459 7939
rect 14090 7936 14096 7948
rect 9447 7908 14096 7936
rect 9447 7905 9459 7908
rect 9401 7899 9459 7905
rect 14090 7896 14096 7908
rect 14148 7896 14154 7948
rect 14182 7896 14188 7948
rect 14240 7936 14246 7948
rect 14645 7939 14703 7945
rect 14645 7936 14657 7939
rect 14240 7908 14657 7936
rect 14240 7896 14246 7908
rect 14645 7905 14657 7908
rect 14691 7936 14703 7939
rect 16114 7936 16120 7948
rect 14691 7908 16120 7936
rect 14691 7905 14703 7908
rect 14645 7899 14703 7905
rect 16114 7896 16120 7908
rect 16172 7896 16178 7948
rect 16850 7896 16856 7948
rect 16908 7936 16914 7948
rect 17129 7939 17187 7945
rect 17129 7936 17141 7939
rect 16908 7908 17141 7936
rect 16908 7896 16914 7908
rect 17129 7905 17141 7908
rect 17175 7905 17187 7939
rect 17236 7936 17264 7976
rect 18432 7976 18696 8004
rect 17405 7939 17463 7945
rect 17405 7936 17417 7939
rect 17236 7908 17417 7936
rect 17129 7899 17187 7905
rect 17405 7905 17417 7908
rect 17451 7936 17463 7939
rect 18432 7936 18460 7976
rect 18690 7964 18696 7976
rect 18748 7964 18754 8016
rect 21542 7964 21548 8016
rect 21600 8004 21606 8016
rect 21729 8007 21787 8013
rect 21729 8004 21741 8007
rect 21600 7976 21741 8004
rect 21600 7964 21606 7976
rect 21729 7973 21741 7976
rect 21775 7973 21787 8007
rect 21729 7967 21787 7973
rect 21818 7964 21824 8016
rect 21876 8004 21882 8016
rect 24596 8004 24624 8044
rect 24673 8041 24685 8075
rect 24719 8072 24731 8075
rect 24762 8072 24768 8084
rect 24719 8044 24768 8072
rect 24719 8041 24731 8044
rect 24673 8035 24731 8041
rect 24762 8032 24768 8044
rect 24820 8032 24826 8084
rect 25958 8032 25964 8084
rect 26016 8072 26022 8084
rect 26016 8044 35894 8072
rect 26016 8032 26022 8044
rect 25317 8007 25375 8013
rect 25317 8004 25329 8007
rect 21876 7976 24072 8004
rect 24596 7976 25329 8004
rect 21876 7964 21882 7976
rect 23937 7939 23995 7945
rect 23937 7936 23949 7939
rect 17451 7908 18460 7936
rect 18524 7908 23949 7936
rect 17451 7905 17463 7908
rect 17405 7899 17463 7905
rect 8754 7868 8760 7880
rect 8220 7840 8760 7868
rect 8754 7828 8760 7840
rect 8812 7828 8818 7880
rect 10962 7828 10968 7880
rect 11020 7868 11026 7880
rect 11020 7840 12434 7868
rect 11020 7828 11026 7840
rect 4672 7772 4752 7800
rect 4672 7760 4678 7772
rect 2685 7735 2743 7741
rect 2685 7701 2697 7735
rect 2731 7732 2743 7735
rect 3142 7732 3148 7744
rect 2731 7704 3148 7732
rect 2731 7701 2743 7704
rect 2685 7695 2743 7701
rect 3142 7692 3148 7704
rect 3200 7692 3206 7744
rect 3329 7735 3387 7741
rect 3329 7701 3341 7735
rect 3375 7732 3387 7735
rect 3418 7732 3424 7744
rect 3375 7704 3424 7732
rect 3375 7701 3387 7704
rect 3329 7695 3387 7701
rect 3418 7692 3424 7704
rect 3476 7692 3482 7744
rect 4724 7732 4752 7772
rect 4801 7803 4859 7809
rect 4801 7769 4813 7803
rect 4847 7800 4859 7803
rect 6914 7800 6920 7812
rect 4847 7772 6920 7800
rect 4847 7769 4859 7772
rect 4801 7763 4859 7769
rect 6914 7760 6920 7772
rect 6972 7760 6978 7812
rect 7009 7803 7067 7809
rect 7009 7769 7021 7803
rect 7055 7800 7067 7803
rect 7098 7800 7104 7812
rect 7055 7772 7104 7800
rect 7055 7769 7067 7772
rect 7009 7763 7067 7769
rect 7098 7760 7104 7772
rect 7156 7760 7162 7812
rect 7466 7760 7472 7812
rect 7524 7760 7530 7812
rect 8294 7760 8300 7812
rect 8352 7800 8358 7812
rect 11977 7803 12035 7809
rect 8352 7772 9890 7800
rect 8352 7760 8358 7772
rect 11977 7769 11989 7803
rect 12023 7769 12035 7803
rect 12406 7800 12434 7840
rect 12894 7828 12900 7880
rect 12952 7868 12958 7880
rect 13354 7868 13360 7880
rect 12952 7840 13360 7868
rect 12952 7828 12958 7840
rect 13354 7828 13360 7840
rect 13412 7868 13418 7880
rect 13541 7871 13599 7877
rect 13541 7868 13553 7871
rect 13412 7840 13553 7868
rect 13412 7828 13418 7840
rect 13541 7837 13553 7840
rect 13587 7837 13599 7871
rect 18524 7854 18552 7908
rect 23937 7905 23949 7908
rect 23983 7905 23995 7939
rect 23937 7899 23995 7905
rect 19978 7868 19984 7880
rect 19939 7840 19984 7868
rect 13541 7831 13599 7837
rect 19978 7828 19984 7840
rect 20036 7828 20042 7880
rect 22370 7828 22376 7880
rect 22428 7868 22434 7880
rect 23201 7871 23259 7877
rect 23201 7868 23213 7871
rect 22428 7840 23213 7868
rect 22428 7828 22434 7840
rect 23201 7837 23213 7840
rect 23247 7868 23259 7871
rect 23658 7868 23664 7880
rect 23247 7840 23664 7868
rect 23247 7837 23259 7840
rect 23201 7831 23259 7837
rect 23658 7828 23664 7840
rect 23716 7828 23722 7880
rect 23845 7871 23903 7877
rect 23845 7837 23857 7871
rect 23891 7868 23903 7871
rect 24044 7868 24072 7976
rect 25317 7973 25329 7976
rect 25363 7973 25375 8007
rect 25317 7967 25375 7973
rect 28994 7964 29000 8016
rect 29052 8004 29058 8016
rect 31662 8004 31668 8016
rect 29052 7976 31668 8004
rect 29052 7964 29058 7976
rect 31662 7964 31668 7976
rect 31720 7964 31726 8016
rect 24210 7896 24216 7948
rect 24268 7936 24274 7948
rect 24762 7936 24768 7948
rect 24268 7908 24768 7936
rect 24268 7896 24274 7908
rect 24762 7896 24768 7908
rect 24820 7896 24826 7948
rect 27246 7936 27252 7948
rect 24872 7908 27108 7936
rect 27207 7908 27252 7936
rect 24486 7868 24492 7880
rect 23891 7840 24492 7868
rect 23891 7837 23903 7840
rect 23845 7831 23903 7837
rect 24486 7828 24492 7840
rect 24544 7828 24550 7880
rect 24581 7871 24639 7877
rect 24581 7837 24593 7871
rect 24627 7837 24639 7871
rect 24581 7831 24639 7837
rect 16666 7800 16672 7812
rect 12406 7772 13400 7800
rect 16146 7772 16672 7800
rect 11977 7763 12035 7769
rect 5350 7732 5356 7744
rect 4724 7704 5356 7732
rect 5350 7692 5356 7704
rect 5408 7692 5414 7744
rect 6086 7732 6092 7744
rect 6047 7704 6092 7732
rect 6086 7692 6092 7704
rect 6144 7692 6150 7744
rect 7650 7692 7656 7744
rect 7708 7732 7714 7744
rect 11992 7732 12020 7763
rect 7708 7704 12020 7732
rect 13372 7732 13400 7772
rect 16666 7760 16672 7772
rect 16724 7760 16730 7812
rect 20257 7803 20315 7809
rect 20257 7769 20269 7803
rect 20303 7769 20315 7803
rect 22002 7800 22008 7812
rect 21482 7772 22008 7800
rect 20257 7763 20315 7769
rect 16298 7732 16304 7744
rect 13372 7704 16304 7732
rect 7708 7692 7714 7704
rect 16298 7692 16304 7704
rect 16356 7692 16362 7744
rect 20272 7732 20300 7763
rect 22002 7760 22008 7772
rect 22060 7760 22066 7812
rect 22922 7760 22928 7812
rect 22980 7800 22986 7812
rect 24596 7800 24624 7831
rect 22980 7772 24624 7800
rect 22980 7760 22986 7772
rect 21266 7732 21272 7744
rect 20272 7704 21272 7732
rect 21266 7692 21272 7704
rect 21324 7692 21330 7744
rect 21542 7692 21548 7744
rect 21600 7732 21606 7744
rect 24872 7732 24900 7908
rect 24946 7828 24952 7880
rect 25004 7868 25010 7880
rect 25225 7871 25283 7877
rect 25225 7868 25237 7871
rect 25004 7840 25237 7868
rect 25004 7828 25010 7840
rect 25225 7837 25237 7840
rect 25271 7837 25283 7871
rect 27080 7868 27108 7908
rect 27246 7896 27252 7908
rect 27304 7896 27310 7948
rect 35866 7936 35894 8044
rect 37737 7939 37795 7945
rect 37737 7936 37749 7939
rect 35866 7908 37749 7936
rect 37737 7905 37749 7908
rect 37783 7905 37795 7939
rect 37737 7899 37795 7905
rect 27709 7871 27767 7877
rect 27709 7868 27721 7871
rect 27080 7840 27721 7868
rect 25225 7831 25283 7837
rect 27709 7837 27721 7840
rect 27755 7837 27767 7871
rect 37458 7868 37464 7880
rect 37419 7840 37464 7868
rect 27709 7831 27767 7837
rect 21600 7704 24900 7732
rect 25240 7732 25268 7831
rect 37458 7828 37464 7840
rect 37516 7828 37522 7880
rect 26234 7800 26240 7812
rect 26195 7772 26240 7800
rect 26234 7760 26240 7772
rect 26292 7760 26298 7812
rect 26329 7803 26387 7809
rect 26329 7769 26341 7803
rect 26375 7800 26387 7803
rect 27801 7803 27859 7809
rect 27801 7800 27813 7803
rect 26375 7772 27813 7800
rect 26375 7769 26387 7772
rect 26329 7763 26387 7769
rect 27801 7769 27813 7772
rect 27847 7769 27859 7803
rect 27801 7763 27859 7769
rect 27430 7732 27436 7744
rect 25240 7704 27436 7732
rect 21600 7692 21606 7704
rect 27430 7692 27436 7704
rect 27488 7692 27494 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 2498 7488 2504 7540
rect 2556 7528 2562 7540
rect 2593 7531 2651 7537
rect 2593 7528 2605 7531
rect 2556 7500 2605 7528
rect 2556 7488 2562 7500
rect 2593 7497 2605 7500
rect 2639 7528 2651 7531
rect 2682 7528 2688 7540
rect 2639 7500 2688 7528
rect 2639 7497 2651 7500
rect 2593 7491 2651 7497
rect 2682 7488 2688 7500
rect 2740 7488 2746 7540
rect 8018 7528 8024 7540
rect 6656 7500 8024 7528
rect 4706 7460 4712 7472
rect 3252 7432 4712 7460
rect 3252 7401 3280 7432
rect 4706 7420 4712 7432
rect 4764 7420 4770 7472
rect 5350 7460 5356 7472
rect 5000 7432 5356 7460
rect 3237 7395 3295 7401
rect 3237 7361 3249 7395
rect 3283 7361 3295 7395
rect 3237 7355 3295 7361
rect 3329 7395 3387 7401
rect 3329 7361 3341 7395
rect 3375 7392 3387 7395
rect 3694 7392 3700 7404
rect 3375 7364 3700 7392
rect 3375 7361 3387 7364
rect 3329 7355 3387 7361
rect 3694 7352 3700 7364
rect 3752 7352 3758 7404
rect 4065 7395 4123 7401
rect 4065 7361 4077 7395
rect 4111 7361 4123 7395
rect 4065 7355 4123 7361
rect 4525 7395 4583 7401
rect 4525 7361 4537 7395
rect 4571 7392 4583 7395
rect 5000 7392 5028 7432
rect 5350 7420 5356 7432
rect 5408 7460 5414 7472
rect 5408 7432 5764 7460
rect 5408 7420 5414 7432
rect 4571 7364 5028 7392
rect 4571 7361 4583 7364
rect 4525 7355 4583 7361
rect 1946 7324 1952 7336
rect 1907 7296 1952 7324
rect 1946 7284 1952 7296
rect 2004 7284 2010 7336
rect 2130 7324 2136 7336
rect 2091 7296 2136 7324
rect 2130 7284 2136 7296
rect 2188 7284 2194 7336
rect 2222 7284 2228 7336
rect 2280 7324 2286 7336
rect 2590 7324 2596 7336
rect 2280 7296 2596 7324
rect 2280 7284 2286 7296
rect 2590 7284 2596 7296
rect 2648 7284 2654 7336
rect 4080 7324 4108 7355
rect 5074 7352 5080 7404
rect 5132 7392 5138 7404
rect 5169 7395 5227 7401
rect 5169 7392 5181 7395
rect 5132 7364 5181 7392
rect 5132 7352 5138 7364
rect 5169 7361 5181 7364
rect 5215 7361 5227 7395
rect 5736 7392 5764 7432
rect 5813 7395 5871 7401
rect 5813 7392 5825 7395
rect 5736 7364 5825 7392
rect 5169 7355 5227 7361
rect 5813 7361 5825 7364
rect 5859 7361 5871 7395
rect 5813 7355 5871 7361
rect 6656 7324 6684 7500
rect 8018 7488 8024 7500
rect 8076 7488 8082 7540
rect 8754 7488 8760 7540
rect 8812 7528 8818 7540
rect 8812 7500 12434 7528
rect 8812 7488 8818 7500
rect 7834 7420 7840 7472
rect 7892 7420 7898 7472
rect 12406 7460 12434 7500
rect 13170 7488 13176 7540
rect 13228 7528 13234 7540
rect 13633 7531 13691 7537
rect 13633 7528 13645 7531
rect 13228 7500 13645 7528
rect 13228 7488 13234 7500
rect 13633 7497 13645 7500
rect 13679 7528 13691 7531
rect 14274 7528 14280 7540
rect 13679 7500 14280 7528
rect 13679 7497 13691 7500
rect 13633 7491 13691 7497
rect 14274 7488 14280 7500
rect 14332 7488 14338 7540
rect 15838 7488 15844 7540
rect 15896 7528 15902 7540
rect 15933 7531 15991 7537
rect 15933 7528 15945 7531
rect 15896 7500 15945 7528
rect 15896 7488 15902 7500
rect 15933 7497 15945 7500
rect 15979 7497 15991 7531
rect 15933 7491 15991 7497
rect 17512 7500 19748 7528
rect 8937 7432 10074 7460
rect 12406 7432 12650 7460
rect 6730 7352 6736 7404
rect 6788 7392 6794 7404
rect 7101 7395 7159 7401
rect 7101 7392 7113 7395
rect 6788 7364 7113 7392
rect 6788 7352 6794 7364
rect 7101 7361 7113 7364
rect 7147 7361 7159 7395
rect 7101 7355 7159 7361
rect 7374 7324 7380 7336
rect 4080 7296 6684 7324
rect 7335 7296 7380 7324
rect 7374 7284 7380 7296
rect 7432 7284 7438 7336
rect 7926 7284 7932 7336
rect 7984 7324 7990 7336
rect 8849 7327 8907 7333
rect 8849 7324 8861 7327
rect 7984 7296 8861 7324
rect 7984 7284 7990 7296
rect 8849 7293 8861 7296
rect 8895 7293 8907 7327
rect 8849 7287 8907 7293
rect 4522 7216 4528 7268
rect 4580 7256 4586 7268
rect 4617 7259 4675 7265
rect 4617 7256 4629 7259
rect 4580 7228 4629 7256
rect 4580 7216 4586 7228
rect 4617 7225 4629 7228
rect 4663 7225 4675 7259
rect 4617 7219 4675 7225
rect 5074 7216 5080 7268
rect 5132 7256 5138 7268
rect 5261 7259 5319 7265
rect 5261 7256 5273 7259
rect 5132 7228 5273 7256
rect 5132 7216 5138 7228
rect 5261 7225 5273 7228
rect 5307 7225 5319 7259
rect 5261 7219 5319 7225
rect 5905 7259 5963 7265
rect 5905 7225 5917 7259
rect 5951 7256 5963 7259
rect 5951 7228 7236 7256
rect 5951 7225 5963 7228
rect 5905 7219 5963 7225
rect 2774 7148 2780 7200
rect 2832 7188 2838 7200
rect 3881 7191 3939 7197
rect 3881 7188 3893 7191
rect 2832 7160 3893 7188
rect 2832 7148 2838 7160
rect 3881 7157 3893 7160
rect 3927 7157 3939 7191
rect 3881 7151 3939 7157
rect 5442 7148 5448 7200
rect 5500 7188 5506 7200
rect 7098 7188 7104 7200
rect 5500 7160 7104 7188
rect 5500 7148 5506 7160
rect 7098 7148 7104 7160
rect 7156 7148 7162 7200
rect 7208 7188 7236 7228
rect 8937 7188 8965 7432
rect 15194 7420 15200 7472
rect 15252 7420 15258 7472
rect 14182 7392 14188 7404
rect 14143 7364 14188 7392
rect 14182 7352 14188 7364
rect 14240 7352 14246 7404
rect 16482 7352 16488 7404
rect 16540 7392 16546 7404
rect 16853 7395 16911 7401
rect 16853 7392 16865 7395
rect 16540 7364 16865 7392
rect 16540 7352 16546 7364
rect 16853 7361 16865 7364
rect 16899 7361 16911 7395
rect 16853 7355 16911 7361
rect 17218 7352 17224 7404
rect 17276 7392 17282 7404
rect 17512 7401 17540 7500
rect 17770 7460 17776 7472
rect 17731 7432 17776 7460
rect 17770 7420 17776 7432
rect 17828 7420 17834 7472
rect 19720 7460 19748 7500
rect 19978 7488 19984 7540
rect 20036 7528 20042 7540
rect 20036 7500 22094 7528
rect 20036 7488 20042 7500
rect 19996 7460 20024 7488
rect 21358 7460 21364 7472
rect 19720 7432 20024 7460
rect 21206 7432 21364 7460
rect 19720 7404 19748 7432
rect 21358 7420 21364 7432
rect 21416 7420 21422 7472
rect 22066 7460 22094 7500
rect 23382 7488 23388 7540
rect 23440 7528 23446 7540
rect 25133 7531 25191 7537
rect 25133 7528 25145 7531
rect 23440 7500 25145 7528
rect 23440 7488 23446 7500
rect 25133 7497 25145 7500
rect 25179 7497 25191 7531
rect 25774 7528 25780 7540
rect 25735 7500 25780 7528
rect 25133 7491 25191 7497
rect 25774 7488 25780 7500
rect 25832 7488 25838 7540
rect 26234 7488 26240 7540
rect 26292 7528 26298 7540
rect 27801 7531 27859 7537
rect 27801 7528 27813 7531
rect 26292 7500 27813 7528
rect 26292 7488 26298 7500
rect 27801 7497 27813 7500
rect 27847 7497 27859 7531
rect 27801 7491 27859 7497
rect 34054 7488 34060 7540
rect 34112 7528 34118 7540
rect 38105 7531 38163 7537
rect 38105 7528 38117 7531
rect 34112 7500 38117 7528
rect 34112 7488 34118 7500
rect 38105 7497 38117 7500
rect 38151 7497 38163 7531
rect 38105 7491 38163 7497
rect 22741 7463 22799 7469
rect 22741 7460 22753 7463
rect 22066 7432 22753 7460
rect 22741 7429 22753 7432
rect 22787 7429 22799 7463
rect 22741 7423 22799 7429
rect 23106 7420 23112 7472
rect 23164 7460 23170 7472
rect 23937 7463 23995 7469
rect 23937 7460 23949 7463
rect 23164 7432 23949 7460
rect 23164 7420 23170 7432
rect 23937 7429 23949 7432
rect 23983 7429 23995 7463
rect 23937 7423 23995 7429
rect 24029 7463 24087 7469
rect 24029 7429 24041 7463
rect 24075 7460 24087 7463
rect 26421 7463 26479 7469
rect 26421 7460 26433 7463
rect 24075 7432 26433 7460
rect 24075 7429 24087 7432
rect 24029 7423 24087 7429
rect 26421 7429 26433 7432
rect 26467 7429 26479 7463
rect 26421 7423 26479 7429
rect 17497 7395 17555 7401
rect 17497 7392 17509 7395
rect 17276 7364 17509 7392
rect 17276 7352 17282 7364
rect 17497 7361 17509 7364
rect 17543 7361 17555 7395
rect 17497 7355 17555 7361
rect 18874 7352 18880 7404
rect 18932 7352 18938 7404
rect 19702 7392 19708 7404
rect 19615 7364 19708 7392
rect 19702 7352 19708 7364
rect 19760 7352 19766 7404
rect 22005 7395 22063 7401
rect 22005 7361 22017 7395
rect 22051 7361 22063 7395
rect 22005 7355 22063 7361
rect 9306 7324 9312 7336
rect 9267 7296 9312 7324
rect 9306 7284 9312 7296
rect 9364 7284 9370 7336
rect 9585 7327 9643 7333
rect 9585 7293 9597 7327
rect 9631 7324 9643 7327
rect 9674 7324 9680 7336
rect 9631 7296 9680 7324
rect 9631 7293 9643 7296
rect 9585 7287 9643 7293
rect 9674 7284 9680 7296
rect 9732 7284 9738 7336
rect 11606 7284 11612 7336
rect 11664 7324 11670 7336
rect 11885 7327 11943 7333
rect 11885 7324 11897 7327
rect 11664 7296 11897 7324
rect 11664 7284 11670 7296
rect 11885 7293 11897 7296
rect 11931 7293 11943 7327
rect 12158 7324 12164 7336
rect 12119 7296 12164 7324
rect 11885 7287 11943 7293
rect 7208 7160 8965 7188
rect 10962 7148 10968 7200
rect 11020 7188 11026 7200
rect 11057 7191 11115 7197
rect 11057 7188 11069 7191
rect 11020 7160 11069 7188
rect 11020 7148 11026 7160
rect 11057 7157 11069 7160
rect 11103 7157 11115 7191
rect 11900 7188 11928 7287
rect 12158 7284 12164 7296
rect 12216 7284 12222 7336
rect 14461 7327 14519 7333
rect 14461 7293 14473 7327
rect 14507 7324 14519 7327
rect 16206 7324 16212 7336
rect 14507 7296 16212 7324
rect 14507 7293 14519 7296
rect 14461 7287 14519 7293
rect 16206 7284 16212 7296
rect 16264 7284 16270 7336
rect 17770 7284 17776 7336
rect 17828 7324 17834 7336
rect 19610 7324 19616 7336
rect 17828 7296 19616 7324
rect 17828 7284 17834 7296
rect 19610 7284 19616 7296
rect 19668 7284 19674 7336
rect 19981 7327 20039 7333
rect 19981 7293 19993 7327
rect 20027 7324 20039 7327
rect 20346 7324 20352 7336
rect 20027 7296 20352 7324
rect 20027 7293 20039 7296
rect 19981 7287 20039 7293
rect 20346 7284 20352 7296
rect 20404 7284 20410 7336
rect 20622 7284 20628 7336
rect 20680 7324 20686 7336
rect 22020 7324 22048 7355
rect 24762 7352 24768 7404
rect 24820 7392 24826 7404
rect 25041 7395 25099 7401
rect 25041 7392 25053 7395
rect 24820 7364 25053 7392
rect 24820 7352 24826 7364
rect 25041 7361 25053 7364
rect 25087 7392 25099 7395
rect 25685 7395 25743 7401
rect 25685 7392 25697 7395
rect 25087 7364 25697 7392
rect 25087 7361 25099 7364
rect 25041 7355 25099 7361
rect 25685 7361 25697 7364
rect 25731 7361 25743 7395
rect 25685 7355 25743 7361
rect 26234 7352 26240 7404
rect 26292 7392 26298 7404
rect 26329 7395 26387 7401
rect 26329 7392 26341 7395
rect 26292 7364 26341 7392
rect 26292 7352 26298 7364
rect 26329 7361 26341 7364
rect 26375 7361 26387 7395
rect 26329 7355 26387 7361
rect 26510 7352 26516 7404
rect 26568 7392 26574 7404
rect 27157 7395 27215 7401
rect 27157 7392 27169 7395
rect 26568 7364 27169 7392
rect 26568 7352 26574 7364
rect 27157 7361 27169 7364
rect 27203 7392 27215 7395
rect 27890 7392 27896 7404
rect 27203 7364 27896 7392
rect 27203 7361 27215 7364
rect 27157 7355 27215 7361
rect 27890 7352 27896 7364
rect 27948 7352 27954 7404
rect 34241 7395 34299 7401
rect 34241 7392 34253 7395
rect 31726 7364 34253 7392
rect 24210 7324 24216 7336
rect 20680 7296 22048 7324
rect 24171 7296 24216 7324
rect 20680 7284 20686 7296
rect 24210 7284 24216 7296
rect 24268 7284 24274 7336
rect 24946 7324 24952 7336
rect 24412 7296 24952 7324
rect 14182 7256 14188 7268
rect 13556 7228 14188 7256
rect 13556 7188 13584 7228
rect 14182 7216 14188 7228
rect 14240 7216 14246 7268
rect 17494 7256 17500 7268
rect 16868 7228 17500 7256
rect 11900 7160 13584 7188
rect 11057 7151 11115 7157
rect 14090 7148 14096 7200
rect 14148 7188 14154 7200
rect 16868 7188 16896 7228
rect 17494 7216 17500 7228
rect 17552 7216 17558 7268
rect 20990 7216 20996 7268
rect 21048 7256 21054 7268
rect 21048 7228 21864 7256
rect 21048 7216 21054 7228
rect 14148 7160 16896 7188
rect 16945 7191 17003 7197
rect 14148 7148 14154 7160
rect 16945 7157 16957 7191
rect 16991 7188 17003 7191
rect 18138 7188 18144 7200
rect 16991 7160 18144 7188
rect 16991 7157 17003 7160
rect 16945 7151 17003 7157
rect 18138 7148 18144 7160
rect 18196 7148 18202 7200
rect 19245 7191 19303 7197
rect 19245 7157 19257 7191
rect 19291 7188 19303 7191
rect 20162 7188 20168 7200
rect 19291 7160 20168 7188
rect 19291 7157 19303 7160
rect 19245 7151 19303 7157
rect 20162 7148 20168 7160
rect 20220 7148 20226 7200
rect 21082 7148 21088 7200
rect 21140 7188 21146 7200
rect 21453 7191 21511 7197
rect 21453 7188 21465 7191
rect 21140 7160 21465 7188
rect 21140 7148 21146 7160
rect 21453 7157 21465 7160
rect 21499 7157 21511 7191
rect 21836 7188 21864 7228
rect 21910 7216 21916 7268
rect 21968 7256 21974 7268
rect 24412 7256 24440 7296
rect 24946 7284 24952 7296
rect 25004 7284 25010 7336
rect 25774 7284 25780 7336
rect 25832 7324 25838 7336
rect 31726 7324 31754 7364
rect 34241 7361 34253 7364
rect 34287 7361 34299 7395
rect 38286 7392 38292 7404
rect 38247 7364 38292 7392
rect 34241 7355 34299 7361
rect 38286 7352 38292 7364
rect 38344 7352 38350 7404
rect 25832 7296 31754 7324
rect 25832 7284 25838 7296
rect 21968 7228 24440 7256
rect 21968 7216 21974 7228
rect 24486 7216 24492 7268
rect 24544 7256 24550 7268
rect 29546 7256 29552 7268
rect 24544 7228 29552 7256
rect 24544 7216 24550 7228
rect 29546 7216 29552 7228
rect 29604 7216 29610 7268
rect 26234 7188 26240 7200
rect 21836 7160 26240 7188
rect 21453 7151 21511 7157
rect 26234 7148 26240 7160
rect 26292 7148 26298 7200
rect 26326 7148 26332 7200
rect 26384 7188 26390 7200
rect 27249 7191 27307 7197
rect 27249 7188 27261 7191
rect 26384 7160 27261 7188
rect 26384 7148 26390 7160
rect 27249 7157 27261 7160
rect 27295 7157 27307 7191
rect 27249 7151 27307 7157
rect 34333 7191 34391 7197
rect 34333 7157 34345 7191
rect 34379 7188 34391 7191
rect 35802 7188 35808 7200
rect 34379 7160 35808 7188
rect 34379 7157 34391 7160
rect 34333 7151 34391 7157
rect 35802 7148 35808 7160
rect 35860 7148 35866 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 2682 6984 2688 6996
rect 2643 6956 2688 6984
rect 2682 6944 2688 6956
rect 2740 6944 2746 6996
rect 7466 6984 7472 6996
rect 5552 6956 7472 6984
rect 1946 6876 1952 6928
rect 2004 6916 2010 6928
rect 5442 6916 5448 6928
rect 2004 6888 5448 6916
rect 2004 6876 2010 6888
rect 5442 6876 5448 6888
rect 5500 6876 5506 6928
rect 2409 6851 2467 6857
rect 2409 6817 2421 6851
rect 2455 6848 2467 6851
rect 2866 6848 2872 6860
rect 2455 6820 2872 6848
rect 2455 6817 2467 6820
rect 2409 6811 2467 6817
rect 2866 6808 2872 6820
rect 2924 6808 2930 6860
rect 4985 6851 5043 6857
rect 4985 6817 4997 6851
rect 5031 6848 5043 6851
rect 5552 6848 5580 6956
rect 7466 6944 7472 6956
rect 7524 6944 7530 6996
rect 7558 6944 7564 6996
rect 7616 6984 7622 6996
rect 10962 6984 10968 6996
rect 7616 6956 10968 6984
rect 7616 6944 7622 6956
rect 10962 6944 10968 6956
rect 11020 6944 11026 6996
rect 11964 6987 12022 6993
rect 11964 6953 11976 6987
rect 12010 6984 12022 6987
rect 12066 6984 12072 6996
rect 12010 6956 12072 6984
rect 12010 6953 12022 6956
rect 11964 6947 12022 6953
rect 12066 6944 12072 6956
rect 12124 6944 12130 6996
rect 12158 6944 12164 6996
rect 12216 6984 12222 6996
rect 17116 6987 17174 6993
rect 17116 6984 17128 6987
rect 12216 6956 17128 6984
rect 12216 6944 12222 6956
rect 17116 6953 17128 6956
rect 17162 6984 17174 6987
rect 17162 6956 18184 6984
rect 17162 6953 17174 6956
rect 17116 6947 17174 6953
rect 6178 6876 6184 6928
rect 6236 6916 6242 6928
rect 6546 6916 6552 6928
rect 6236 6888 6552 6916
rect 6236 6876 6242 6888
rect 6546 6876 6552 6888
rect 6604 6876 6610 6928
rect 6656 6888 6960 6916
rect 5031 6820 5580 6848
rect 5629 6851 5687 6857
rect 5031 6817 5043 6820
rect 4985 6811 5043 6817
rect 5629 6817 5641 6851
rect 5675 6848 5687 6851
rect 6656 6848 6684 6888
rect 5675 6820 6684 6848
rect 5675 6817 5687 6820
rect 5629 6811 5687 6817
rect 6730 6808 6736 6860
rect 6788 6848 6794 6860
rect 6825 6851 6883 6857
rect 6825 6848 6837 6851
rect 6788 6820 6837 6848
rect 6788 6808 6794 6820
rect 6825 6817 6837 6820
rect 6871 6817 6883 6851
rect 6932 6848 6960 6888
rect 13262 6876 13268 6928
rect 13320 6916 13326 6928
rect 13722 6916 13728 6928
rect 13320 6888 13728 6916
rect 13320 6876 13326 6888
rect 13722 6876 13728 6888
rect 13780 6916 13786 6928
rect 18156 6916 18184 6956
rect 18874 6944 18880 6996
rect 18932 6984 18938 6996
rect 26234 6984 26240 6996
rect 18932 6956 26240 6984
rect 18932 6944 18938 6956
rect 26234 6944 26240 6956
rect 26292 6944 26298 6996
rect 26528 6956 28994 6984
rect 21542 6916 21548 6928
rect 13780 6888 14596 6916
rect 18156 6888 19840 6916
rect 13780 6876 13786 6888
rect 8573 6851 8631 6857
rect 6932 6820 8524 6848
rect 6825 6811 6883 6817
rect 1762 6780 1768 6792
rect 1723 6752 1768 6780
rect 1762 6740 1768 6752
rect 1820 6740 1826 6792
rect 2222 6780 2228 6792
rect 2183 6752 2228 6780
rect 2222 6740 2228 6752
rect 2280 6740 2286 6792
rect 3326 6740 3332 6792
rect 3384 6780 3390 6792
rect 4249 6783 4307 6789
rect 4249 6780 4261 6783
rect 3384 6752 4261 6780
rect 3384 6740 3390 6752
rect 4249 6749 4261 6752
rect 4295 6749 4307 6783
rect 4249 6743 4307 6749
rect 4338 6740 4344 6792
rect 4396 6780 4402 6792
rect 4893 6783 4951 6789
rect 4396 6752 4441 6780
rect 4396 6740 4402 6752
rect 4893 6749 4905 6783
rect 4939 6780 4951 6783
rect 5074 6780 5080 6792
rect 4939 6752 5080 6780
rect 4939 6749 4951 6752
rect 4893 6743 4951 6749
rect 2958 6672 2964 6724
rect 3016 6712 3022 6724
rect 3694 6712 3700 6724
rect 3016 6684 3700 6712
rect 3016 6672 3022 6684
rect 3694 6672 3700 6684
rect 3752 6712 3758 6724
rect 4908 6712 4936 6743
rect 5074 6740 5080 6752
rect 5132 6740 5138 6792
rect 5534 6780 5540 6792
rect 5495 6752 5540 6780
rect 5534 6740 5540 6752
rect 5592 6740 5598 6792
rect 5718 6740 5724 6792
rect 5776 6780 5782 6792
rect 6181 6783 6239 6789
rect 6181 6780 6193 6783
rect 5776 6752 6193 6780
rect 5776 6740 5782 6752
rect 6181 6749 6193 6752
rect 6227 6749 6239 6783
rect 6181 6743 6239 6749
rect 6273 6783 6331 6789
rect 6273 6749 6285 6783
rect 6319 6749 6331 6783
rect 6273 6743 6331 6749
rect 3752 6684 4936 6712
rect 6288 6712 6316 6743
rect 7006 6712 7012 6724
rect 6288 6684 7012 6712
rect 3752 6672 3758 6684
rect 7006 6672 7012 6684
rect 7064 6672 7070 6724
rect 7101 6715 7159 6721
rect 7101 6681 7113 6715
rect 7147 6681 7159 6715
rect 7101 6675 7159 6681
rect 1486 6604 1492 6656
rect 1544 6644 1550 6656
rect 1581 6647 1639 6653
rect 1581 6644 1593 6647
rect 1544 6616 1593 6644
rect 1544 6604 1550 6616
rect 1581 6613 1593 6616
rect 1627 6613 1639 6647
rect 1581 6607 1639 6613
rect 6822 6604 6828 6656
rect 6880 6644 6886 6656
rect 7116 6644 7144 6675
rect 7558 6672 7564 6724
rect 7616 6672 7622 6724
rect 8496 6712 8524 6820
rect 8573 6817 8585 6851
rect 8619 6848 8631 6851
rect 12066 6848 12072 6860
rect 8619 6820 12072 6848
rect 8619 6817 8631 6820
rect 8573 6811 8631 6817
rect 12066 6808 12072 6820
rect 12124 6808 12130 6860
rect 12342 6808 12348 6860
rect 12400 6848 12406 6860
rect 12400 6820 13860 6848
rect 12400 6808 12406 6820
rect 8662 6740 8668 6792
rect 8720 6780 8726 6792
rect 9677 6783 9735 6789
rect 9677 6780 9689 6783
rect 8720 6752 9689 6780
rect 8720 6740 8726 6752
rect 9677 6749 9689 6752
rect 9723 6749 9735 6783
rect 9677 6743 9735 6749
rect 10134 6740 10140 6792
rect 10192 6780 10198 6792
rect 10321 6783 10379 6789
rect 10321 6780 10333 6783
rect 10192 6752 10333 6780
rect 10192 6740 10198 6752
rect 10321 6749 10333 6752
rect 10367 6749 10379 6783
rect 10321 6743 10379 6749
rect 11149 6783 11207 6789
rect 11149 6749 11161 6783
rect 11195 6780 11207 6783
rect 11698 6780 11704 6792
rect 11195 6752 11704 6780
rect 11195 6749 11207 6752
rect 11149 6743 11207 6749
rect 11698 6740 11704 6752
rect 11756 6740 11762 6792
rect 8496 6684 11928 6712
rect 6880 6616 7144 6644
rect 6880 6604 6886 6616
rect 8478 6604 8484 6656
rect 8536 6644 8542 6656
rect 9398 6644 9404 6656
rect 8536 6616 9404 6644
rect 8536 6604 8542 6616
rect 9398 6604 9404 6616
rect 9456 6604 9462 6656
rect 9766 6644 9772 6656
rect 9727 6616 9772 6644
rect 9766 6604 9772 6616
rect 9824 6604 9830 6656
rect 11900 6644 11928 6684
rect 11974 6672 11980 6724
rect 12032 6712 12038 6724
rect 12032 6684 12296 6712
rect 12032 6672 12038 6684
rect 12066 6644 12072 6656
rect 11900 6616 12072 6644
rect 12066 6604 12072 6616
rect 12124 6604 12130 6656
rect 12268 6644 12296 6684
rect 12434 6672 12440 6724
rect 12492 6672 12498 6724
rect 13449 6647 13507 6653
rect 13449 6644 13461 6647
rect 12268 6616 13461 6644
rect 13449 6613 13461 6616
rect 13495 6613 13507 6647
rect 13832 6644 13860 6820
rect 14182 6808 14188 6860
rect 14240 6848 14246 6860
rect 14461 6851 14519 6857
rect 14461 6848 14473 6851
rect 14240 6820 14473 6848
rect 14240 6808 14246 6820
rect 14461 6817 14473 6820
rect 14507 6817 14519 6851
rect 14568 6848 14596 6888
rect 14737 6851 14795 6857
rect 14737 6848 14749 6851
rect 14568 6820 14749 6848
rect 14461 6811 14519 6817
rect 14737 6817 14749 6820
rect 14783 6817 14795 6851
rect 14737 6811 14795 6817
rect 16022 6808 16028 6860
rect 16080 6848 16086 6860
rect 16209 6851 16267 6857
rect 16209 6848 16221 6851
rect 16080 6820 16221 6848
rect 16080 6808 16086 6820
rect 16209 6817 16221 6820
rect 16255 6817 16267 6851
rect 16209 6811 16267 6817
rect 16853 6851 16911 6857
rect 16853 6817 16865 6851
rect 16899 6848 16911 6851
rect 17218 6848 17224 6860
rect 16899 6820 17224 6848
rect 16899 6817 16911 6820
rect 16853 6811 16911 6817
rect 17218 6808 17224 6820
rect 17276 6808 17282 6860
rect 17494 6808 17500 6860
rect 17552 6848 17558 6860
rect 18877 6851 18935 6857
rect 18877 6848 18889 6851
rect 17552 6820 18889 6848
rect 17552 6808 17558 6820
rect 18877 6817 18889 6820
rect 18923 6817 18935 6851
rect 18877 6811 18935 6817
rect 18892 6780 18920 6811
rect 19426 6808 19432 6860
rect 19484 6848 19490 6860
rect 19702 6848 19708 6860
rect 19484 6820 19708 6848
rect 19484 6808 19490 6820
rect 19702 6808 19708 6820
rect 19760 6808 19766 6860
rect 19812 6848 19840 6888
rect 21008 6888 21548 6916
rect 21008 6848 21036 6888
rect 21542 6876 21548 6888
rect 21600 6876 21606 6928
rect 25958 6916 25964 6928
rect 21652 6888 22140 6916
rect 19812 6820 21036 6848
rect 21174 6808 21180 6860
rect 21232 6848 21238 6860
rect 21652 6848 21680 6888
rect 22002 6848 22008 6860
rect 21232 6820 21680 6848
rect 21963 6820 22008 6848
rect 21232 6808 21238 6820
rect 22002 6808 22008 6820
rect 22060 6808 22066 6860
rect 22112 6848 22140 6888
rect 24872 6888 25964 6916
rect 24872 6848 24900 6888
rect 25958 6876 25964 6888
rect 26016 6876 26022 6928
rect 25222 6848 25228 6860
rect 22112 6820 23244 6848
rect 19610 6780 19616 6792
rect 18892 6752 19616 6780
rect 19610 6740 19616 6752
rect 19668 6740 19674 6792
rect 21266 6740 21272 6792
rect 21324 6780 21330 6792
rect 21913 6783 21971 6789
rect 21324 6752 21680 6780
rect 21324 6740 21330 6752
rect 14844 6684 15226 6712
rect 14844 6644 14872 6684
rect 18138 6672 18144 6724
rect 18196 6672 18202 6724
rect 19978 6712 19984 6724
rect 19939 6684 19984 6712
rect 19978 6672 19984 6684
rect 20036 6672 20042 6724
rect 21542 6712 21548 6724
rect 21206 6684 21548 6712
rect 21542 6672 21548 6684
rect 21600 6672 21606 6724
rect 21652 6712 21680 6752
rect 21913 6749 21925 6783
rect 21959 6780 21971 6783
rect 22370 6780 22376 6792
rect 21959 6752 22376 6780
rect 21959 6749 21971 6752
rect 21913 6743 21971 6749
rect 22370 6740 22376 6752
rect 22428 6740 22434 6792
rect 22557 6783 22615 6789
rect 22557 6749 22569 6783
rect 22603 6780 22615 6783
rect 23014 6780 23020 6792
rect 22603 6752 23020 6780
rect 22603 6749 22615 6752
rect 22557 6743 22615 6749
rect 23014 6740 23020 6752
rect 23072 6740 23078 6792
rect 23216 6789 23244 6820
rect 24044 6820 24900 6848
rect 25183 6820 25228 6848
rect 24044 6789 24072 6820
rect 25222 6808 25228 6820
rect 25280 6848 25286 6860
rect 26142 6848 26148 6860
rect 25280 6820 26148 6848
rect 25280 6808 25286 6820
rect 26142 6808 26148 6820
rect 26200 6808 26206 6860
rect 26528 6857 26556 6956
rect 26970 6916 26976 6928
rect 26804 6888 26976 6916
rect 26513 6851 26571 6857
rect 26513 6817 26525 6851
rect 26559 6817 26571 6851
rect 26513 6811 26571 6817
rect 26694 6808 26700 6860
rect 26752 6848 26758 6860
rect 26804 6857 26832 6888
rect 26970 6876 26976 6888
rect 27028 6876 27034 6928
rect 26789 6851 26847 6857
rect 26789 6848 26801 6851
rect 26752 6820 26801 6848
rect 26752 6808 26758 6820
rect 26789 6817 26801 6820
rect 26835 6817 26847 6851
rect 28966 6848 28994 6956
rect 30466 6848 30472 6860
rect 28966 6820 30472 6848
rect 26789 6811 26847 6817
rect 30466 6808 30472 6820
rect 30524 6808 30530 6860
rect 23201 6783 23259 6789
rect 23201 6749 23213 6783
rect 23247 6749 23259 6783
rect 23201 6743 23259 6749
rect 24029 6783 24087 6789
rect 24029 6749 24041 6783
rect 24075 6749 24087 6783
rect 24029 6743 24087 6749
rect 26326 6740 26332 6792
rect 26384 6740 26390 6792
rect 27982 6780 27988 6792
rect 27943 6752 27988 6780
rect 27982 6740 27988 6752
rect 28040 6740 28046 6792
rect 28442 6740 28448 6792
rect 28500 6780 28506 6792
rect 28629 6783 28687 6789
rect 28629 6780 28641 6783
rect 28500 6752 28641 6780
rect 28500 6740 28506 6752
rect 28629 6749 28641 6752
rect 28675 6749 28687 6783
rect 28629 6743 28687 6749
rect 24946 6712 24952 6724
rect 21652 6684 23888 6712
rect 24907 6684 24952 6712
rect 13832 6616 14872 6644
rect 13449 6607 13507 6613
rect 17402 6604 17408 6656
rect 17460 6644 17466 6656
rect 21453 6647 21511 6653
rect 21453 6644 21465 6647
rect 17460 6616 21465 6644
rect 17460 6604 17466 6616
rect 21453 6613 21465 6616
rect 21499 6644 21511 6647
rect 22002 6644 22008 6656
rect 21499 6616 22008 6644
rect 21499 6613 21511 6616
rect 21453 6607 21511 6613
rect 22002 6604 22008 6616
rect 22060 6604 22066 6656
rect 22186 6604 22192 6656
rect 22244 6644 22250 6656
rect 22649 6647 22707 6653
rect 22649 6644 22661 6647
rect 22244 6616 22661 6644
rect 22244 6604 22250 6616
rect 22649 6613 22661 6616
rect 22695 6613 22707 6647
rect 22649 6607 22707 6613
rect 23106 6604 23112 6656
rect 23164 6644 23170 6656
rect 23860 6653 23888 6684
rect 24946 6672 24952 6684
rect 25004 6672 25010 6724
rect 25041 6715 25099 6721
rect 25041 6681 25053 6715
rect 25087 6681 25099 6715
rect 26344 6712 26372 6740
rect 26582 6715 26640 6721
rect 26582 6712 26594 6715
rect 26344 6684 26594 6712
rect 25041 6675 25099 6681
rect 26582 6681 26594 6684
rect 26628 6681 26640 6715
rect 26582 6675 26640 6681
rect 23293 6647 23351 6653
rect 23293 6644 23305 6647
rect 23164 6616 23305 6644
rect 23164 6604 23170 6616
rect 23293 6613 23305 6616
rect 23339 6613 23351 6647
rect 23293 6607 23351 6613
rect 23845 6647 23903 6653
rect 23845 6613 23857 6647
rect 23891 6613 23903 6647
rect 25056 6644 25084 6675
rect 28077 6647 28135 6653
rect 28077 6644 28089 6647
rect 25056 6616 28089 6644
rect 23845 6607 23903 6613
rect 28077 6613 28089 6616
rect 28123 6613 28135 6647
rect 28718 6644 28724 6656
rect 28679 6616 28724 6644
rect 28077 6607 28135 6613
rect 28718 6604 28724 6616
rect 28776 6604 28782 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 5902 6440 5908 6452
rect 5863 6412 5908 6440
rect 5902 6400 5908 6412
rect 5960 6400 5966 6452
rect 9950 6440 9956 6452
rect 6564 6412 9956 6440
rect 2958 6372 2964 6384
rect 2919 6344 2964 6372
rect 2958 6332 2964 6344
rect 3016 6332 3022 6384
rect 3881 6375 3939 6381
rect 3881 6341 3893 6375
rect 3927 6372 3939 6375
rect 4062 6372 4068 6384
rect 3927 6344 4068 6372
rect 3927 6341 3939 6344
rect 3881 6335 3939 6341
rect 4062 6332 4068 6344
rect 4120 6332 4126 6384
rect 6564 6381 6592 6412
rect 9950 6400 9956 6412
rect 10008 6400 10014 6452
rect 12710 6440 12716 6452
rect 10244 6412 12716 6440
rect 6549 6375 6607 6381
rect 6549 6341 6561 6375
rect 6595 6341 6607 6375
rect 6549 6335 6607 6341
rect 7098 6332 7104 6384
rect 7156 6372 7162 6384
rect 8110 6372 8116 6384
rect 7156 6344 8116 6372
rect 7156 6332 7162 6344
rect 8110 6332 8116 6344
rect 8168 6332 8174 6384
rect 9214 6372 9220 6384
rect 8680 6344 9220 6372
rect 2133 6307 2191 6313
rect 2133 6273 2145 6307
rect 2179 6273 2191 6307
rect 2133 6267 2191 6273
rect 4525 6307 4583 6313
rect 4525 6273 4537 6307
rect 4571 6304 4583 6307
rect 5169 6307 5227 6313
rect 5169 6304 5181 6307
rect 4571 6276 5181 6304
rect 4571 6273 4583 6276
rect 4525 6267 4583 6273
rect 5169 6273 5181 6276
rect 5215 6304 5227 6307
rect 5534 6304 5540 6316
rect 5215 6276 5540 6304
rect 5215 6273 5227 6276
rect 5169 6267 5227 6273
rect 2148 6168 2176 6267
rect 2222 6196 2228 6248
rect 2280 6236 2286 6248
rect 2869 6239 2927 6245
rect 2869 6236 2881 6239
rect 2280 6208 2881 6236
rect 2280 6196 2286 6208
rect 2869 6205 2881 6208
rect 2915 6205 2927 6239
rect 2869 6199 2927 6205
rect 4540 6168 4568 6267
rect 5534 6264 5540 6276
rect 5592 6304 5598 6316
rect 5718 6304 5724 6316
rect 5592 6276 5724 6304
rect 5592 6264 5598 6276
rect 5718 6264 5724 6276
rect 5776 6304 5782 6316
rect 5813 6307 5871 6313
rect 5813 6304 5825 6307
rect 5776 6276 5825 6304
rect 5776 6264 5782 6276
rect 5813 6273 5825 6276
rect 5859 6273 5871 6307
rect 5813 6267 5871 6273
rect 7024 6276 7972 6304
rect 5261 6239 5319 6245
rect 5261 6205 5273 6239
rect 5307 6236 5319 6239
rect 7024 6236 7052 6276
rect 5307 6208 7052 6236
rect 5307 6205 5319 6208
rect 5261 6199 5319 6205
rect 7098 6196 7104 6248
rect 7156 6236 7162 6248
rect 7285 6239 7343 6245
rect 7285 6236 7297 6239
rect 7156 6208 7297 6236
rect 7156 6196 7162 6208
rect 7285 6205 7297 6208
rect 7331 6205 7343 6239
rect 7944 6236 7972 6276
rect 8018 6264 8024 6316
rect 8076 6304 8082 6316
rect 8570 6304 8576 6316
rect 8076 6276 8576 6304
rect 8076 6264 8082 6276
rect 8570 6264 8576 6276
rect 8628 6264 8634 6316
rect 8680 6313 8708 6344
rect 9214 6332 9220 6344
rect 9272 6332 9278 6384
rect 9398 6332 9404 6384
rect 9456 6332 9462 6384
rect 8665 6307 8723 6313
rect 8665 6273 8677 6307
rect 8711 6273 8723 6307
rect 8665 6267 8723 6273
rect 10244 6236 10272 6412
rect 12710 6400 12716 6412
rect 12768 6400 12774 6452
rect 15194 6440 15200 6452
rect 13924 6412 15200 6440
rect 10318 6332 10324 6384
rect 10376 6372 10382 6384
rect 11977 6375 12035 6381
rect 11977 6372 11989 6375
rect 10376 6344 11989 6372
rect 10376 6332 10382 6344
rect 11977 6341 11989 6344
rect 12023 6341 12035 6375
rect 11977 6335 12035 6341
rect 12434 6332 12440 6384
rect 12492 6332 12498 6384
rect 10778 6264 10784 6316
rect 10836 6304 10842 6316
rect 10965 6307 11023 6313
rect 10965 6304 10977 6307
rect 10836 6276 10977 6304
rect 10836 6264 10842 6276
rect 10965 6273 10977 6276
rect 11011 6273 11023 6307
rect 10965 6267 11023 6273
rect 7944 6208 10272 6236
rect 10413 6239 10471 6245
rect 7285 6199 7343 6205
rect 10413 6205 10425 6239
rect 10459 6236 10471 6239
rect 11514 6236 11520 6248
rect 10459 6208 11520 6236
rect 10459 6205 10471 6208
rect 10413 6199 10471 6205
rect 2148 6140 4568 6168
rect 4617 6171 4675 6177
rect 4617 6137 4629 6171
rect 4663 6168 4675 6171
rect 8478 6168 8484 6180
rect 4663 6140 8484 6168
rect 4663 6137 4675 6140
rect 4617 6131 4675 6137
rect 8478 6128 8484 6140
rect 8536 6128 8542 6180
rect 8662 6128 8668 6180
rect 8720 6168 8726 6180
rect 8720 6140 8800 6168
rect 8720 6128 8726 6140
rect 2225 6103 2283 6109
rect 2225 6069 2237 6103
rect 2271 6100 2283 6103
rect 6546 6100 6552 6112
rect 2271 6072 6552 6100
rect 2271 6069 2283 6072
rect 2225 6063 2283 6069
rect 6546 6060 6552 6072
rect 6604 6060 6610 6112
rect 8772 6100 8800 6140
rect 9950 6128 9956 6180
rect 10008 6168 10014 6180
rect 10428 6168 10456 6199
rect 11514 6196 11520 6208
rect 11572 6196 11578 6248
rect 11698 6236 11704 6248
rect 11659 6208 11704 6236
rect 11698 6196 11704 6208
rect 11756 6196 11762 6248
rect 13924 6236 13952 6412
rect 15194 6400 15200 6412
rect 15252 6400 15258 6452
rect 15749 6443 15807 6449
rect 15749 6409 15761 6443
rect 15795 6440 15807 6443
rect 16758 6440 16764 6452
rect 15795 6412 16764 6440
rect 15795 6409 15807 6412
rect 15749 6403 15807 6409
rect 16758 6400 16764 6412
rect 16816 6400 16822 6452
rect 19058 6440 19064 6452
rect 17512 6412 19064 6440
rect 14182 6372 14188 6384
rect 14016 6344 14188 6372
rect 14016 6313 14044 6344
rect 14182 6332 14188 6344
rect 14240 6332 14246 6384
rect 14277 6375 14335 6381
rect 14277 6341 14289 6375
rect 14323 6372 14335 6375
rect 14366 6372 14372 6384
rect 14323 6344 14372 6372
rect 14323 6341 14335 6344
rect 14277 6335 14335 6341
rect 14366 6332 14372 6344
rect 14424 6332 14430 6384
rect 15286 6332 15292 6384
rect 15344 6332 15350 6384
rect 17512 6381 17540 6412
rect 19058 6400 19064 6412
rect 19116 6400 19122 6452
rect 19334 6400 19340 6452
rect 19392 6440 19398 6452
rect 20254 6440 20260 6452
rect 19392 6412 20260 6440
rect 19392 6400 19398 6412
rect 20254 6400 20260 6412
rect 20312 6400 20318 6452
rect 23382 6440 23388 6452
rect 20364 6412 23388 6440
rect 17497 6375 17555 6381
rect 17497 6341 17509 6375
rect 17543 6341 17555 6375
rect 20364 6372 20392 6412
rect 23382 6400 23388 6412
rect 23440 6400 23446 6452
rect 23676 6412 27752 6440
rect 22002 6372 22008 6384
rect 18722 6344 20392 6372
rect 21206 6344 22008 6372
rect 17497 6335 17555 6341
rect 22002 6332 22008 6344
rect 22060 6332 22066 6384
rect 23014 6332 23020 6384
rect 23072 6372 23078 6384
rect 23676 6372 23704 6412
rect 23072 6344 23704 6372
rect 23753 6375 23811 6381
rect 23072 6332 23078 6344
rect 23753 6341 23765 6375
rect 23799 6372 23811 6375
rect 24026 6372 24032 6384
rect 23799 6344 24032 6372
rect 23799 6341 23811 6344
rect 23753 6335 23811 6341
rect 24026 6332 24032 6344
rect 24084 6332 24090 6384
rect 25314 6372 25320 6384
rect 25275 6344 25320 6372
rect 25314 6332 25320 6344
rect 25372 6332 25378 6384
rect 25409 6375 25467 6381
rect 25409 6341 25421 6375
rect 25455 6372 25467 6375
rect 27522 6372 27528 6384
rect 25455 6344 27528 6372
rect 25455 6341 25467 6344
rect 25409 6335 25467 6341
rect 27522 6332 27528 6344
rect 27580 6332 27586 6384
rect 27724 6372 27752 6412
rect 27798 6400 27804 6452
rect 27856 6440 27862 6452
rect 27985 6443 28043 6449
rect 27985 6440 27997 6443
rect 27856 6412 27997 6440
rect 27856 6400 27862 6412
rect 27985 6409 27997 6412
rect 28031 6409 28043 6443
rect 27985 6403 28043 6409
rect 31478 6372 31484 6384
rect 27724 6344 31484 6372
rect 31478 6332 31484 6344
rect 31536 6332 31542 6384
rect 14001 6307 14059 6313
rect 14001 6273 14013 6307
rect 14047 6273 14059 6307
rect 17218 6304 17224 6316
rect 17179 6276 17224 6304
rect 14001 6267 14059 6273
rect 17218 6264 17224 6276
rect 17276 6264 17282 6316
rect 19334 6304 19340 6316
rect 18708 6276 19340 6304
rect 18708 6236 18736 6276
rect 19334 6264 19340 6276
rect 19392 6264 19398 6316
rect 19426 6264 19432 6316
rect 19484 6304 19490 6316
rect 19705 6307 19763 6313
rect 19705 6304 19717 6307
rect 19484 6276 19717 6304
rect 19484 6264 19490 6276
rect 19705 6273 19717 6276
rect 19751 6273 19763 6307
rect 19705 6267 19763 6273
rect 22094 6264 22100 6316
rect 22152 6304 22158 6316
rect 22373 6307 22431 6313
rect 22373 6304 22385 6307
rect 22152 6276 22385 6304
rect 22152 6264 22158 6276
rect 22373 6273 22385 6276
rect 22419 6273 22431 6307
rect 27154 6304 27160 6316
rect 27115 6276 27160 6304
rect 22373 6267 22431 6273
rect 27154 6264 27160 6276
rect 27212 6264 27218 6316
rect 27246 6264 27252 6316
rect 27304 6304 27310 6316
rect 27433 6307 27491 6313
rect 27433 6304 27445 6307
rect 27304 6276 27445 6304
rect 27304 6264 27310 6276
rect 27433 6273 27445 6276
rect 27479 6273 27491 6307
rect 27433 6267 27491 6273
rect 27893 6307 27951 6313
rect 27893 6273 27905 6307
rect 27939 6273 27951 6307
rect 27893 6267 27951 6273
rect 28537 6307 28595 6313
rect 28537 6273 28549 6307
rect 28583 6273 28595 6307
rect 30190 6304 30196 6316
rect 30151 6276 30196 6304
rect 28537 6267 28595 6273
rect 11808 6208 13952 6236
rect 14108 6208 18736 6236
rect 18969 6239 19027 6245
rect 10008 6140 10456 6168
rect 11057 6171 11115 6177
rect 10008 6128 10014 6140
rect 11057 6137 11069 6171
rect 11103 6168 11115 6171
rect 11808 6168 11836 6208
rect 11103 6140 11836 6168
rect 13449 6171 13507 6177
rect 11103 6137 11115 6140
rect 11057 6131 11115 6137
rect 13449 6137 13461 6171
rect 13495 6168 13507 6171
rect 14108 6168 14136 6208
rect 18969 6205 18981 6239
rect 19015 6236 19027 6239
rect 19981 6239 20039 6245
rect 19981 6236 19993 6239
rect 19015 6208 19993 6236
rect 19015 6205 19027 6208
rect 18969 6199 19027 6205
rect 19981 6205 19993 6208
rect 20027 6236 20039 6239
rect 22830 6236 22836 6248
rect 20027 6208 22836 6236
rect 20027 6205 20039 6208
rect 19981 6199 20039 6205
rect 22830 6196 22836 6208
rect 22888 6196 22894 6248
rect 23658 6236 23664 6248
rect 23619 6208 23664 6236
rect 23658 6196 23664 6208
rect 23716 6196 23722 6248
rect 23750 6196 23756 6248
rect 23808 6236 23814 6248
rect 23937 6239 23995 6245
rect 23937 6236 23949 6239
rect 23808 6208 23949 6236
rect 23808 6196 23814 6208
rect 23937 6205 23949 6208
rect 23983 6236 23995 6239
rect 24946 6236 24952 6248
rect 23983 6208 24952 6236
rect 23983 6205 23995 6208
rect 23937 6199 23995 6205
rect 24946 6196 24952 6208
rect 25004 6236 25010 6248
rect 25593 6239 25651 6245
rect 25593 6236 25605 6239
rect 25004 6208 25605 6236
rect 25004 6196 25010 6208
rect 25593 6205 25605 6208
rect 25639 6205 25651 6239
rect 25593 6199 25651 6205
rect 26510 6196 26516 6248
rect 26568 6236 26574 6248
rect 27908 6236 27936 6267
rect 26568 6208 27936 6236
rect 28552 6236 28580 6267
rect 30190 6264 30196 6276
rect 30248 6264 30254 6316
rect 35802 6264 35808 6316
rect 35860 6304 35866 6316
rect 36817 6307 36875 6313
rect 36817 6304 36829 6307
rect 35860 6276 36829 6304
rect 35860 6264 35866 6276
rect 36817 6273 36829 6276
rect 36863 6273 36875 6307
rect 36817 6267 36875 6273
rect 34606 6236 34612 6248
rect 28552 6208 34612 6236
rect 26568 6196 26574 6208
rect 34606 6196 34612 6208
rect 34664 6196 34670 6248
rect 19702 6168 19708 6180
rect 13495 6140 14136 6168
rect 18524 6140 19708 6168
rect 13495 6137 13507 6140
rect 13449 6131 13507 6137
rect 8922 6103 8980 6109
rect 8922 6100 8934 6103
rect 8772 6072 8934 6100
rect 8922 6069 8934 6072
rect 8968 6069 8980 6103
rect 8922 6063 8980 6069
rect 9582 6060 9588 6112
rect 9640 6100 9646 6112
rect 13170 6100 13176 6112
rect 9640 6072 13176 6100
rect 9640 6060 9646 6072
rect 13170 6060 13176 6072
rect 13228 6060 13234 6112
rect 13630 6060 13636 6112
rect 13688 6100 13694 6112
rect 18524 6100 18552 6140
rect 19702 6128 19708 6140
rect 19760 6128 19766 6180
rect 21453 6171 21511 6177
rect 21453 6137 21465 6171
rect 21499 6168 21511 6171
rect 21634 6168 21640 6180
rect 21499 6140 21640 6168
rect 21499 6137 21511 6140
rect 21453 6131 21511 6137
rect 21634 6128 21640 6140
rect 21692 6128 21698 6180
rect 22278 6128 22284 6180
rect 22336 6168 22342 6180
rect 23842 6168 23848 6180
rect 22336 6140 23848 6168
rect 22336 6128 22342 6140
rect 23842 6128 23848 6140
rect 23900 6128 23906 6180
rect 25314 6128 25320 6180
rect 25372 6168 25378 6180
rect 28629 6171 28687 6177
rect 28629 6168 28641 6171
rect 25372 6140 28641 6168
rect 25372 6128 25378 6140
rect 28629 6137 28641 6140
rect 28675 6137 28687 6171
rect 28629 6131 28687 6137
rect 13688 6072 18552 6100
rect 13688 6060 13694 6072
rect 19334 6060 19340 6112
rect 19392 6100 19398 6112
rect 21910 6100 21916 6112
rect 19392 6072 21916 6100
rect 19392 6060 19398 6072
rect 21910 6060 21916 6072
rect 21968 6060 21974 6112
rect 22557 6103 22615 6109
rect 22557 6069 22569 6103
rect 22603 6100 22615 6103
rect 23014 6100 23020 6112
rect 22603 6072 23020 6100
rect 22603 6069 22615 6072
rect 22557 6063 22615 6069
rect 23014 6060 23020 6072
rect 23072 6060 23078 6112
rect 23198 6060 23204 6112
rect 23256 6100 23262 6112
rect 25958 6100 25964 6112
rect 23256 6072 25964 6100
rect 23256 6060 23262 6072
rect 25958 6060 25964 6072
rect 26016 6060 26022 6112
rect 26326 6060 26332 6112
rect 26384 6100 26390 6112
rect 28258 6100 28264 6112
rect 26384 6072 28264 6100
rect 26384 6060 26390 6072
rect 28258 6060 28264 6072
rect 28316 6060 28322 6112
rect 30009 6103 30067 6109
rect 30009 6069 30021 6103
rect 30055 6100 30067 6103
rect 33410 6100 33416 6112
rect 30055 6072 33416 6100
rect 30055 6069 30067 6072
rect 30009 6063 30067 6069
rect 33410 6060 33416 6072
rect 33468 6060 33474 6112
rect 36633 6103 36691 6109
rect 36633 6069 36645 6103
rect 36679 6100 36691 6103
rect 38010 6100 38016 6112
rect 36679 6072 38016 6100
rect 36679 6069 36691 6072
rect 36633 6063 36691 6069
rect 38010 6060 38016 6072
rect 38068 6060 38074 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 2222 5856 2228 5908
rect 2280 5896 2286 5908
rect 2685 5899 2743 5905
rect 2685 5896 2697 5899
rect 2280 5868 2697 5896
rect 2280 5856 2286 5868
rect 2685 5865 2697 5868
rect 2731 5865 2743 5899
rect 2685 5859 2743 5865
rect 4788 5899 4846 5905
rect 4788 5865 4800 5899
rect 4834 5896 4846 5899
rect 5994 5896 6000 5908
rect 4834 5868 6000 5896
rect 4834 5865 4846 5868
rect 4788 5859 4846 5865
rect 5994 5856 6000 5868
rect 6052 5856 6058 5908
rect 6270 5896 6276 5908
rect 6231 5868 6276 5896
rect 6270 5856 6276 5868
rect 6328 5856 6334 5908
rect 7742 5896 7748 5908
rect 6656 5868 7748 5896
rect 1949 5831 2007 5837
rect 1949 5797 1961 5831
rect 1995 5828 2007 5831
rect 3234 5828 3240 5840
rect 1995 5800 3240 5828
rect 1995 5797 2007 5800
rect 1949 5791 2007 5797
rect 3234 5788 3240 5800
rect 3292 5788 3298 5840
rect 6656 5828 6684 5868
rect 7742 5856 7748 5868
rect 7800 5856 7806 5908
rect 8110 5856 8116 5908
rect 8168 5896 8174 5908
rect 8168 5868 13584 5896
rect 8168 5856 8174 5868
rect 8478 5828 8484 5840
rect 6288 5800 6684 5828
rect 8439 5800 8484 5828
rect 2133 5695 2191 5701
rect 2133 5661 2145 5695
rect 2179 5692 2191 5695
rect 2222 5692 2228 5704
rect 2179 5664 2228 5692
rect 2179 5661 2191 5664
rect 2133 5655 2191 5661
rect 2222 5652 2228 5664
rect 2280 5652 2286 5704
rect 2406 5652 2412 5704
rect 2464 5692 2470 5704
rect 2593 5695 2651 5701
rect 2593 5692 2605 5695
rect 2464 5664 2605 5692
rect 2464 5652 2470 5664
rect 2593 5661 2605 5664
rect 2639 5661 2651 5695
rect 2593 5655 2651 5661
rect 3237 5695 3295 5701
rect 3237 5661 3249 5695
rect 3283 5692 3295 5695
rect 3326 5692 3332 5704
rect 3283 5664 3332 5692
rect 3283 5661 3295 5664
rect 3237 5655 3295 5661
rect 3326 5652 3332 5664
rect 3384 5652 3390 5704
rect 4522 5692 4528 5704
rect 4483 5664 4528 5692
rect 4522 5652 4528 5664
rect 4580 5652 4586 5704
rect 5258 5584 5264 5636
rect 5316 5584 5322 5636
rect 6288 5624 6316 5800
rect 8478 5788 8484 5800
rect 8536 5788 8542 5840
rect 11057 5831 11115 5837
rect 11057 5797 11069 5831
rect 11103 5828 11115 5831
rect 11330 5828 11336 5840
rect 11103 5800 11336 5828
rect 11103 5797 11115 5800
rect 11057 5791 11115 5797
rect 11330 5788 11336 5800
rect 11388 5788 11394 5840
rect 11974 5788 11980 5840
rect 12032 5788 12038 5840
rect 13556 5828 13584 5868
rect 14366 5856 14372 5908
rect 14424 5896 14430 5908
rect 14424 5868 22232 5896
rect 14424 5856 14430 5868
rect 22204 5828 22232 5868
rect 22278 5856 22284 5908
rect 22336 5896 22342 5908
rect 22373 5899 22431 5905
rect 22373 5896 22385 5899
rect 22336 5868 22385 5896
rect 22336 5856 22342 5868
rect 22373 5865 22385 5868
rect 22419 5865 22431 5899
rect 22373 5859 22431 5865
rect 22462 5856 22468 5908
rect 22520 5896 22526 5908
rect 26326 5896 26332 5908
rect 22520 5868 26332 5896
rect 22520 5856 22526 5868
rect 26326 5856 26332 5868
rect 26384 5856 26390 5908
rect 26602 5856 26608 5908
rect 26660 5896 26666 5908
rect 26881 5899 26939 5905
rect 26881 5896 26893 5899
rect 26660 5868 26893 5896
rect 26660 5856 26666 5868
rect 26881 5865 26893 5868
rect 26927 5865 26939 5899
rect 27522 5896 27528 5908
rect 27483 5868 27528 5896
rect 26881 5859 26939 5865
rect 27522 5856 27528 5868
rect 27580 5856 27586 5908
rect 31846 5828 31852 5840
rect 13556 5800 14504 5828
rect 6546 5720 6552 5772
rect 6604 5720 6610 5772
rect 6730 5760 6736 5772
rect 6691 5732 6736 5760
rect 6730 5720 6736 5732
rect 6788 5720 6794 5772
rect 7006 5720 7012 5772
rect 7064 5760 7070 5772
rect 8294 5760 8300 5772
rect 7064 5732 8300 5760
rect 7064 5720 7070 5732
rect 8294 5720 8300 5732
rect 8352 5720 8358 5772
rect 9306 5760 9312 5772
rect 9219 5732 9312 5760
rect 9306 5720 9312 5732
rect 9364 5760 9370 5772
rect 11992 5760 12020 5788
rect 12253 5763 12311 5769
rect 12253 5760 12265 5763
rect 9364 5732 11836 5760
rect 11992 5732 12265 5760
rect 9364 5720 9370 5732
rect 6196 5596 6316 5624
rect 3329 5559 3387 5565
rect 3329 5525 3341 5559
rect 3375 5556 3387 5559
rect 6196 5556 6224 5596
rect 3375 5528 6224 5556
rect 6564 5556 6592 5720
rect 11808 5704 11836 5732
rect 12253 5729 12265 5732
rect 12299 5729 12311 5763
rect 12253 5723 12311 5729
rect 13722 5720 13728 5772
rect 13780 5760 13786 5772
rect 13780 5732 13825 5760
rect 13780 5720 13786 5732
rect 14182 5720 14188 5772
rect 14240 5760 14246 5772
rect 14369 5763 14427 5769
rect 14369 5760 14381 5763
rect 14240 5732 14381 5760
rect 14240 5720 14246 5732
rect 14369 5729 14381 5732
rect 14415 5729 14427 5763
rect 14476 5760 14504 5800
rect 15672 5800 17264 5828
rect 15672 5760 15700 5800
rect 14476 5732 15700 5760
rect 16117 5763 16175 5769
rect 14369 5723 14427 5729
rect 16117 5729 16129 5763
rect 16163 5760 16175 5763
rect 16206 5760 16212 5772
rect 16163 5732 16212 5760
rect 16163 5729 16175 5732
rect 16117 5723 16175 5729
rect 16206 5720 16212 5732
rect 16264 5720 16270 5772
rect 17126 5760 17132 5772
rect 17087 5732 17132 5760
rect 17126 5720 17132 5732
rect 17184 5720 17190 5772
rect 17236 5760 17264 5800
rect 18432 5800 19932 5828
rect 22204 5800 31852 5828
rect 18432 5760 18460 5800
rect 17236 5732 18460 5760
rect 18877 5763 18935 5769
rect 18877 5729 18889 5763
rect 18923 5760 18935 5763
rect 18966 5760 18972 5772
rect 18923 5732 18972 5760
rect 18923 5729 18935 5732
rect 18877 5723 18935 5729
rect 18966 5720 18972 5732
rect 19024 5720 19030 5772
rect 19426 5720 19432 5772
rect 19484 5760 19490 5772
rect 19797 5763 19855 5769
rect 19797 5760 19809 5763
rect 19484 5732 19809 5760
rect 19484 5720 19490 5732
rect 19797 5729 19809 5732
rect 19843 5729 19855 5763
rect 19904 5760 19932 5800
rect 31846 5788 31852 5800
rect 31904 5788 31910 5840
rect 21910 5760 21916 5772
rect 19904 5732 21916 5760
rect 19797 5723 19855 5729
rect 21910 5720 21916 5732
rect 21968 5720 21974 5772
rect 23014 5760 23020 5772
rect 22975 5732 23020 5760
rect 23014 5720 23020 5732
rect 23072 5720 23078 5772
rect 23658 5720 23664 5772
rect 23716 5760 23722 5772
rect 24673 5763 24731 5769
rect 24673 5760 24685 5763
rect 23716 5732 24685 5760
rect 23716 5720 23722 5732
rect 24673 5729 24685 5732
rect 24719 5760 24731 5763
rect 28718 5760 28724 5772
rect 24719 5732 28724 5760
rect 24719 5729 24731 5732
rect 24673 5723 24731 5729
rect 28718 5720 28724 5732
rect 28776 5720 28782 5772
rect 28810 5720 28816 5772
rect 28868 5760 28874 5772
rect 28868 5732 35894 5760
rect 28868 5720 28874 5732
rect 11790 5652 11796 5704
rect 11848 5692 11854 5704
rect 11977 5695 12035 5701
rect 11977 5692 11989 5695
rect 11848 5664 11989 5692
rect 11848 5652 11854 5664
rect 11977 5661 11989 5664
rect 12023 5661 12035 5695
rect 21450 5692 21456 5704
rect 21206 5664 21456 5692
rect 11977 5655 12035 5661
rect 21450 5652 21456 5664
rect 21508 5652 21514 5704
rect 22186 5652 22192 5704
rect 22244 5692 22250 5704
rect 22281 5695 22339 5701
rect 22281 5692 22293 5695
rect 22244 5664 22293 5692
rect 22244 5652 22250 5664
rect 22281 5661 22293 5664
rect 22327 5661 22339 5695
rect 22281 5655 22339 5661
rect 25590 5652 25596 5704
rect 25648 5692 25654 5704
rect 26145 5695 26203 5701
rect 26145 5692 26157 5695
rect 25648 5664 26157 5692
rect 25648 5652 25654 5664
rect 26145 5661 26157 5664
rect 26191 5661 26203 5695
rect 26145 5655 26203 5661
rect 26234 5652 26240 5704
rect 26292 5692 26298 5704
rect 26292 5664 26337 5692
rect 26292 5652 26298 5664
rect 26418 5652 26424 5704
rect 26476 5692 26482 5704
rect 26789 5695 26847 5701
rect 26789 5692 26801 5695
rect 26476 5664 26801 5692
rect 26476 5652 26482 5664
rect 26789 5661 26801 5664
rect 26835 5692 26847 5695
rect 27154 5692 27160 5704
rect 26835 5664 27160 5692
rect 26835 5661 26847 5664
rect 26789 5655 26847 5661
rect 27154 5652 27160 5664
rect 27212 5652 27218 5704
rect 27430 5692 27436 5704
rect 27391 5664 27436 5692
rect 27430 5652 27436 5664
rect 27488 5652 27494 5704
rect 27982 5652 27988 5704
rect 28040 5692 28046 5704
rect 28077 5695 28135 5701
rect 28077 5692 28089 5695
rect 28040 5664 28089 5692
rect 28040 5652 28046 5664
rect 28077 5661 28089 5664
rect 28123 5661 28135 5695
rect 29730 5692 29736 5704
rect 29691 5664 29736 5692
rect 28077 5655 28135 5661
rect 29730 5652 29736 5664
rect 29788 5652 29794 5704
rect 35866 5692 35894 5732
rect 38013 5695 38071 5701
rect 38013 5692 38025 5695
rect 35866 5664 38025 5692
rect 38013 5661 38025 5664
rect 38059 5661 38071 5695
rect 38013 5655 38071 5661
rect 6638 5584 6644 5636
rect 6696 5624 6702 5636
rect 7009 5627 7067 5633
rect 7009 5624 7021 5627
rect 6696 5596 7021 5624
rect 6696 5584 6702 5596
rect 7009 5593 7021 5596
rect 7055 5593 7067 5627
rect 9585 5627 9643 5633
rect 9585 5624 9597 5627
rect 7009 5587 7067 5593
rect 7116 5596 7498 5624
rect 8312 5596 9597 5624
rect 7116 5556 7144 5596
rect 6564 5528 7144 5556
rect 3375 5525 3387 5528
rect 3329 5519 3387 5525
rect 7190 5516 7196 5568
rect 7248 5556 7254 5568
rect 8312 5556 8340 5596
rect 9585 5593 9597 5596
rect 9631 5593 9643 5627
rect 9585 5587 9643 5593
rect 9692 5596 10074 5624
rect 7248 5528 8340 5556
rect 7248 5516 7254 5528
rect 9030 5516 9036 5568
rect 9088 5556 9094 5568
rect 9692 5556 9720 5596
rect 12710 5584 12716 5636
rect 12768 5584 12774 5636
rect 14645 5627 14703 5633
rect 14645 5593 14657 5627
rect 14691 5593 14703 5627
rect 14645 5587 14703 5593
rect 9088 5528 9720 5556
rect 9088 5516 9094 5528
rect 11146 5516 11152 5568
rect 11204 5556 11210 5568
rect 14366 5556 14372 5568
rect 11204 5528 14372 5556
rect 11204 5516 11210 5528
rect 14366 5516 14372 5528
rect 14424 5516 14430 5568
rect 14660 5556 14688 5587
rect 15102 5584 15108 5636
rect 15160 5584 15166 5636
rect 17402 5624 17408 5636
rect 17363 5596 17408 5624
rect 17402 5584 17408 5596
rect 17460 5584 17466 5636
rect 20073 5627 20131 5633
rect 18630 5596 20024 5624
rect 15930 5556 15936 5568
rect 14660 5528 15936 5556
rect 15930 5516 15936 5528
rect 15988 5516 15994 5568
rect 18046 5516 18052 5568
rect 18104 5556 18110 5568
rect 18966 5556 18972 5568
rect 18104 5528 18972 5556
rect 18104 5516 18110 5528
rect 18966 5516 18972 5528
rect 19024 5516 19030 5568
rect 19996 5556 20024 5596
rect 20073 5593 20085 5627
rect 20119 5624 20131 5627
rect 20346 5624 20352 5636
rect 20119 5596 20352 5624
rect 20119 5593 20131 5596
rect 20073 5587 20131 5593
rect 20346 5584 20352 5596
rect 20404 5584 20410 5636
rect 23014 5624 23020 5636
rect 21376 5596 23020 5624
rect 21376 5556 21404 5596
rect 23014 5584 23020 5596
rect 23072 5584 23078 5636
rect 23106 5584 23112 5636
rect 23164 5624 23170 5636
rect 23661 5627 23719 5633
rect 23164 5596 23209 5624
rect 23164 5584 23170 5596
rect 23661 5593 23673 5627
rect 23707 5624 23719 5627
rect 24302 5624 24308 5636
rect 23707 5596 24308 5624
rect 23707 5593 23719 5596
rect 23661 5587 23719 5593
rect 24302 5584 24308 5596
rect 24360 5584 24366 5636
rect 24765 5627 24823 5633
rect 24765 5593 24777 5627
rect 24811 5593 24823 5627
rect 25682 5624 25688 5636
rect 25643 5596 25688 5624
rect 24765 5587 24823 5593
rect 21542 5556 21548 5568
rect 19996 5528 21404 5556
rect 21503 5528 21548 5556
rect 21542 5516 21548 5528
rect 21600 5516 21606 5568
rect 22462 5516 22468 5568
rect 22520 5556 22526 5568
rect 24394 5556 24400 5568
rect 22520 5528 24400 5556
rect 22520 5516 22526 5528
rect 24394 5516 24400 5528
rect 24452 5516 24458 5568
rect 24780 5556 24808 5587
rect 25682 5584 25688 5596
rect 25740 5624 25746 5636
rect 25740 5596 26372 5624
rect 25740 5584 25746 5596
rect 26234 5556 26240 5568
rect 24780 5528 26240 5556
rect 26234 5516 26240 5528
rect 26292 5516 26298 5568
rect 26344 5556 26372 5596
rect 27982 5556 27988 5568
rect 26344 5528 27988 5556
rect 27982 5516 27988 5528
rect 28040 5516 28046 5568
rect 28166 5556 28172 5568
rect 28127 5528 28172 5556
rect 28166 5516 28172 5528
rect 28224 5516 28230 5568
rect 28718 5556 28724 5568
rect 28679 5528 28724 5556
rect 28718 5516 28724 5528
rect 28776 5516 28782 5568
rect 29822 5556 29828 5568
rect 29783 5528 29828 5556
rect 29822 5516 29828 5528
rect 29880 5516 29886 5568
rect 38194 5556 38200 5568
rect 38155 5528 38200 5556
rect 38194 5516 38200 5528
rect 38252 5516 38258 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 1673 5355 1731 5361
rect 1673 5321 1685 5355
rect 1719 5352 1731 5355
rect 2130 5352 2136 5364
rect 1719 5324 2136 5352
rect 1719 5321 1731 5324
rect 1673 5315 1731 5321
rect 2130 5312 2136 5324
rect 2188 5312 2194 5364
rect 2409 5355 2467 5361
rect 2409 5321 2421 5355
rect 2455 5352 2467 5355
rect 2958 5352 2964 5364
rect 2455 5324 2964 5352
rect 2455 5321 2467 5324
rect 2409 5315 2467 5321
rect 2958 5312 2964 5324
rect 3016 5312 3022 5364
rect 3697 5355 3755 5361
rect 3697 5321 3709 5355
rect 3743 5352 3755 5355
rect 14550 5352 14556 5364
rect 3743 5324 9260 5352
rect 3743 5321 3755 5324
rect 3697 5315 3755 5321
rect 2222 5284 2228 5296
rect 1596 5256 2228 5284
rect 1596 5225 1624 5256
rect 2222 5244 2228 5256
rect 2280 5284 2286 5296
rect 4614 5284 4620 5296
rect 2280 5256 2774 5284
rect 2280 5244 2286 5256
rect 1581 5219 1639 5225
rect 1581 5185 1593 5219
rect 1627 5185 1639 5219
rect 2314 5216 2320 5228
rect 2275 5188 2320 5216
rect 1581 5179 1639 5185
rect 2314 5176 2320 5188
rect 2372 5176 2378 5228
rect 2746 5080 2774 5256
rect 4264 5256 4620 5284
rect 3145 5219 3203 5225
rect 3145 5185 3157 5219
rect 3191 5216 3203 5219
rect 3326 5216 3332 5228
rect 3191 5188 3332 5216
rect 3191 5185 3203 5188
rect 3145 5179 3203 5185
rect 3326 5176 3332 5188
rect 3384 5176 3390 5228
rect 3602 5216 3608 5228
rect 3563 5188 3608 5216
rect 3602 5176 3608 5188
rect 3660 5176 3666 5228
rect 4264 5225 4292 5256
rect 4614 5244 4620 5256
rect 4672 5244 4678 5296
rect 6086 5284 6092 5296
rect 5750 5256 6092 5284
rect 6086 5244 6092 5256
rect 6144 5244 6150 5296
rect 7190 5284 7196 5296
rect 6564 5256 7196 5284
rect 4249 5219 4307 5225
rect 4249 5185 4261 5219
rect 4295 5185 4307 5219
rect 4249 5179 4307 5185
rect 5994 5176 6000 5228
rect 6052 5216 6058 5228
rect 6564 5225 6592 5256
rect 7190 5244 7196 5256
rect 7248 5244 7254 5296
rect 7466 5284 7472 5296
rect 7427 5256 7472 5284
rect 7466 5244 7472 5256
rect 7524 5244 7530 5296
rect 7558 5244 7564 5296
rect 7616 5284 7622 5296
rect 7616 5256 7958 5284
rect 7616 5244 7622 5256
rect 6549 5219 6607 5225
rect 6549 5216 6561 5219
rect 6052 5188 6561 5216
rect 6052 5176 6058 5188
rect 6549 5185 6561 5188
rect 6595 5185 6607 5219
rect 6549 5179 6607 5185
rect 4522 5108 4528 5160
rect 4580 5148 4586 5160
rect 7190 5148 7196 5160
rect 4580 5120 4625 5148
rect 7151 5120 7196 5148
rect 4580 5108 4586 5120
rect 7190 5108 7196 5120
rect 7248 5108 7254 5160
rect 9232 5148 9260 5324
rect 9692 5324 14556 5352
rect 9692 5293 9720 5324
rect 14550 5312 14556 5324
rect 14608 5312 14614 5364
rect 14642 5312 14648 5364
rect 14700 5352 14706 5364
rect 15930 5352 15936 5364
rect 14700 5324 15792 5352
rect 15891 5324 15936 5352
rect 14700 5312 14706 5324
rect 9677 5287 9735 5293
rect 9677 5253 9689 5287
rect 9723 5253 9735 5287
rect 9677 5247 9735 5253
rect 9950 5244 9956 5296
rect 10008 5284 10014 5296
rect 10008 5256 10166 5284
rect 10008 5244 10014 5256
rect 13446 5244 13452 5296
rect 13504 5284 13510 5296
rect 13725 5287 13783 5293
rect 13725 5284 13737 5287
rect 13504 5256 13737 5284
rect 13504 5244 13510 5256
rect 13725 5253 13737 5256
rect 13771 5253 13783 5287
rect 13725 5247 13783 5253
rect 13814 5244 13820 5296
rect 13872 5284 13878 5296
rect 15764 5284 15792 5324
rect 15930 5312 15936 5324
rect 15988 5312 15994 5364
rect 16114 5312 16120 5364
rect 16172 5352 16178 5364
rect 20070 5352 20076 5364
rect 16172 5324 20076 5352
rect 16172 5312 16178 5324
rect 20070 5312 20076 5324
rect 20128 5312 20134 5364
rect 21910 5352 21916 5364
rect 20180 5324 21916 5352
rect 17221 5287 17279 5293
rect 17221 5284 17233 5287
rect 13872 5256 14950 5284
rect 15764 5256 17233 5284
rect 13872 5244 13878 5256
rect 17221 5253 17233 5256
rect 17267 5253 17279 5287
rect 20180 5284 20208 5324
rect 21910 5312 21916 5324
rect 21968 5312 21974 5364
rect 28537 5355 28595 5361
rect 28537 5352 28549 5355
rect 25332 5324 28549 5352
rect 21634 5284 21640 5296
rect 18446 5256 20208 5284
rect 21022 5256 21640 5284
rect 17221 5247 17279 5253
rect 21634 5244 21640 5256
rect 21692 5244 21698 5296
rect 21726 5244 21732 5296
rect 21784 5284 21790 5296
rect 21784 5256 22508 5284
rect 21784 5244 21790 5256
rect 9306 5176 9312 5228
rect 9364 5216 9370 5228
rect 9401 5219 9459 5225
rect 9401 5216 9413 5219
rect 9364 5188 9413 5216
rect 9364 5176 9370 5188
rect 9401 5185 9413 5188
rect 9447 5185 9459 5219
rect 13538 5216 13544 5228
rect 13110 5188 13544 5216
rect 9401 5179 9459 5185
rect 13538 5176 13544 5188
rect 13596 5176 13602 5228
rect 18874 5216 18880 5228
rect 18432 5188 18880 5216
rect 10042 5148 10048 5160
rect 9232 5120 10048 5148
rect 10042 5108 10048 5120
rect 10100 5108 10106 5160
rect 11146 5148 11152 5160
rect 11107 5120 11152 5148
rect 11146 5108 11152 5120
rect 11204 5108 11210 5160
rect 11698 5148 11704 5160
rect 11659 5120 11704 5148
rect 11698 5108 11704 5120
rect 11756 5108 11762 5160
rect 11977 5151 12035 5157
rect 11977 5117 11989 5151
rect 12023 5148 12035 5151
rect 14182 5148 14188 5160
rect 12023 5120 14044 5148
rect 14143 5120 14188 5148
rect 12023 5117 12035 5120
rect 11977 5111 12035 5117
rect 2746 5052 4384 5080
rect 2866 4972 2872 5024
rect 2924 5012 2930 5024
rect 2961 5015 3019 5021
rect 2961 5012 2973 5015
rect 2924 4984 2973 5012
rect 2924 4972 2930 4984
rect 2961 4981 2973 4984
rect 3007 4981 3019 5015
rect 4356 5012 4384 5052
rect 5534 5040 5540 5092
rect 5592 5080 5598 5092
rect 5997 5083 6055 5089
rect 5997 5080 6009 5083
rect 5592 5052 6009 5080
rect 5592 5040 5598 5052
rect 5997 5049 6009 5052
rect 6043 5080 6055 5083
rect 6822 5080 6828 5092
rect 6043 5052 6828 5080
rect 6043 5049 6055 5052
rect 5997 5043 6055 5049
rect 6822 5040 6828 5052
rect 6880 5040 6886 5092
rect 8864 5052 9536 5080
rect 5902 5012 5908 5024
rect 4356 4984 5908 5012
rect 2961 4975 3019 4981
rect 5902 4972 5908 4984
rect 5960 4972 5966 5024
rect 6641 5015 6699 5021
rect 6641 4981 6653 5015
rect 6687 5012 6699 5015
rect 8864 5012 8892 5052
rect 6687 4984 8892 5012
rect 8941 5015 8999 5021
rect 6687 4981 6699 4984
rect 6641 4975 6699 4981
rect 8941 4981 8953 5015
rect 8987 5012 8999 5015
rect 9122 5012 9128 5024
rect 8987 4984 9128 5012
rect 8987 4981 8999 4984
rect 8941 4975 8999 4981
rect 9122 4972 9128 4984
rect 9180 4972 9186 5024
rect 9508 5012 9536 5052
rect 13814 5012 13820 5024
rect 9508 4984 13820 5012
rect 13814 4972 13820 4984
rect 13872 4972 13878 5024
rect 14016 5012 14044 5120
rect 14182 5108 14188 5120
rect 14240 5108 14246 5160
rect 14458 5148 14464 5160
rect 14419 5120 14464 5148
rect 14458 5108 14464 5120
rect 14516 5108 14522 5160
rect 14550 5108 14556 5160
rect 14608 5148 14614 5160
rect 14608 5120 15516 5148
rect 14608 5108 14614 5120
rect 15488 5080 15516 5120
rect 15654 5108 15660 5160
rect 15712 5148 15718 5160
rect 16114 5148 16120 5160
rect 15712 5120 16120 5148
rect 15712 5108 15718 5120
rect 16114 5108 16120 5120
rect 16172 5108 16178 5160
rect 16942 5148 16948 5160
rect 16903 5120 16948 5148
rect 16942 5108 16948 5120
rect 17000 5108 17006 5160
rect 18432 5148 18460 5188
rect 18874 5176 18880 5188
rect 18932 5176 18938 5228
rect 19426 5176 19432 5228
rect 19484 5216 19490 5228
rect 22480 5225 22508 5256
rect 22554 5244 22560 5296
rect 22612 5284 22618 5296
rect 23293 5287 23351 5293
rect 23293 5284 23305 5287
rect 22612 5256 23305 5284
rect 22612 5244 22618 5256
rect 23293 5253 23305 5256
rect 23339 5253 23351 5287
rect 23293 5247 23351 5253
rect 19521 5219 19579 5225
rect 19521 5216 19533 5219
rect 19484 5188 19533 5216
rect 19484 5176 19490 5188
rect 19521 5185 19533 5188
rect 19567 5185 19579 5219
rect 19521 5179 19579 5185
rect 22465 5219 22523 5225
rect 22465 5185 22477 5219
rect 22511 5185 22523 5219
rect 22465 5179 22523 5185
rect 24578 5176 24584 5228
rect 24636 5216 24642 5228
rect 24673 5219 24731 5225
rect 24673 5216 24685 5219
rect 24636 5188 24685 5216
rect 24636 5176 24642 5188
rect 24673 5185 24685 5188
rect 24719 5185 24731 5219
rect 25332 5216 25360 5324
rect 28537 5321 28549 5324
rect 28583 5321 28595 5355
rect 28537 5315 28595 5321
rect 25685 5287 25743 5293
rect 25685 5253 25697 5287
rect 25731 5284 25743 5287
rect 28166 5284 28172 5296
rect 25731 5256 28172 5284
rect 25731 5253 25743 5256
rect 25685 5247 25743 5253
rect 28166 5244 28172 5256
rect 28224 5244 28230 5296
rect 28626 5244 28632 5296
rect 28684 5284 28690 5296
rect 28684 5256 29776 5284
rect 28684 5244 28690 5256
rect 24673 5179 24731 5185
rect 25240 5188 25360 5216
rect 17052 5120 18460 5148
rect 18693 5151 18751 5157
rect 17052 5080 17080 5120
rect 18693 5117 18705 5151
rect 18739 5148 18751 5151
rect 19334 5148 19340 5160
rect 18739 5120 19340 5148
rect 18739 5117 18751 5120
rect 18693 5111 18751 5117
rect 19334 5108 19340 5120
rect 19392 5108 19398 5160
rect 19797 5151 19855 5157
rect 19797 5117 19809 5151
rect 19843 5148 19855 5151
rect 21266 5148 21272 5160
rect 19843 5120 21272 5148
rect 19843 5117 19855 5120
rect 19797 5111 19855 5117
rect 21266 5108 21272 5120
rect 21324 5148 21330 5160
rect 22922 5148 22928 5160
rect 21324 5120 22928 5148
rect 21324 5108 21330 5120
rect 22922 5108 22928 5120
rect 22980 5108 22986 5160
rect 23198 5148 23204 5160
rect 23159 5120 23204 5148
rect 23198 5108 23204 5120
rect 23256 5108 23262 5160
rect 24026 5148 24032 5160
rect 23987 5120 24032 5148
rect 24026 5108 24032 5120
rect 24084 5108 24090 5160
rect 19518 5080 19524 5092
rect 15488 5052 17080 5080
rect 18248 5052 19524 5080
rect 16298 5012 16304 5024
rect 14016 4984 16304 5012
rect 16298 4972 16304 4984
rect 16356 5012 16362 5024
rect 18248 5012 18276 5052
rect 19518 5040 19524 5052
rect 19576 5040 19582 5092
rect 21910 5080 21916 5092
rect 20824 5052 21916 5080
rect 16356 4984 18276 5012
rect 16356 4972 16362 4984
rect 18782 4972 18788 5024
rect 18840 5012 18846 5024
rect 20824 5012 20852 5052
rect 21910 5040 21916 5052
rect 21968 5040 21974 5092
rect 22002 5040 22008 5092
rect 22060 5080 22066 5092
rect 25240 5080 25268 5188
rect 26786 5176 26792 5228
rect 26844 5216 26850 5228
rect 27157 5219 27215 5225
rect 27157 5216 27169 5219
rect 26844 5188 27169 5216
rect 26844 5176 26850 5188
rect 27157 5185 27169 5188
rect 27203 5185 27215 5219
rect 27157 5179 27215 5185
rect 27801 5219 27859 5225
rect 27801 5185 27813 5219
rect 27847 5216 27859 5219
rect 27847 5188 28304 5216
rect 27847 5185 27859 5188
rect 27801 5179 27859 5185
rect 25593 5151 25651 5157
rect 25593 5117 25605 5151
rect 25639 5117 25651 5151
rect 25593 5111 25651 5117
rect 22060 5052 25268 5080
rect 25608 5080 25636 5111
rect 25682 5108 25688 5160
rect 25740 5148 25746 5160
rect 25869 5151 25927 5157
rect 25869 5148 25881 5151
rect 25740 5120 25881 5148
rect 25740 5108 25746 5120
rect 25869 5117 25881 5120
rect 25915 5117 25927 5151
rect 28276 5148 28304 5188
rect 28350 5176 28356 5228
rect 28408 5216 28414 5228
rect 28445 5219 28503 5225
rect 28445 5216 28457 5219
rect 28408 5188 28457 5216
rect 28408 5176 28414 5188
rect 28445 5185 28457 5188
rect 28491 5216 28503 5219
rect 28994 5216 29000 5228
rect 28491 5188 29000 5216
rect 28491 5185 28503 5188
rect 28445 5179 28503 5185
rect 28994 5176 29000 5188
rect 29052 5176 29058 5228
rect 29089 5219 29147 5225
rect 29089 5185 29101 5219
rect 29135 5216 29147 5219
rect 29178 5216 29184 5228
rect 29135 5188 29184 5216
rect 29135 5185 29147 5188
rect 29089 5179 29147 5185
rect 29178 5176 29184 5188
rect 29236 5176 29242 5228
rect 29748 5225 29776 5256
rect 29733 5219 29791 5225
rect 29733 5185 29745 5219
rect 29779 5185 29791 5219
rect 30374 5216 30380 5228
rect 30335 5188 30380 5216
rect 29733 5179 29791 5185
rect 30374 5176 30380 5188
rect 30432 5176 30438 5228
rect 32950 5148 32956 5160
rect 25869 5111 25927 5117
rect 25976 5120 27936 5148
rect 28276 5120 32956 5148
rect 25976 5080 26004 5120
rect 27908 5089 27936 5120
rect 32950 5108 32956 5120
rect 33008 5108 33014 5160
rect 25608 5052 26004 5080
rect 27893 5083 27951 5089
rect 22060 5040 22066 5052
rect 27893 5049 27905 5083
rect 27939 5049 27951 5083
rect 27893 5043 27951 5049
rect 28258 5040 28264 5092
rect 28316 5080 28322 5092
rect 30006 5080 30012 5092
rect 28316 5052 30012 5080
rect 28316 5040 28322 5052
rect 30006 5040 30012 5052
rect 30064 5040 30070 5092
rect 18840 4984 20852 5012
rect 18840 4972 18846 4984
rect 20898 4972 20904 5024
rect 20956 5012 20962 5024
rect 21269 5015 21327 5021
rect 21269 5012 21281 5015
rect 20956 4984 21281 5012
rect 20956 4972 20962 4984
rect 21269 4981 21281 4984
rect 21315 5012 21327 5015
rect 22370 5012 22376 5024
rect 21315 4984 22376 5012
rect 21315 4981 21327 4984
rect 21269 4975 21327 4981
rect 22370 4972 22376 4984
rect 22428 4972 22434 5024
rect 22557 5015 22615 5021
rect 22557 4981 22569 5015
rect 22603 5012 22615 5015
rect 23290 5012 23296 5024
rect 22603 4984 23296 5012
rect 22603 4981 22615 4984
rect 22557 4975 22615 4981
rect 23290 4972 23296 4984
rect 23348 4972 23354 5024
rect 23382 4972 23388 5024
rect 23440 5012 23446 5024
rect 24765 5015 24823 5021
rect 24765 5012 24777 5015
rect 23440 4984 24777 5012
rect 23440 4972 23446 4984
rect 24765 4981 24777 4984
rect 24811 4981 24823 5015
rect 24765 4975 24823 4981
rect 26786 4972 26792 5024
rect 26844 5012 26850 5024
rect 27249 5015 27307 5021
rect 27249 5012 27261 5015
rect 26844 4984 27261 5012
rect 26844 4972 26850 4984
rect 27249 4981 27261 4984
rect 27295 4981 27307 5015
rect 27249 4975 27307 4981
rect 27522 4972 27528 5024
rect 27580 5012 27586 5024
rect 29181 5015 29239 5021
rect 29181 5012 29193 5015
rect 27580 4984 29193 5012
rect 27580 4972 27586 4984
rect 29181 4981 29193 4984
rect 29227 4981 29239 5015
rect 29181 4975 29239 4981
rect 29270 4972 29276 5024
rect 29328 5012 29334 5024
rect 29825 5015 29883 5021
rect 29825 5012 29837 5015
rect 29328 4984 29837 5012
rect 29328 4972 29334 4984
rect 29825 4981 29837 4984
rect 29871 4981 29883 5015
rect 29825 4975 29883 4981
rect 30469 5015 30527 5021
rect 30469 4981 30481 5015
rect 30515 5012 30527 5015
rect 30558 5012 30564 5024
rect 30515 4984 30564 5012
rect 30515 4981 30527 4984
rect 30469 4975 30527 4981
rect 30558 4972 30564 4984
rect 30616 4972 30622 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 7558 4808 7564 4820
rect 4632 4780 7564 4808
rect 3786 4740 3792 4752
rect 2608 4712 3792 4740
rect 1578 4604 1584 4616
rect 1539 4576 1584 4604
rect 1578 4564 1584 4576
rect 1636 4564 1642 4616
rect 2608 4613 2636 4712
rect 3786 4700 3792 4712
rect 3844 4700 3850 4752
rect 2685 4675 2743 4681
rect 2685 4641 2697 4675
rect 2731 4672 2743 4675
rect 4632 4672 4660 4780
rect 7558 4768 7564 4780
rect 7616 4768 7622 4820
rect 8294 4768 8300 4820
rect 8352 4808 8358 4820
rect 9950 4808 9956 4820
rect 8352 4780 9956 4808
rect 8352 4768 8358 4780
rect 9950 4768 9956 4780
rect 10008 4768 10014 4820
rect 10502 4768 10508 4820
rect 10560 4808 10566 4820
rect 18782 4808 18788 4820
rect 10560 4780 18788 4808
rect 10560 4768 10566 4780
rect 18782 4768 18788 4780
rect 18840 4768 18846 4820
rect 19784 4811 19842 4817
rect 19784 4777 19796 4811
rect 19830 4808 19842 4811
rect 19830 4780 21864 4808
rect 19830 4777 19842 4780
rect 19784 4771 19842 4777
rect 5902 4700 5908 4752
rect 5960 4740 5966 4752
rect 6273 4743 6331 4749
rect 6273 4740 6285 4743
rect 5960 4712 6285 4740
rect 5960 4700 5966 4712
rect 6273 4709 6285 4712
rect 6319 4740 6331 4743
rect 6319 4712 6868 4740
rect 6319 4709 6331 4712
rect 6273 4703 6331 4709
rect 2731 4644 4660 4672
rect 4801 4675 4859 4681
rect 2731 4641 2743 4644
rect 2685 4635 2743 4641
rect 4801 4641 4813 4675
rect 4847 4672 4859 4675
rect 4890 4672 4896 4684
rect 4847 4644 4896 4672
rect 4847 4641 4859 4644
rect 4801 4635 4859 4641
rect 4890 4632 4896 4644
rect 4948 4632 4954 4684
rect 6730 4672 6736 4684
rect 6691 4644 6736 4672
rect 6730 4632 6736 4644
rect 6788 4632 6794 4684
rect 6840 4672 6868 4712
rect 8202 4700 8208 4752
rect 8260 4740 8266 4752
rect 9490 4740 9496 4752
rect 8260 4712 9496 4740
rect 8260 4700 8266 4712
rect 9490 4700 9496 4712
rect 9548 4700 9554 4752
rect 11333 4743 11391 4749
rect 11333 4709 11345 4743
rect 11379 4740 11391 4743
rect 14458 4740 14464 4752
rect 11379 4712 11928 4740
rect 11379 4709 11391 4712
rect 11333 4703 11391 4709
rect 7009 4675 7067 4681
rect 7009 4672 7021 4675
rect 6840 4644 7021 4672
rect 7009 4641 7021 4644
rect 7055 4641 7067 4675
rect 7009 4635 7067 4641
rect 7374 4632 7380 4684
rect 7432 4672 7438 4684
rect 9582 4672 9588 4684
rect 7432 4644 9588 4672
rect 7432 4632 7438 4644
rect 9582 4632 9588 4644
rect 9640 4632 9646 4684
rect 9861 4675 9919 4681
rect 9861 4641 9873 4675
rect 9907 4672 9919 4675
rect 11146 4672 11152 4684
rect 9907 4644 11152 4672
rect 9907 4641 9919 4644
rect 9861 4635 9919 4641
rect 11146 4632 11152 4644
rect 11204 4632 11210 4684
rect 11790 4672 11796 4684
rect 11751 4644 11796 4672
rect 11790 4632 11796 4644
rect 11848 4632 11854 4684
rect 11900 4672 11928 4712
rect 13096 4712 14464 4740
rect 13096 4672 13124 4712
rect 14458 4700 14464 4712
rect 14516 4700 14522 4752
rect 16298 4740 16304 4752
rect 16259 4712 16304 4740
rect 16298 4700 16304 4712
rect 16356 4700 16362 4752
rect 21266 4740 21272 4752
rect 21227 4712 21272 4740
rect 21266 4700 21272 4712
rect 21324 4700 21330 4752
rect 11900 4644 13124 4672
rect 13262 4632 13268 4684
rect 13320 4672 13326 4684
rect 17310 4672 17316 4684
rect 13320 4644 17316 4672
rect 13320 4632 13326 4644
rect 17310 4632 17316 4644
rect 17368 4632 17374 4684
rect 18785 4675 18843 4681
rect 18785 4641 18797 4675
rect 18831 4672 18843 4675
rect 19242 4672 19248 4684
rect 18831 4644 19248 4672
rect 18831 4641 18843 4644
rect 18785 4635 18843 4641
rect 19242 4632 19248 4644
rect 19300 4632 19306 4684
rect 19521 4675 19579 4681
rect 19521 4641 19533 4675
rect 19567 4672 19579 4675
rect 21836 4672 21864 4780
rect 22002 4768 22008 4820
rect 22060 4808 22066 4820
rect 22060 4780 29776 4808
rect 22060 4768 22066 4780
rect 25682 4700 25688 4752
rect 25740 4740 25746 4752
rect 26694 4740 26700 4752
rect 25740 4712 26700 4740
rect 25740 4700 25746 4712
rect 26694 4700 26700 4712
rect 26752 4700 26758 4752
rect 26878 4700 26884 4752
rect 26936 4740 26942 4752
rect 26936 4712 27016 4740
rect 26936 4700 26942 4712
rect 24118 4672 24124 4684
rect 19567 4644 21772 4672
rect 21836 4644 24124 4672
rect 19567 4641 19579 4644
rect 19521 4635 19579 4641
rect 2593 4607 2651 4613
rect 2593 4573 2605 4607
rect 2639 4573 2651 4607
rect 3234 4604 3240 4616
rect 3195 4576 3240 4604
rect 2593 4567 2651 4573
rect 3234 4564 3240 4576
rect 3292 4564 3298 4616
rect 4522 4604 4528 4616
rect 4483 4576 4528 4604
rect 4522 4564 4528 4576
rect 4580 4564 4586 4616
rect 14274 4564 14280 4616
rect 14332 4604 14338 4616
rect 14553 4607 14611 4613
rect 14553 4604 14565 4607
rect 14332 4576 14565 4604
rect 14332 4564 14338 4576
rect 14553 4573 14565 4576
rect 14599 4573 14611 4607
rect 14553 4567 14611 4573
rect 16942 4564 16948 4616
rect 17000 4604 17006 4616
rect 17037 4607 17095 4613
rect 17037 4604 17049 4607
rect 17000 4576 17049 4604
rect 17000 4564 17006 4576
rect 17037 4573 17049 4576
rect 17083 4573 17095 4607
rect 17037 4567 17095 4573
rect 19150 4564 19156 4616
rect 19208 4604 19214 4616
rect 19536 4604 19564 4635
rect 21744 4616 21772 4644
rect 24118 4632 24124 4644
rect 24176 4632 24182 4684
rect 24946 4672 24952 4684
rect 24907 4644 24952 4672
rect 24946 4632 24952 4644
rect 25004 4632 25010 4684
rect 25774 4672 25780 4684
rect 25735 4644 25780 4672
rect 25774 4632 25780 4644
rect 25832 4632 25838 4684
rect 26234 4632 26240 4684
rect 26292 4672 26298 4684
rect 26786 4672 26792 4684
rect 26292 4644 26792 4672
rect 26292 4632 26298 4644
rect 26786 4632 26792 4644
rect 26844 4632 26850 4684
rect 26988 4681 27016 4712
rect 28810 4700 28816 4752
rect 28868 4740 28874 4752
rect 28868 4712 28913 4740
rect 28868 4700 28874 4712
rect 26973 4675 27031 4681
rect 26973 4641 26985 4675
rect 27019 4641 27031 4675
rect 26973 4635 27031 4641
rect 27798 4632 27804 4684
rect 27856 4672 27862 4684
rect 29270 4672 29276 4684
rect 27856 4644 29276 4672
rect 27856 4632 27862 4644
rect 29270 4632 29276 4644
rect 29328 4632 29334 4684
rect 21726 4604 21732 4616
rect 19208 4576 19564 4604
rect 21687 4576 21732 4604
rect 19208 4564 19214 4576
rect 21726 4564 21732 4576
rect 21784 4564 21790 4616
rect 26418 4564 26424 4616
rect 26476 4564 26482 4616
rect 28077 4607 28135 4613
rect 28077 4573 28089 4607
rect 28123 4604 28135 4607
rect 28166 4604 28172 4616
rect 28123 4576 28172 4604
rect 28123 4573 28135 4576
rect 28077 4567 28135 4573
rect 28166 4564 28172 4576
rect 28224 4564 28230 4616
rect 28350 4564 28356 4616
rect 28408 4604 28414 4616
rect 29748 4613 29776 4780
rect 30006 4768 30012 4820
rect 30064 4808 30070 4820
rect 30469 4811 30527 4817
rect 30469 4808 30481 4811
rect 30064 4780 30481 4808
rect 30064 4768 30070 4780
rect 30469 4777 30481 4780
rect 30515 4777 30527 4811
rect 31754 4808 31760 4820
rect 31715 4780 31760 4808
rect 30469 4771 30527 4777
rect 31754 4768 31760 4780
rect 31812 4768 31818 4820
rect 37826 4768 37832 4820
rect 37884 4808 37890 4820
rect 38197 4811 38255 4817
rect 38197 4808 38209 4811
rect 37884 4780 38209 4808
rect 37884 4768 37890 4780
rect 38197 4777 38209 4780
rect 38243 4777 38255 4811
rect 38197 4771 38255 4777
rect 29840 4712 32352 4740
rect 28721 4607 28779 4613
rect 28721 4604 28733 4607
rect 28408 4576 28733 4604
rect 28408 4564 28414 4576
rect 28721 4573 28733 4576
rect 28767 4573 28779 4607
rect 28721 4567 28779 4573
rect 29733 4607 29791 4613
rect 29733 4573 29745 4607
rect 29779 4573 29791 4607
rect 29733 4567 29791 4573
rect 5810 4496 5816 4548
rect 5868 4496 5874 4548
rect 6196 4508 6868 4536
rect 1762 4468 1768 4480
rect 1723 4440 1768 4468
rect 1762 4428 1768 4440
rect 1820 4428 1826 4480
rect 3329 4471 3387 4477
rect 3329 4437 3341 4471
rect 3375 4468 3387 4471
rect 6196 4468 6224 4508
rect 3375 4440 6224 4468
rect 6840 4468 6868 4508
rect 6914 4496 6920 4548
rect 6972 4536 6978 4548
rect 6972 4508 7498 4536
rect 8312 4508 8616 4536
rect 6972 4496 6978 4508
rect 8312 4468 8340 4508
rect 6840 4440 8340 4468
rect 3375 4437 3387 4440
rect 3329 4431 3387 4437
rect 8386 4428 8392 4480
rect 8444 4468 8450 4480
rect 8481 4471 8539 4477
rect 8481 4468 8493 4471
rect 8444 4440 8493 4468
rect 8444 4428 8450 4440
rect 8481 4437 8493 4440
rect 8527 4437 8539 4471
rect 8588 4468 8616 4508
rect 9968 4508 10350 4536
rect 9968 4468 9996 4508
rect 11790 4496 11796 4548
rect 11848 4536 11854 4548
rect 12066 4536 12072 4548
rect 11848 4508 12072 4536
rect 11848 4496 11854 4508
rect 12066 4496 12072 4508
rect 12124 4496 12130 4548
rect 12176 4508 12558 4536
rect 13372 4508 14780 4536
rect 8588 4440 9996 4468
rect 8481 4431 8539 4437
rect 10042 4428 10048 4480
rect 10100 4468 10106 4480
rect 12176 4468 12204 4508
rect 10100 4440 12204 4468
rect 10100 4428 10106 4440
rect 12250 4428 12256 4480
rect 12308 4468 12314 4480
rect 13372 4468 13400 4508
rect 13538 4468 13544 4480
rect 12308 4440 13400 4468
rect 13499 4440 13544 4468
rect 12308 4428 12314 4440
rect 13538 4428 13544 4440
rect 13596 4428 13602 4480
rect 14752 4468 14780 4508
rect 14826 4496 14832 4548
rect 14884 4536 14890 4548
rect 14884 4508 14929 4536
rect 14884 4496 14890 4508
rect 15102 4496 15108 4548
rect 15160 4536 15166 4548
rect 17218 4536 17224 4548
rect 15160 4508 15318 4536
rect 16500 4508 17224 4536
rect 15160 4496 15166 4508
rect 16500 4468 16528 4508
rect 17218 4496 17224 4508
rect 17276 4496 17282 4548
rect 17313 4539 17371 4545
rect 17313 4505 17325 4539
rect 17359 4505 17371 4539
rect 21174 4536 21180 4548
rect 18538 4508 20208 4536
rect 21022 4508 21180 4536
rect 17313 4499 17371 4505
rect 14752 4440 16528 4468
rect 16574 4428 16580 4480
rect 16632 4468 16638 4480
rect 17328 4468 17356 4499
rect 18690 4468 18696 4480
rect 16632 4440 18696 4468
rect 16632 4428 16638 4440
rect 18690 4428 18696 4440
rect 18748 4428 18754 4480
rect 18874 4428 18880 4480
rect 18932 4468 18938 4480
rect 19978 4468 19984 4480
rect 18932 4440 19984 4468
rect 18932 4428 18938 4440
rect 19978 4428 19984 4440
rect 20036 4428 20042 4480
rect 20180 4468 20208 4508
rect 21174 4496 21180 4508
rect 21232 4496 21238 4548
rect 21542 4496 21548 4548
rect 21600 4536 21606 4548
rect 22005 4539 22063 4545
rect 22005 4536 22017 4539
rect 21600 4508 22017 4536
rect 21600 4496 21606 4508
rect 22005 4505 22017 4508
rect 22051 4505 22063 4539
rect 24762 4536 24768 4548
rect 23230 4508 24768 4536
rect 22005 4499 22063 4505
rect 24762 4496 24768 4508
rect 24820 4496 24826 4548
rect 25034 4539 25092 4545
rect 25034 4505 25046 4539
rect 25080 4536 25092 4539
rect 25498 4536 25504 4548
rect 25080 4508 25504 4536
rect 25080 4505 25092 4508
rect 25034 4499 25092 4505
rect 25498 4496 25504 4508
rect 25556 4496 25562 4548
rect 26436 4536 26464 4564
rect 26605 4539 26663 4545
rect 26605 4536 26617 4539
rect 26436 4508 26617 4536
rect 26605 4505 26617 4508
rect 26651 4505 26663 4539
rect 26605 4499 26663 4505
rect 26697 4539 26755 4545
rect 26697 4505 26709 4539
rect 26743 4536 26755 4539
rect 27798 4536 27804 4548
rect 26743 4508 27804 4536
rect 26743 4505 26755 4508
rect 26697 4499 26755 4505
rect 27798 4496 27804 4508
rect 27856 4496 27862 4548
rect 28258 4496 28264 4548
rect 28316 4536 28322 4548
rect 29840 4536 29868 4712
rect 30374 4604 30380 4616
rect 30335 4576 30380 4604
rect 30374 4564 30380 4576
rect 30432 4564 30438 4616
rect 31205 4607 31263 4613
rect 31205 4573 31217 4607
rect 31251 4573 31263 4607
rect 31662 4604 31668 4616
rect 31623 4576 31668 4604
rect 31205 4567 31263 4573
rect 28316 4508 29868 4536
rect 31220 4536 31248 4567
rect 31662 4564 31668 4576
rect 31720 4564 31726 4616
rect 32324 4613 32352 4712
rect 32309 4607 32367 4613
rect 32309 4573 32321 4607
rect 32355 4573 32367 4607
rect 32309 4567 32367 4573
rect 33505 4607 33563 4613
rect 33505 4573 33517 4607
rect 33551 4604 33563 4607
rect 34698 4604 34704 4616
rect 33551 4576 34704 4604
rect 33551 4573 33563 4576
rect 33505 4567 33563 4573
rect 34698 4564 34704 4576
rect 34756 4564 34762 4616
rect 33042 4536 33048 4548
rect 31220 4508 33048 4536
rect 28316 4496 28322 4508
rect 33042 4496 33048 4508
rect 33100 4496 33106 4548
rect 38102 4536 38108 4548
rect 38063 4508 38108 4536
rect 38102 4496 38108 4508
rect 38160 4496 38166 4548
rect 20714 4468 20720 4480
rect 20180 4440 20720 4468
rect 20714 4428 20720 4440
rect 20772 4428 20778 4480
rect 20806 4428 20812 4480
rect 20864 4468 20870 4480
rect 21910 4468 21916 4480
rect 20864 4440 21916 4468
rect 20864 4428 20870 4440
rect 21910 4428 21916 4440
rect 21968 4428 21974 4480
rect 22278 4428 22284 4480
rect 22336 4468 22342 4480
rect 23477 4471 23535 4477
rect 23477 4468 23489 4471
rect 22336 4440 23489 4468
rect 22336 4428 22342 4440
rect 23477 4437 23489 4440
rect 23523 4437 23535 4471
rect 23477 4431 23535 4437
rect 26234 4428 26240 4480
rect 26292 4468 26298 4480
rect 28169 4471 28227 4477
rect 28169 4468 28181 4471
rect 26292 4440 28181 4468
rect 26292 4428 26298 4440
rect 28169 4437 28181 4440
rect 28215 4437 28227 4471
rect 28169 4431 28227 4437
rect 28902 4428 28908 4480
rect 28960 4468 28966 4480
rect 29825 4471 29883 4477
rect 29825 4468 29837 4471
rect 28960 4440 29837 4468
rect 28960 4428 28966 4440
rect 29825 4437 29837 4440
rect 29871 4437 29883 4471
rect 31018 4468 31024 4480
rect 30979 4440 31024 4468
rect 29825 4431 29883 4437
rect 31018 4428 31024 4440
rect 31076 4428 31082 4480
rect 32401 4471 32459 4477
rect 32401 4437 32413 4471
rect 32447 4468 32459 4471
rect 33502 4468 33508 4480
rect 32447 4440 33508 4468
rect 32447 4437 32459 4440
rect 32401 4431 32459 4437
rect 33502 4428 33508 4440
rect 33560 4428 33566 4480
rect 33594 4428 33600 4480
rect 33652 4468 33658 4480
rect 33652 4440 33697 4468
rect 33652 4428 33658 4440
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 4062 4224 4068 4276
rect 4120 4264 4126 4276
rect 8018 4264 8024 4276
rect 4120 4236 8024 4264
rect 4120 4224 4126 4236
rect 8018 4224 8024 4236
rect 8076 4224 8082 4276
rect 8110 4224 8116 4276
rect 8168 4264 8174 4276
rect 12250 4264 12256 4276
rect 8168 4236 12256 4264
rect 8168 4224 8174 4236
rect 12250 4224 12256 4236
rect 12308 4224 12314 4276
rect 12618 4264 12624 4276
rect 12406 4236 12624 4264
rect 3234 4196 3240 4208
rect 2056 4168 3240 4196
rect 2056 4137 2084 4168
rect 3234 4156 3240 4168
rect 3292 4156 3298 4208
rect 3694 4196 3700 4208
rect 3344 4168 3700 4196
rect 3344 4137 3372 4168
rect 3694 4156 3700 4168
rect 3752 4156 3758 4208
rect 3988 4168 4844 4196
rect 2041 4131 2099 4137
rect 2041 4097 2053 4131
rect 2087 4097 2099 4131
rect 2041 4091 2099 4097
rect 2685 4131 2743 4137
rect 2685 4097 2697 4131
rect 2731 4128 2743 4131
rect 3329 4131 3387 4137
rect 2731 4100 2820 4128
rect 2731 4097 2743 4100
rect 2685 4091 2743 4097
rect 2133 4063 2191 4069
rect 2133 4029 2145 4063
rect 2179 4029 2191 4063
rect 2792 4060 2820 4100
rect 3329 4097 3341 4131
rect 3375 4097 3387 4131
rect 3329 4091 3387 4097
rect 3510 4088 3516 4140
rect 3568 4128 3574 4140
rect 3988 4128 4016 4168
rect 4154 4128 4160 4140
rect 3568 4100 4016 4128
rect 4115 4100 4160 4128
rect 3568 4088 3574 4100
rect 4154 4088 4160 4100
rect 4212 4088 4218 4140
rect 4617 4131 4675 4137
rect 4617 4128 4629 4131
rect 4264 4100 4629 4128
rect 3234 4060 3240 4072
rect 2792 4032 3240 4060
rect 2133 4023 2191 4029
rect 2148 3992 2176 4023
rect 3234 4020 3240 4032
rect 3292 4060 3298 4072
rect 4264 4060 4292 4100
rect 4617 4097 4629 4100
rect 4663 4128 4675 4131
rect 4706 4128 4712 4140
rect 4663 4100 4712 4128
rect 4663 4097 4675 4100
rect 4617 4091 4675 4097
rect 4706 4088 4712 4100
rect 4764 4088 4770 4140
rect 4816 4128 4844 4168
rect 5810 4156 5816 4208
rect 5868 4196 5874 4208
rect 6454 4196 6460 4208
rect 5868 4168 6460 4196
rect 5868 4156 5874 4168
rect 6454 4156 6460 4168
rect 6512 4156 6518 4208
rect 7926 4156 7932 4208
rect 7984 4156 7990 4208
rect 9861 4199 9919 4205
rect 8680 4168 9812 4196
rect 5261 4131 5319 4137
rect 5261 4128 5273 4131
rect 4816 4100 5273 4128
rect 5261 4097 5273 4100
rect 5307 4097 5319 4131
rect 7098 4128 7104 4140
rect 7059 4100 7104 4128
rect 5261 4091 5319 4097
rect 7098 4088 7104 4100
rect 7156 4088 7162 4140
rect 7006 4060 7012 4072
rect 3292 4032 4292 4060
rect 4632 4032 7012 4060
rect 3292 4020 3298 4032
rect 4632 3992 4660 4032
rect 7006 4020 7012 4032
rect 7064 4020 7070 4072
rect 7377 4063 7435 4069
rect 7377 4029 7389 4063
rect 7423 4060 7435 4063
rect 7926 4060 7932 4072
rect 7423 4032 7932 4060
rect 7423 4029 7435 4032
rect 7377 4023 7435 4029
rect 7926 4020 7932 4032
rect 7984 4020 7990 4072
rect 8018 4020 8024 4072
rect 8076 4060 8082 4072
rect 8680 4060 8708 4168
rect 9122 4128 9128 4140
rect 9083 4100 9128 4128
rect 9122 4088 9128 4100
rect 9180 4088 9186 4140
rect 9784 4128 9812 4168
rect 9861 4165 9873 4199
rect 9907 4196 9919 4199
rect 10134 4196 10140 4208
rect 9907 4168 10140 4196
rect 9907 4165 9919 4168
rect 9861 4159 9919 4165
rect 10134 4156 10140 4168
rect 10192 4156 10198 4208
rect 12406 4196 12434 4236
rect 12618 4224 12624 4236
rect 12676 4224 12682 4276
rect 13262 4224 13268 4276
rect 13320 4264 13326 4276
rect 13320 4236 16988 4264
rect 13320 4224 13326 4236
rect 10244 4168 12434 4196
rect 10244 4128 10272 4168
rect 12526 4156 12532 4208
rect 12584 4196 12590 4208
rect 16960 4205 16988 4236
rect 17310 4224 17316 4276
rect 17368 4264 17374 4276
rect 22738 4264 22744 4276
rect 17368 4236 22744 4264
rect 17368 4224 17374 4236
rect 22738 4224 22744 4236
rect 22796 4224 22802 4276
rect 24762 4264 24768 4276
rect 23124 4236 24768 4264
rect 16945 4199 17003 4205
rect 12584 4168 12742 4196
rect 13556 4168 15318 4196
rect 12584 4156 12590 4168
rect 9784 4100 10272 4128
rect 11698 4088 11704 4140
rect 11756 4128 11762 4140
rect 11977 4131 12035 4137
rect 11977 4128 11989 4131
rect 11756 4100 11989 4128
rect 11756 4088 11762 4100
rect 11977 4097 11989 4100
rect 12023 4097 12035 4131
rect 11977 4091 12035 4097
rect 8076 4032 8708 4060
rect 8956 4032 10003 4060
rect 8076 4020 8082 4032
rect 2148 3964 4660 3992
rect 4709 3995 4767 4001
rect 4709 3961 4721 3995
rect 4755 3992 4767 3995
rect 4755 3964 7236 3992
rect 4755 3961 4767 3964
rect 4709 3955 4767 3961
rect 2777 3927 2835 3933
rect 2777 3893 2789 3927
rect 2823 3924 2835 3927
rect 2958 3924 2964 3936
rect 2823 3896 2964 3924
rect 2823 3893 2835 3896
rect 2777 3887 2835 3893
rect 2958 3884 2964 3896
rect 3016 3884 3022 3936
rect 3421 3927 3479 3933
rect 3421 3893 3433 3927
rect 3467 3924 3479 3927
rect 3786 3924 3792 3936
rect 3467 3896 3792 3924
rect 3467 3893 3479 3896
rect 3421 3887 3479 3893
rect 3786 3884 3792 3896
rect 3844 3884 3850 3936
rect 3973 3927 4031 3933
rect 3973 3893 3985 3927
rect 4019 3924 4031 3927
rect 5074 3924 5080 3936
rect 4019 3896 5080 3924
rect 4019 3893 4031 3896
rect 3973 3887 4031 3893
rect 5074 3884 5080 3896
rect 5132 3884 5138 3936
rect 5166 3884 5172 3936
rect 5224 3924 5230 3936
rect 5445 3927 5503 3933
rect 5445 3924 5457 3927
rect 5224 3896 5457 3924
rect 5224 3884 5230 3896
rect 5445 3893 5457 3896
rect 5491 3893 5503 3927
rect 7208 3924 7236 3964
rect 8386 3952 8392 4004
rect 8444 3992 8450 4004
rect 8956 3992 8984 4032
rect 8444 3964 8984 3992
rect 8444 3952 8450 3964
rect 9214 3952 9220 4004
rect 9272 3992 9278 4004
rect 9674 3992 9680 4004
rect 9272 3964 9680 3992
rect 9272 3952 9278 3964
rect 9674 3952 9680 3964
rect 9732 3952 9738 4004
rect 9975 3992 10003 4032
rect 10042 4020 10048 4072
rect 10100 4060 10106 4072
rect 10597 4063 10655 4069
rect 10597 4060 10609 4063
rect 10100 4032 10609 4060
rect 10100 4020 10106 4032
rect 10597 4029 10609 4032
rect 10643 4029 10655 4063
rect 10597 4023 10655 4029
rect 11054 4020 11060 4072
rect 11112 4060 11118 4072
rect 12253 4063 12311 4069
rect 12253 4060 12265 4063
rect 11112 4032 12265 4060
rect 11112 4020 11118 4032
rect 12253 4029 12265 4032
rect 12299 4029 12311 4063
rect 12253 4023 12311 4029
rect 12618 4020 12624 4072
rect 12676 4060 12682 4072
rect 13556 4060 13584 4168
rect 16945 4165 16957 4199
rect 16991 4165 17003 4199
rect 16945 4159 17003 4165
rect 17218 4156 17224 4208
rect 17276 4196 17282 4208
rect 18874 4196 18880 4208
rect 17276 4168 18880 4196
rect 17276 4156 17282 4168
rect 18874 4156 18880 4168
rect 18932 4156 18938 4208
rect 23124 4196 23152 4236
rect 24762 4224 24768 4236
rect 24820 4224 24826 4276
rect 25774 4224 25780 4276
rect 25832 4264 25838 4276
rect 26878 4264 26884 4276
rect 25832 4236 26884 4264
rect 25832 4224 25838 4236
rect 26878 4224 26884 4236
rect 26936 4224 26942 4276
rect 26970 4224 26976 4276
rect 27028 4264 27034 4276
rect 27028 4236 28672 4264
rect 27028 4224 27034 4236
rect 23290 4196 23296 4208
rect 19826 4168 23152 4196
rect 23251 4168 23296 4196
rect 23290 4156 23296 4168
rect 23348 4156 23354 4208
rect 24857 4199 24915 4205
rect 24857 4165 24869 4199
rect 24903 4196 24915 4199
rect 25038 4196 25044 4208
rect 24903 4168 25044 4196
rect 24903 4165 24915 4168
rect 24857 4159 24915 4165
rect 25038 4156 25044 4168
rect 25096 4156 25102 4208
rect 26062 4199 26120 4205
rect 26062 4165 26074 4199
rect 26108 4196 26120 4199
rect 27522 4196 27528 4208
rect 26108 4168 27528 4196
rect 26108 4165 26120 4168
rect 26062 4159 26120 4165
rect 27522 4156 27528 4168
rect 27580 4156 27586 4208
rect 27982 4156 27988 4208
rect 28040 4196 28046 4208
rect 28537 4199 28595 4205
rect 28537 4196 28549 4199
rect 28040 4168 28549 4196
rect 28040 4156 28046 4168
rect 28537 4165 28549 4168
rect 28583 4165 28595 4199
rect 28644 4196 28672 4236
rect 28994 4224 29000 4276
rect 29052 4264 29058 4276
rect 30650 4264 30656 4276
rect 29052 4236 30656 4264
rect 29052 4224 29058 4236
rect 30650 4224 30656 4236
rect 30708 4224 30714 4276
rect 33594 4196 33600 4208
rect 28644 4168 33600 4196
rect 28537 4159 28595 4165
rect 33594 4156 33600 4168
rect 33652 4156 33658 4208
rect 18046 4128 18052 4140
rect 16224 4100 18052 4128
rect 12676 4032 13584 4060
rect 12676 4020 12682 4032
rect 14274 4020 14280 4072
rect 14332 4060 14338 4072
rect 14553 4063 14611 4069
rect 14553 4060 14565 4063
rect 14332 4032 14565 4060
rect 14332 4020 14338 4032
rect 14553 4029 14565 4032
rect 14599 4029 14611 4063
rect 14553 4023 14611 4029
rect 14829 4063 14887 4069
rect 14829 4029 14841 4063
rect 14875 4060 14887 4063
rect 16224 4060 16252 4100
rect 18046 4088 18052 4100
rect 18104 4088 18110 4140
rect 20530 4088 20536 4140
rect 20588 4128 20594 4140
rect 20625 4131 20683 4137
rect 20625 4128 20637 4131
rect 20588 4100 20637 4128
rect 20588 4088 20594 4100
rect 20625 4097 20637 4100
rect 20671 4097 20683 4131
rect 20625 4091 20683 4097
rect 20714 4088 20720 4140
rect 20772 4128 20778 4140
rect 20772 4100 20817 4128
rect 20772 4088 20778 4100
rect 21082 4088 21088 4140
rect 21140 4128 21146 4140
rect 21269 4131 21327 4137
rect 21269 4128 21281 4131
rect 21140 4100 21281 4128
rect 21140 4088 21146 4100
rect 21269 4097 21281 4100
rect 21315 4097 21327 4131
rect 21269 4091 21327 4097
rect 21358 4088 21364 4140
rect 21416 4128 21422 4140
rect 21416 4100 21461 4128
rect 21416 4088 21422 4100
rect 21910 4088 21916 4140
rect 21968 4128 21974 4140
rect 22465 4131 22523 4137
rect 22465 4128 22477 4131
rect 21968 4100 22477 4128
rect 21968 4088 21974 4100
rect 22465 4097 22477 4100
rect 22511 4097 22523 4131
rect 22465 4091 22523 4097
rect 22554 4088 22560 4140
rect 22612 4128 22618 4140
rect 27154 4128 27160 4140
rect 22612 4100 22657 4128
rect 27115 4100 27160 4128
rect 22612 4088 22618 4100
rect 27154 4088 27160 4100
rect 27212 4088 27218 4140
rect 27801 4131 27859 4137
rect 27801 4097 27813 4131
rect 27847 4128 27859 4131
rect 27890 4128 27896 4140
rect 27847 4100 27896 4128
rect 27847 4097 27859 4100
rect 27801 4091 27859 4097
rect 27890 4088 27896 4100
rect 27948 4088 27954 4140
rect 28166 4088 28172 4140
rect 28224 4128 28230 4140
rect 28350 4128 28356 4140
rect 28224 4100 28356 4128
rect 28224 4088 28230 4100
rect 28350 4088 28356 4100
rect 28408 4128 28414 4140
rect 28445 4131 28503 4137
rect 28445 4128 28457 4131
rect 28408 4100 28457 4128
rect 28408 4088 28414 4100
rect 28445 4097 28457 4100
rect 28491 4097 28503 4131
rect 28445 4091 28503 4097
rect 28994 4088 29000 4140
rect 29052 4128 29058 4140
rect 29089 4131 29147 4137
rect 29089 4128 29101 4131
rect 29052 4100 29101 4128
rect 29052 4088 29058 4100
rect 29089 4097 29101 4100
rect 29135 4097 29147 4131
rect 29730 4128 29736 4140
rect 29691 4100 29736 4128
rect 29089 4091 29147 4097
rect 29730 4088 29736 4100
rect 29788 4088 29794 4140
rect 30006 4088 30012 4140
rect 30064 4128 30070 4140
rect 30377 4131 30435 4137
rect 30377 4128 30389 4131
rect 30064 4100 30389 4128
rect 30064 4088 30070 4100
rect 30377 4097 30389 4100
rect 30423 4097 30435 4131
rect 30377 4091 30435 4097
rect 30466 4088 30472 4140
rect 30524 4128 30530 4140
rect 30524 4100 30569 4128
rect 30524 4088 30530 4100
rect 30650 4088 30656 4140
rect 30708 4128 30714 4140
rect 31021 4131 31079 4137
rect 31021 4128 31033 4131
rect 30708 4100 31033 4128
rect 30708 4088 30714 4100
rect 31021 4097 31033 4100
rect 31067 4128 31079 4131
rect 31570 4128 31576 4140
rect 31067 4100 31576 4128
rect 31067 4097 31079 4100
rect 31021 4091 31079 4097
rect 31570 4088 31576 4100
rect 31628 4088 31634 4140
rect 32490 4128 32496 4140
rect 32451 4100 32496 4128
rect 32490 4088 32496 4100
rect 32548 4088 32554 4140
rect 33502 4088 33508 4140
rect 33560 4128 33566 4140
rect 33873 4131 33931 4137
rect 33873 4128 33885 4131
rect 33560 4100 33885 4128
rect 33560 4088 33566 4100
rect 33873 4097 33885 4100
rect 33919 4097 33931 4131
rect 33873 4091 33931 4097
rect 14875 4032 16252 4060
rect 16301 4063 16359 4069
rect 14875 4029 14887 4032
rect 14829 4023 14887 4029
rect 16301 4029 16313 4063
rect 16347 4060 16359 4063
rect 16574 4060 16580 4072
rect 16347 4032 16580 4060
rect 16347 4029 16359 4032
rect 16301 4023 16359 4029
rect 16574 4020 16580 4032
rect 16632 4020 16638 4072
rect 16942 4020 16948 4072
rect 17000 4060 17006 4072
rect 17681 4063 17739 4069
rect 17681 4060 17693 4063
rect 17000 4032 17693 4060
rect 17000 4020 17006 4032
rect 17681 4029 17693 4032
rect 17727 4060 17739 4063
rect 18325 4063 18383 4069
rect 18325 4060 18337 4063
rect 17727 4032 18337 4060
rect 17727 4029 17739 4032
rect 17681 4023 17739 4029
rect 11330 3992 11336 4004
rect 9975 3964 11336 3992
rect 11330 3952 11336 3964
rect 11388 3952 11394 4004
rect 13354 3924 13360 3936
rect 7208 3896 13360 3924
rect 5445 3887 5503 3893
rect 13354 3884 13360 3896
rect 13412 3884 13418 3936
rect 13446 3884 13452 3936
rect 13504 3924 13510 3936
rect 13725 3927 13783 3933
rect 13725 3924 13737 3927
rect 13504 3896 13737 3924
rect 13504 3884 13510 3896
rect 13725 3893 13737 3896
rect 13771 3893 13783 3927
rect 13725 3887 13783 3893
rect 14550 3884 14556 3936
rect 14608 3924 14614 3936
rect 16758 3924 16764 3936
rect 14608 3896 16764 3924
rect 14608 3884 14614 3896
rect 16758 3884 16764 3896
rect 16816 3884 16822 3936
rect 18156 3924 18184 4032
rect 18325 4029 18337 4032
rect 18371 4029 18383 4063
rect 18601 4063 18659 4069
rect 18601 4060 18613 4063
rect 18325 4023 18383 4029
rect 18432 4032 18613 4060
rect 18230 3952 18236 4004
rect 18288 3992 18294 4004
rect 18432 3992 18460 4032
rect 18601 4029 18613 4032
rect 18647 4029 18659 4063
rect 18601 4023 18659 4029
rect 18690 4020 18696 4072
rect 18748 4060 18754 4072
rect 20806 4060 20812 4072
rect 18748 4032 20812 4060
rect 18748 4020 18754 4032
rect 20806 4020 20812 4032
rect 20864 4020 20870 4072
rect 23198 4060 23204 4072
rect 23159 4032 23204 4060
rect 23198 4020 23204 4032
rect 23256 4020 23262 4072
rect 24118 4060 24124 4072
rect 24079 4032 24124 4060
rect 24118 4020 24124 4032
rect 24176 4020 24182 4072
rect 24394 4020 24400 4072
rect 24452 4060 24458 4072
rect 24765 4063 24823 4069
rect 24765 4060 24777 4063
rect 24452 4032 24777 4060
rect 24452 4020 24458 4032
rect 24765 4029 24777 4032
rect 24811 4029 24823 4063
rect 24765 4023 24823 4029
rect 24854 4020 24860 4072
rect 24912 4060 24918 4072
rect 25041 4063 25099 4069
rect 25041 4060 25053 4063
rect 24912 4032 25053 4060
rect 24912 4020 24918 4032
rect 25041 4029 25053 4032
rect 25087 4060 25099 4063
rect 25961 4063 26019 4069
rect 25961 4060 25973 4063
rect 25087 4032 25973 4060
rect 25087 4029 25099 4032
rect 25041 4023 25099 4029
rect 25961 4029 25973 4032
rect 26007 4029 26019 4063
rect 25961 4023 26019 4029
rect 26050 4020 26056 4072
rect 26108 4060 26114 4072
rect 27249 4063 27307 4069
rect 27249 4060 27261 4063
rect 26108 4032 27261 4060
rect 26108 4020 26114 4032
rect 27249 4029 27261 4032
rect 27295 4029 27307 4063
rect 27249 4023 27307 4029
rect 27614 4020 27620 4072
rect 27672 4060 27678 4072
rect 29181 4063 29239 4069
rect 29181 4060 29193 4063
rect 27672 4032 29193 4060
rect 27672 4020 27678 4032
rect 29181 4029 29193 4032
rect 29227 4029 29239 4063
rect 29181 4023 29239 4029
rect 18288 3964 18460 3992
rect 18288 3952 18294 3964
rect 21082 3952 21088 4004
rect 21140 3992 21146 4004
rect 23750 3992 23756 4004
rect 21140 3964 23756 3992
rect 21140 3952 21146 3964
rect 23750 3952 23756 3964
rect 23808 3992 23814 4004
rect 25590 3992 25596 4004
rect 23808 3964 25596 3992
rect 23808 3952 23814 3964
rect 25590 3952 25596 3964
rect 25648 3952 25654 4004
rect 26418 3952 26424 4004
rect 26476 3992 26482 4004
rect 26513 3995 26571 4001
rect 26513 3992 26525 3995
rect 26476 3964 26525 3992
rect 26476 3952 26482 3964
rect 26513 3961 26525 3964
rect 26559 3961 26571 3995
rect 29825 3995 29883 4001
rect 29825 3992 29837 3995
rect 26513 3955 26571 3961
rect 26620 3964 29837 3992
rect 19150 3924 19156 3936
rect 18156 3896 19156 3924
rect 19150 3884 19156 3896
rect 19208 3884 19214 3936
rect 19978 3884 19984 3936
rect 20036 3924 20042 3936
rect 20073 3927 20131 3933
rect 20073 3924 20085 3927
rect 20036 3896 20085 3924
rect 20036 3884 20042 3896
rect 20073 3893 20085 3896
rect 20119 3893 20131 3927
rect 20073 3887 20131 3893
rect 22646 3884 22652 3936
rect 22704 3924 22710 3936
rect 25314 3924 25320 3936
rect 22704 3896 25320 3924
rect 22704 3884 22710 3896
rect 25314 3884 25320 3896
rect 25372 3884 25378 3936
rect 25958 3884 25964 3936
rect 26016 3924 26022 3936
rect 26620 3924 26648 3964
rect 29825 3961 29837 3964
rect 29871 3961 29883 3995
rect 29825 3955 29883 3961
rect 30926 3952 30932 4004
rect 30984 3992 30990 4004
rect 33778 3992 33784 4004
rect 30984 3964 33784 3992
rect 30984 3952 30990 3964
rect 33778 3952 33784 3964
rect 33836 3952 33842 4004
rect 26016 3896 26648 3924
rect 26016 3884 26022 3896
rect 26786 3884 26792 3936
rect 26844 3924 26850 3936
rect 27893 3927 27951 3933
rect 27893 3924 27905 3927
rect 26844 3896 27905 3924
rect 26844 3884 26850 3896
rect 27893 3893 27905 3896
rect 27939 3893 27951 3927
rect 27893 3887 27951 3893
rect 27982 3884 27988 3936
rect 28040 3924 28046 3936
rect 30006 3924 30012 3936
rect 28040 3896 30012 3924
rect 28040 3884 28046 3896
rect 30006 3884 30012 3896
rect 30064 3884 30070 3936
rect 30282 3884 30288 3936
rect 30340 3924 30346 3936
rect 31113 3927 31171 3933
rect 31113 3924 31125 3927
rect 30340 3896 31125 3924
rect 30340 3884 30346 3896
rect 31113 3893 31125 3896
rect 31159 3893 31171 3927
rect 32306 3924 32312 3936
rect 32267 3896 32312 3924
rect 31113 3887 31171 3893
rect 32306 3884 32312 3896
rect 32364 3884 32370 3936
rect 33689 3927 33747 3933
rect 33689 3893 33701 3927
rect 33735 3924 33747 3927
rect 34790 3924 34796 3936
rect 33735 3896 34796 3924
rect 33735 3893 33747 3896
rect 33689 3887 33747 3893
rect 34790 3884 34796 3896
rect 34848 3884 34854 3936
rect 37182 3884 37188 3936
rect 37240 3924 37246 3936
rect 38289 3927 38347 3933
rect 38289 3924 38301 3927
rect 37240 3896 38301 3924
rect 37240 3884 37246 3896
rect 38289 3893 38301 3896
rect 38335 3893 38347 3927
rect 38289 3887 38347 3893
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 4062 3720 4068 3732
rect 4023 3692 4068 3720
rect 4062 3680 4068 3692
rect 4120 3680 4126 3732
rect 4522 3680 4528 3732
rect 4580 3720 4586 3732
rect 6914 3720 6920 3732
rect 4580 3692 6920 3720
rect 4580 3680 4586 3692
rect 6914 3680 6920 3692
rect 6972 3680 6978 3732
rect 7088 3723 7146 3729
rect 7088 3689 7100 3723
rect 7134 3720 7146 3723
rect 8573 3723 8631 3729
rect 7134 3692 8524 3720
rect 7134 3689 7146 3692
rect 7088 3683 7146 3689
rect 6365 3655 6423 3661
rect 3160 3624 4752 3652
rect 2222 3584 2228 3596
rect 2183 3556 2228 3584
rect 2222 3544 2228 3556
rect 2280 3544 2286 3596
rect 2685 3587 2743 3593
rect 2685 3553 2697 3587
rect 2731 3584 2743 3587
rect 3160 3584 3188 3624
rect 2731 3556 3188 3584
rect 2731 3553 2743 3556
rect 2685 3547 2743 3553
rect 4522 3544 4528 3596
rect 4580 3584 4586 3596
rect 4614 3584 4620 3596
rect 4580 3556 4620 3584
rect 4580 3544 4586 3556
rect 4614 3544 4620 3556
rect 4672 3544 4678 3596
rect 4724 3584 4752 3624
rect 6365 3621 6377 3655
rect 6411 3652 6423 3655
rect 6546 3652 6552 3664
rect 6411 3624 6552 3652
rect 6411 3621 6423 3624
rect 6365 3615 6423 3621
rect 6546 3612 6552 3624
rect 6604 3612 6610 3664
rect 8202 3612 8208 3664
rect 8260 3652 8266 3664
rect 8496 3652 8524 3692
rect 8573 3689 8585 3723
rect 8619 3720 8631 3723
rect 9490 3720 9496 3732
rect 8619 3692 9496 3720
rect 8619 3689 8631 3692
rect 8573 3683 8631 3689
rect 9490 3680 9496 3692
rect 9548 3680 9554 3732
rect 10302 3723 10360 3729
rect 10302 3720 10314 3723
rect 10152 3692 10314 3720
rect 9122 3652 9128 3664
rect 8260 3624 8432 3652
rect 8496 3624 9128 3652
rect 8260 3612 8266 3624
rect 6730 3584 6736 3596
rect 4724 3556 6736 3584
rect 6730 3544 6736 3556
rect 6788 3544 6794 3596
rect 6825 3587 6883 3593
rect 6825 3553 6837 3587
rect 6871 3584 6883 3587
rect 7190 3584 7196 3596
rect 6871 3556 7196 3584
rect 6871 3553 6883 3556
rect 6825 3547 6883 3553
rect 7190 3544 7196 3556
rect 7248 3544 7254 3596
rect 8404 3584 8432 3624
rect 9122 3612 9128 3624
rect 9180 3612 9186 3664
rect 9950 3612 9956 3664
rect 10008 3652 10014 3664
rect 10152 3652 10180 3692
rect 10302 3689 10314 3692
rect 10348 3689 10360 3723
rect 10302 3683 10360 3689
rect 10686 3680 10692 3732
rect 10744 3720 10750 3732
rect 11793 3723 11851 3729
rect 10744 3692 11376 3720
rect 10744 3680 10750 3692
rect 10008 3624 10180 3652
rect 11348 3652 11376 3692
rect 11793 3689 11805 3723
rect 11839 3720 11851 3723
rect 11882 3720 11888 3732
rect 11839 3692 11888 3720
rect 11839 3689 11851 3692
rect 11793 3683 11851 3689
rect 11882 3680 11888 3692
rect 11940 3680 11946 3732
rect 12894 3680 12900 3732
rect 12952 3720 12958 3732
rect 16022 3720 16028 3732
rect 12952 3692 15608 3720
rect 15983 3692 16028 3720
rect 12952 3680 12958 3692
rect 14182 3652 14188 3664
rect 11348 3624 14188 3652
rect 10008 3612 10014 3624
rect 14182 3612 14188 3624
rect 14240 3612 14246 3664
rect 15580 3652 15608 3692
rect 16022 3680 16028 3692
rect 16080 3680 16086 3732
rect 16485 3723 16543 3729
rect 16485 3689 16497 3723
rect 16531 3720 16543 3723
rect 22186 3720 22192 3732
rect 16531 3692 22192 3720
rect 16531 3689 16543 3692
rect 16485 3683 16543 3689
rect 22186 3680 22192 3692
rect 22244 3680 22250 3732
rect 23842 3720 23848 3732
rect 22480 3692 23428 3720
rect 23803 3692 23848 3720
rect 20898 3652 20904 3664
rect 15580 3624 17264 3652
rect 12526 3584 12532 3596
rect 8404 3556 12532 3584
rect 12526 3544 12532 3556
rect 12584 3544 12590 3596
rect 13262 3584 13268 3596
rect 12820 3556 13268 3584
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3516 1639 3519
rect 2240 3516 2268 3544
rect 2590 3516 2596 3528
rect 1627 3488 2268 3516
rect 2551 3488 2596 3516
rect 1627 3485 1639 3488
rect 1581 3479 1639 3485
rect 2590 3476 2596 3488
rect 2648 3476 2654 3528
rect 3237 3519 3295 3525
rect 3237 3485 3249 3519
rect 3283 3516 3295 3519
rect 3694 3516 3700 3528
rect 3283 3488 3700 3516
rect 3283 3485 3295 3488
rect 3237 3479 3295 3485
rect 3694 3476 3700 3488
rect 3752 3476 3758 3528
rect 3970 3516 3976 3528
rect 3931 3488 3976 3516
rect 3970 3476 3976 3488
rect 4028 3476 4034 3528
rect 9582 3476 9588 3528
rect 9640 3516 9646 3528
rect 10042 3516 10048 3528
rect 9640 3488 10048 3516
rect 9640 3476 9646 3488
rect 10042 3476 10048 3488
rect 10100 3476 10106 3528
rect 12820 3525 12848 3556
rect 13262 3544 13268 3556
rect 13320 3544 13326 3596
rect 16942 3544 16948 3596
rect 17000 3584 17006 3596
rect 17129 3587 17187 3593
rect 17129 3584 17141 3587
rect 17000 3556 17141 3584
rect 17000 3544 17006 3556
rect 17129 3553 17141 3556
rect 17175 3553 17187 3587
rect 17236 3584 17264 3624
rect 20732 3624 20904 3652
rect 18414 3584 18420 3596
rect 17236 3556 18420 3584
rect 17129 3547 17187 3553
rect 18414 3544 18420 3556
rect 18472 3544 18478 3596
rect 19150 3544 19156 3596
rect 19208 3584 19214 3596
rect 19429 3587 19487 3593
rect 19429 3584 19441 3587
rect 19208 3556 19441 3584
rect 19208 3544 19214 3556
rect 19429 3553 19441 3556
rect 19475 3553 19487 3587
rect 19429 3547 19487 3553
rect 19705 3587 19763 3593
rect 19705 3553 19717 3587
rect 19751 3584 19763 3587
rect 20732 3584 20760 3624
rect 20898 3612 20904 3624
rect 20956 3612 20962 3664
rect 22480 3584 22508 3692
rect 23400 3652 23428 3692
rect 23842 3680 23848 3692
rect 23900 3680 23906 3732
rect 24486 3680 24492 3732
rect 24544 3720 24550 3732
rect 24544 3692 27200 3720
rect 24544 3680 24550 3692
rect 26694 3652 26700 3664
rect 23400 3624 26700 3652
rect 26694 3612 26700 3624
rect 26752 3612 26758 3664
rect 22646 3584 22652 3596
rect 19751 3556 20760 3584
rect 20824 3556 22508 3584
rect 22607 3556 22652 3584
rect 19751 3553 19763 3556
rect 19705 3547 19763 3553
rect 12807 3519 12865 3525
rect 12807 3485 12819 3519
rect 12853 3485 12865 3519
rect 14274 3516 14280 3528
rect 14187 3488 14280 3516
rect 12807 3479 12865 3485
rect 14274 3476 14280 3488
rect 14332 3476 14338 3528
rect 16669 3519 16727 3525
rect 16669 3485 16681 3519
rect 16715 3485 16727 3519
rect 16669 3479 16727 3485
rect 3329 3451 3387 3457
rect 3329 3417 3341 3451
rect 3375 3448 3387 3451
rect 4798 3448 4804 3460
rect 3375 3420 4804 3448
rect 3375 3417 3387 3420
rect 3329 3411 3387 3417
rect 4798 3408 4804 3420
rect 4856 3408 4862 3460
rect 4893 3451 4951 3457
rect 4893 3417 4905 3451
rect 4939 3448 4951 3451
rect 4982 3448 4988 3460
rect 4939 3420 4988 3448
rect 4939 3417 4951 3420
rect 4893 3411 4951 3417
rect 4982 3408 4988 3420
rect 5040 3408 5046 3460
rect 5626 3408 5632 3460
rect 5684 3408 5690 3460
rect 6840 3420 7590 3448
rect 1762 3380 1768 3392
rect 1723 3352 1768 3380
rect 1762 3340 1768 3352
rect 1820 3340 1826 3392
rect 2958 3340 2964 3392
rect 3016 3380 3022 3392
rect 6840 3380 6868 3420
rect 8754 3408 8760 3460
rect 8812 3448 8818 3460
rect 9217 3451 9275 3457
rect 9217 3448 9229 3451
rect 8812 3420 9229 3448
rect 8812 3408 8818 3420
rect 9217 3417 9229 3420
rect 9263 3417 9275 3451
rect 9398 3448 9404 3460
rect 9359 3420 9404 3448
rect 9217 3411 9275 3417
rect 9398 3408 9404 3420
rect 9456 3408 9462 3460
rect 9858 3408 9864 3460
rect 9916 3448 9922 3460
rect 9916 3420 10810 3448
rect 9916 3408 9922 3420
rect 12618 3408 12624 3460
rect 12676 3448 12682 3460
rect 13170 3448 13176 3460
rect 12676 3420 13176 3448
rect 12676 3408 12682 3420
rect 13170 3408 13176 3420
rect 13228 3408 13234 3460
rect 13633 3451 13691 3457
rect 13633 3417 13645 3451
rect 13679 3448 13691 3451
rect 13906 3448 13912 3460
rect 13679 3420 13912 3448
rect 13679 3417 13691 3420
rect 13633 3411 13691 3417
rect 13906 3408 13912 3420
rect 13964 3448 13970 3460
rect 14292 3448 14320 3476
rect 13964 3420 14320 3448
rect 13964 3408 13970 3420
rect 14458 3408 14464 3460
rect 14516 3448 14522 3460
rect 14553 3451 14611 3457
rect 14553 3448 14565 3451
rect 14516 3420 14565 3448
rect 14516 3408 14522 3420
rect 14553 3417 14565 3420
rect 14599 3417 14611 3451
rect 14553 3411 14611 3417
rect 14660 3420 15042 3448
rect 3016 3352 6868 3380
rect 3016 3340 3022 3352
rect 6914 3340 6920 3392
rect 6972 3380 6978 3392
rect 12342 3380 12348 3392
rect 6972 3352 12348 3380
rect 6972 3340 6978 3352
rect 12342 3340 12348 3352
rect 12400 3340 12406 3392
rect 13354 3340 13360 3392
rect 13412 3380 13418 3392
rect 14660 3380 14688 3420
rect 13412 3352 14688 3380
rect 16684 3380 16712 3479
rect 18506 3476 18512 3528
rect 18564 3476 18570 3528
rect 20824 3502 20852 3556
rect 22646 3544 22652 3556
rect 22704 3544 22710 3596
rect 22738 3544 22744 3596
rect 22796 3584 22802 3596
rect 26786 3584 26792 3596
rect 22796 3556 26792 3584
rect 22796 3544 22802 3556
rect 26786 3544 26792 3556
rect 26844 3544 26850 3596
rect 27062 3584 27068 3596
rect 27023 3556 27068 3584
rect 27062 3544 27068 3556
rect 27120 3544 27126 3596
rect 27172 3584 27200 3692
rect 27522 3680 27528 3732
rect 27580 3720 27586 3732
rect 29270 3720 29276 3732
rect 27580 3692 29276 3720
rect 27580 3680 27586 3692
rect 29270 3680 29276 3692
rect 29328 3680 29334 3732
rect 29454 3680 29460 3732
rect 29512 3720 29518 3732
rect 30742 3720 30748 3732
rect 29512 3692 30748 3720
rect 29512 3680 29518 3692
rect 30742 3680 30748 3692
rect 30800 3680 30806 3732
rect 32950 3720 32956 3732
rect 31726 3692 32628 3720
rect 32911 3692 32956 3720
rect 27246 3612 27252 3664
rect 27304 3652 27310 3664
rect 29822 3652 29828 3664
rect 27304 3624 29828 3652
rect 27304 3612 27310 3624
rect 29822 3612 29828 3624
rect 29880 3612 29886 3664
rect 31726 3652 31754 3692
rect 29932 3624 31754 3652
rect 32600 3652 32628 3692
rect 32950 3680 32956 3692
rect 33008 3680 33014 3732
rect 33597 3655 33655 3661
rect 33597 3652 33609 3655
rect 32600 3624 33609 3652
rect 27172 3556 28212 3584
rect 21910 3516 21916 3528
rect 21823 3488 21916 3516
rect 21910 3476 21916 3488
rect 21968 3516 21974 3528
rect 22278 3516 22284 3528
rect 21968 3488 22284 3516
rect 21968 3476 21974 3488
rect 22278 3476 22284 3488
rect 22336 3476 22342 3528
rect 23290 3476 23296 3528
rect 23348 3516 23354 3528
rect 23750 3516 23756 3528
rect 23348 3488 23393 3516
rect 23711 3488 23756 3516
rect 23348 3476 23354 3488
rect 23750 3476 23756 3488
rect 23808 3476 23814 3528
rect 25314 3476 25320 3528
rect 25372 3516 25378 3528
rect 25372 3488 25417 3516
rect 25372 3476 25378 3488
rect 17402 3448 17408 3460
rect 17363 3420 17408 3448
rect 17402 3408 17408 3420
rect 17460 3408 17466 3460
rect 21450 3448 21456 3460
rect 21411 3420 21456 3448
rect 21450 3408 21456 3420
rect 21508 3408 21514 3460
rect 22738 3448 22744 3460
rect 22699 3420 22744 3448
rect 22738 3408 22744 3420
rect 22796 3408 22802 3460
rect 24670 3448 24676 3460
rect 24631 3420 24676 3448
rect 24670 3408 24676 3420
rect 24728 3408 24734 3460
rect 24765 3451 24823 3457
rect 24765 3417 24777 3451
rect 24811 3417 24823 3451
rect 25866 3448 25872 3460
rect 25827 3420 25872 3448
rect 24765 3411 24823 3417
rect 18782 3380 18788 3392
rect 16684 3352 18788 3380
rect 13412 3340 13418 3352
rect 18782 3340 18788 3352
rect 18840 3340 18846 3392
rect 18877 3383 18935 3389
rect 18877 3349 18889 3383
rect 18923 3380 18935 3383
rect 19334 3380 19340 3392
rect 18923 3352 19340 3380
rect 18923 3349 18935 3352
rect 18877 3343 18935 3349
rect 19334 3340 19340 3352
rect 19392 3340 19398 3392
rect 22005 3383 22063 3389
rect 22005 3349 22017 3383
rect 22051 3380 22063 3383
rect 24780 3380 24808 3411
rect 25866 3408 25872 3420
rect 25924 3408 25930 3460
rect 25958 3408 25964 3460
rect 26016 3448 26022 3460
rect 26016 3420 26061 3448
rect 26016 3408 26022 3420
rect 26234 3408 26240 3460
rect 26292 3448 26298 3460
rect 26513 3451 26571 3457
rect 26513 3448 26525 3451
rect 26292 3420 26525 3448
rect 26292 3408 26298 3420
rect 26513 3417 26525 3420
rect 26559 3448 26571 3451
rect 27062 3448 27068 3460
rect 26559 3420 27068 3448
rect 26559 3417 26571 3420
rect 26513 3411 26571 3417
rect 27062 3408 27068 3420
rect 27120 3408 27126 3460
rect 27157 3451 27215 3457
rect 27157 3417 27169 3451
rect 27203 3448 27215 3451
rect 27338 3448 27344 3460
rect 27203 3420 27344 3448
rect 27203 3417 27215 3420
rect 27157 3411 27215 3417
rect 27338 3408 27344 3420
rect 27396 3408 27402 3460
rect 28074 3448 28080 3460
rect 28035 3420 28080 3448
rect 28074 3408 28080 3420
rect 28132 3408 28138 3460
rect 28184 3448 28212 3556
rect 28442 3544 28448 3596
rect 28500 3584 28506 3596
rect 29932 3584 29960 3624
rect 33597 3621 33609 3624
rect 33643 3621 33655 3655
rect 33597 3615 33655 3621
rect 32306 3584 32312 3596
rect 28500 3556 29960 3584
rect 30392 3556 32312 3584
rect 28500 3544 28506 3556
rect 28350 3476 28356 3528
rect 28408 3516 28414 3528
rect 28537 3519 28595 3525
rect 28537 3516 28549 3519
rect 28408 3488 28549 3516
rect 28408 3476 28414 3488
rect 28537 3485 28549 3488
rect 28583 3516 28595 3519
rect 28810 3516 28816 3528
rect 28583 3488 28816 3516
rect 28583 3485 28595 3488
rect 28537 3479 28595 3485
rect 28810 3476 28816 3488
rect 28868 3476 28874 3528
rect 28994 3476 29000 3528
rect 29052 3516 29058 3528
rect 30392 3525 30420 3556
rect 32306 3544 32312 3556
rect 32364 3544 32370 3596
rect 29733 3519 29791 3525
rect 29733 3516 29745 3519
rect 29052 3488 29745 3516
rect 29052 3476 29058 3488
rect 29733 3485 29745 3488
rect 29779 3485 29791 3519
rect 29733 3479 29791 3485
rect 30377 3519 30435 3525
rect 30377 3485 30389 3519
rect 30423 3485 30435 3519
rect 30377 3479 30435 3485
rect 30742 3476 30748 3528
rect 30800 3516 30806 3528
rect 31021 3519 31079 3525
rect 31021 3516 31033 3519
rect 30800 3488 31033 3516
rect 30800 3476 30806 3488
rect 31021 3485 31033 3488
rect 31067 3516 31079 3519
rect 31294 3516 31300 3528
rect 31067 3488 31300 3516
rect 31067 3485 31079 3488
rect 31021 3479 31079 3485
rect 31294 3476 31300 3488
rect 31352 3476 31358 3528
rect 31849 3519 31907 3525
rect 31849 3485 31861 3519
rect 31895 3485 31907 3519
rect 31849 3479 31907 3485
rect 31864 3448 31892 3479
rect 31938 3476 31944 3528
rect 31996 3516 32002 3528
rect 33137 3519 33195 3525
rect 33137 3516 33149 3519
rect 31996 3488 33149 3516
rect 31996 3476 32002 3488
rect 33137 3485 33149 3488
rect 33183 3485 33195 3519
rect 33778 3516 33784 3528
rect 33739 3488 33784 3516
rect 33137 3479 33195 3485
rect 33778 3476 33784 3488
rect 33836 3476 33842 3528
rect 38010 3516 38016 3528
rect 37971 3488 38016 3516
rect 38010 3476 38016 3488
rect 38068 3476 38074 3528
rect 28184 3420 31892 3448
rect 22051 3352 24808 3380
rect 22051 3349 22063 3352
rect 22005 3343 22063 3349
rect 24854 3340 24860 3392
rect 24912 3380 24918 3392
rect 27982 3380 27988 3392
rect 24912 3352 27988 3380
rect 24912 3340 24918 3352
rect 27982 3340 27988 3352
rect 28040 3340 28046 3392
rect 28534 3340 28540 3392
rect 28592 3380 28598 3392
rect 28629 3383 28687 3389
rect 28629 3380 28641 3383
rect 28592 3352 28641 3380
rect 28592 3340 28598 3352
rect 28629 3349 28641 3352
rect 28675 3349 28687 3383
rect 28629 3343 28687 3349
rect 28810 3340 28816 3392
rect 28868 3380 28874 3392
rect 29454 3380 29460 3392
rect 28868 3352 29460 3380
rect 28868 3340 28874 3352
rect 29454 3340 29460 3352
rect 29512 3340 29518 3392
rect 29638 3340 29644 3392
rect 29696 3380 29702 3392
rect 29825 3383 29883 3389
rect 29825 3380 29837 3383
rect 29696 3352 29837 3380
rect 29696 3340 29702 3352
rect 29825 3349 29837 3352
rect 29871 3349 29883 3383
rect 30466 3380 30472 3392
rect 30427 3352 30472 3380
rect 29825 3343 29883 3349
rect 30466 3340 30472 3352
rect 30524 3340 30530 3392
rect 31110 3380 31116 3392
rect 31071 3352 31116 3380
rect 31110 3340 31116 3352
rect 31168 3340 31174 3392
rect 31478 3340 31484 3392
rect 31536 3380 31542 3392
rect 31665 3383 31723 3389
rect 31665 3380 31677 3383
rect 31536 3352 31677 3380
rect 31536 3340 31542 3352
rect 31665 3349 31677 3352
rect 31711 3349 31723 3383
rect 31665 3343 31723 3349
rect 31754 3340 31760 3392
rect 31812 3380 31818 3392
rect 32309 3383 32367 3389
rect 32309 3380 32321 3383
rect 31812 3352 32321 3380
rect 31812 3340 31818 3352
rect 32309 3349 32321 3352
rect 32355 3349 32367 3383
rect 38194 3380 38200 3392
rect 38155 3352 38200 3380
rect 32309 3343 32367 3349
rect 38194 3340 38200 3352
rect 38252 3340 38258 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 2774 3176 2780 3188
rect 1596 3148 2780 3176
rect 1596 3049 1624 3148
rect 2774 3136 2780 3148
rect 2832 3136 2838 3188
rect 3053 3179 3111 3185
rect 3053 3145 3065 3179
rect 3099 3176 3111 3179
rect 3142 3176 3148 3188
rect 3099 3148 3148 3176
rect 3099 3145 3111 3148
rect 3053 3139 3111 3145
rect 3142 3136 3148 3148
rect 3200 3136 3206 3188
rect 3786 3136 3792 3188
rect 3844 3176 3850 3188
rect 5534 3176 5540 3188
rect 3844 3148 5540 3176
rect 3844 3136 3850 3148
rect 5534 3136 5540 3148
rect 5592 3136 5598 3188
rect 5997 3179 6055 3185
rect 5997 3145 6009 3179
rect 6043 3176 6055 3179
rect 6362 3176 6368 3188
rect 6043 3148 6368 3176
rect 6043 3145 6055 3148
rect 5997 3139 6055 3145
rect 6362 3136 6368 3148
rect 6420 3136 6426 3188
rect 11882 3176 11888 3188
rect 6564 3148 11888 3176
rect 2406 3108 2412 3120
rect 2367 3080 2412 3108
rect 2406 3068 2412 3080
rect 2464 3068 2470 3120
rect 4614 3108 4620 3120
rect 4264 3080 4620 3108
rect 1581 3043 1639 3049
rect 1581 3009 1593 3043
rect 1627 3009 1639 3043
rect 1581 3003 1639 3009
rect 2317 3043 2375 3049
rect 2317 3009 2329 3043
rect 2363 3040 2375 3043
rect 2866 3040 2872 3052
rect 2363 3012 2872 3040
rect 2363 3009 2375 3012
rect 2317 3003 2375 3009
rect 2866 3000 2872 3012
rect 2924 3000 2930 3052
rect 2961 3043 3019 3049
rect 2961 3009 2973 3043
rect 3007 3040 3019 3043
rect 3234 3040 3240 3052
rect 3007 3012 3240 3040
rect 3007 3009 3019 3012
rect 2961 3003 3019 3009
rect 3234 3000 3240 3012
rect 3292 3000 3298 3052
rect 3786 3040 3792 3052
rect 3747 3012 3792 3040
rect 3786 3000 3792 3012
rect 3844 3000 3850 3052
rect 4264 3049 4292 3080
rect 4614 3068 4620 3080
rect 4672 3068 4678 3120
rect 4798 3068 4804 3120
rect 4856 3108 4862 3120
rect 4856 3080 5014 3108
rect 4856 3068 4862 3080
rect 6564 3049 6592 3148
rect 11882 3136 11888 3148
rect 11940 3136 11946 3188
rect 23198 3176 23204 3188
rect 12544 3148 23204 3176
rect 8110 3068 8116 3120
rect 8168 3108 8174 3120
rect 8168 3080 8213 3108
rect 8168 3068 8174 3080
rect 8570 3068 8576 3120
rect 8628 3068 8634 3120
rect 11146 3068 11152 3120
rect 11204 3108 11210 3120
rect 12544 3108 12572 3148
rect 23198 3136 23204 3148
rect 23256 3136 23262 3188
rect 23753 3179 23811 3185
rect 23753 3145 23765 3179
rect 23799 3176 23811 3179
rect 24026 3176 24032 3188
rect 23799 3148 24032 3176
rect 23799 3145 23811 3148
rect 23753 3139 23811 3145
rect 24026 3136 24032 3148
rect 24084 3136 24090 3188
rect 26234 3176 26240 3188
rect 24320 3148 26240 3176
rect 11204 3080 12572 3108
rect 12636 3080 13216 3108
rect 11204 3068 11210 3080
rect 4249 3043 4307 3049
rect 4249 3009 4261 3043
rect 4295 3009 4307 3043
rect 4249 3003 4307 3009
rect 6549 3043 6607 3049
rect 6549 3009 6561 3043
rect 6595 3009 6607 3043
rect 6549 3003 6607 3009
rect 7190 3000 7196 3052
rect 7248 3040 7254 3052
rect 7742 3040 7748 3052
rect 7248 3012 7748 3040
rect 7248 3000 7254 3012
rect 7742 3000 7748 3012
rect 7800 3040 7806 3052
rect 7837 3043 7895 3049
rect 7837 3040 7849 3043
rect 7800 3012 7849 3040
rect 7800 3000 7806 3012
rect 7837 3009 7849 3012
rect 7883 3009 7895 3043
rect 10226 3040 10232 3052
rect 7837 3003 7895 3009
rect 9646 3012 10232 3040
rect 4522 2972 4528 2984
rect 4483 2944 4528 2972
rect 4522 2932 4528 2944
rect 4580 2932 4586 2984
rect 5074 2932 5080 2984
rect 5132 2972 5138 2984
rect 9646 2972 9674 3012
rect 10226 3000 10232 3012
rect 10284 3000 10290 3052
rect 10321 3043 10379 3049
rect 10321 3009 10333 3043
rect 10367 3040 10379 3043
rect 10502 3040 10508 3052
rect 10367 3012 10508 3040
rect 10367 3009 10379 3012
rect 10321 3003 10379 3009
rect 10502 3000 10508 3012
rect 10560 3000 10566 3052
rect 10870 3000 10876 3052
rect 10928 3040 10934 3052
rect 10965 3043 11023 3049
rect 10965 3040 10977 3043
rect 10928 3012 10977 3040
rect 10928 3000 10934 3012
rect 10965 3009 10977 3012
rect 11011 3009 11023 3043
rect 10965 3003 11023 3009
rect 12161 3043 12219 3049
rect 12161 3009 12173 3043
rect 12207 3040 12219 3043
rect 12636 3040 12664 3080
rect 12207 3012 12664 3040
rect 12713 3043 12771 3049
rect 12207 3009 12219 3012
rect 12161 3003 12219 3009
rect 12713 3009 12725 3043
rect 12759 3009 12771 3043
rect 12894 3040 12900 3052
rect 12855 3012 12900 3040
rect 12713 3003 12771 3009
rect 5132 2944 9674 2972
rect 9861 2975 9919 2981
rect 5132 2932 5138 2944
rect 9861 2941 9873 2975
rect 9907 2941 9919 2975
rect 9861 2935 9919 2941
rect 10413 2975 10471 2981
rect 10413 2941 10425 2975
rect 10459 2972 10471 2975
rect 10594 2972 10600 2984
rect 10459 2944 10600 2972
rect 10459 2941 10471 2944
rect 10413 2935 10471 2941
rect 5920 2876 7972 2904
rect 658 2796 664 2848
rect 716 2836 722 2848
rect 1765 2839 1823 2845
rect 1765 2836 1777 2839
rect 716 2808 1777 2836
rect 716 2796 722 2808
rect 1765 2805 1777 2808
rect 1811 2805 1823 2839
rect 1765 2799 1823 2805
rect 3605 2839 3663 2845
rect 3605 2805 3617 2839
rect 3651 2836 3663 2839
rect 5920 2836 5948 2876
rect 3651 2808 5948 2836
rect 3651 2805 3663 2808
rect 3605 2799 3663 2805
rect 6454 2796 6460 2848
rect 6512 2836 6518 2848
rect 6733 2839 6791 2845
rect 6733 2836 6745 2839
rect 6512 2808 6745 2836
rect 6512 2796 6518 2808
rect 6733 2805 6745 2808
rect 6779 2805 6791 2839
rect 6733 2799 6791 2805
rect 7098 2796 7104 2848
rect 7156 2836 7162 2848
rect 7650 2836 7656 2848
rect 7156 2808 7656 2836
rect 7156 2796 7162 2808
rect 7650 2796 7656 2808
rect 7708 2796 7714 2848
rect 7944 2836 7972 2876
rect 9122 2864 9128 2916
rect 9180 2904 9186 2916
rect 9876 2904 9904 2935
rect 10594 2932 10600 2944
rect 10652 2932 10658 2984
rect 11057 2975 11115 2981
rect 11057 2941 11069 2975
rect 11103 2972 11115 2975
rect 11146 2972 11152 2984
rect 11103 2944 11152 2972
rect 11103 2941 11115 2944
rect 11057 2935 11115 2941
rect 11146 2932 11152 2944
rect 11204 2932 11210 2984
rect 11974 2904 11980 2916
rect 9180 2876 9904 2904
rect 10336 2876 11192 2904
rect 11935 2876 11980 2904
rect 9180 2864 9186 2876
rect 10336 2836 10364 2876
rect 7944 2808 10364 2836
rect 11164 2836 11192 2876
rect 11974 2864 11980 2876
rect 12032 2864 12038 2916
rect 12728 2904 12756 3003
rect 12894 3000 12900 3012
rect 12952 3000 12958 3052
rect 13188 2972 13216 3080
rect 13538 3068 13544 3120
rect 13596 3108 13602 3120
rect 13633 3111 13691 3117
rect 13633 3108 13645 3111
rect 13596 3080 13645 3108
rect 13596 3068 13602 3080
rect 13633 3077 13645 3080
rect 13679 3077 13691 3111
rect 15010 3108 15016 3120
rect 14858 3080 15016 3108
rect 13633 3071 13691 3077
rect 15010 3068 15016 3080
rect 15068 3068 15074 3120
rect 16298 3108 16304 3120
rect 16259 3080 16304 3108
rect 16298 3068 16304 3080
rect 16356 3068 16362 3120
rect 19058 3108 19064 3120
rect 18538 3080 19064 3108
rect 19058 3068 19064 3080
rect 19116 3068 19122 3120
rect 19150 3068 19156 3120
rect 19208 3068 19214 3120
rect 24320 3117 24348 3148
rect 26234 3136 26240 3148
rect 26292 3136 26298 3188
rect 27430 3136 27436 3188
rect 27488 3176 27494 3188
rect 32401 3179 32459 3185
rect 32401 3176 32413 3179
rect 27488 3148 32413 3176
rect 27488 3136 27494 3148
rect 32401 3145 32413 3148
rect 32447 3145 32459 3179
rect 33042 3176 33048 3188
rect 33003 3148 33048 3176
rect 32401 3139 32459 3145
rect 33042 3136 33048 3148
rect 33100 3136 33106 3188
rect 34698 3136 34704 3188
rect 34756 3176 34762 3188
rect 36725 3179 36783 3185
rect 36725 3176 36737 3179
rect 34756 3148 36737 3176
rect 34756 3136 34762 3148
rect 36725 3145 36737 3148
rect 36771 3145 36783 3179
rect 36725 3139 36783 3145
rect 24305 3111 24363 3117
rect 24305 3077 24317 3111
rect 24351 3077 24363 3111
rect 24305 3071 24363 3077
rect 24397 3111 24455 3117
rect 24397 3077 24409 3111
rect 24443 3108 24455 3111
rect 25961 3111 26019 3117
rect 24443 3080 25728 3108
rect 24443 3077 24455 3080
rect 24397 3071 24455 3077
rect 13262 3000 13268 3052
rect 13320 3040 13326 3052
rect 13357 3043 13415 3049
rect 13357 3040 13369 3043
rect 13320 3012 13369 3040
rect 13320 3000 13326 3012
rect 13357 3009 13369 3012
rect 13403 3009 13415 3043
rect 16114 3040 16120 3052
rect 16075 3012 16120 3040
rect 13357 3003 13415 3009
rect 16114 3000 16120 3012
rect 16172 3000 16178 3052
rect 16942 3000 16948 3052
rect 17000 3040 17006 3052
rect 17037 3043 17095 3049
rect 17037 3040 17049 3043
rect 17000 3012 17049 3040
rect 17000 3000 17006 3012
rect 17037 3009 17049 3012
rect 17083 3009 17095 3043
rect 17037 3003 17095 3009
rect 18966 3000 18972 3052
rect 19024 3040 19030 3052
rect 19168 3040 19196 3068
rect 19245 3043 19303 3049
rect 19245 3040 19257 3043
rect 19024 3012 19257 3040
rect 19024 3000 19030 3012
rect 19245 3009 19257 3012
rect 19291 3009 19303 3043
rect 19245 3003 19303 3009
rect 14826 2972 14832 2984
rect 13188 2944 14832 2972
rect 14826 2932 14832 2944
rect 14884 2932 14890 2984
rect 14918 2932 14924 2984
rect 14976 2972 14982 2984
rect 15105 2975 15163 2981
rect 15105 2972 15117 2975
rect 14976 2944 15117 2972
rect 14976 2932 14982 2944
rect 15105 2941 15117 2944
rect 15151 2941 15163 2975
rect 15105 2935 15163 2941
rect 17313 2975 17371 2981
rect 17313 2941 17325 2975
rect 17359 2972 17371 2975
rect 19150 2972 19156 2984
rect 17359 2944 19156 2972
rect 17359 2941 17371 2944
rect 17313 2935 17371 2941
rect 19150 2932 19156 2944
rect 19208 2932 19214 2984
rect 19518 2972 19524 2984
rect 19431 2944 19524 2972
rect 19518 2932 19524 2944
rect 19576 2972 19582 2984
rect 20530 2972 20536 2984
rect 19576 2944 20536 2972
rect 19576 2932 19582 2944
rect 20530 2932 20536 2944
rect 20588 2932 20594 2984
rect 20640 2904 20668 3026
rect 21726 3000 21732 3052
rect 21784 3040 21790 3052
rect 22005 3043 22063 3049
rect 22005 3040 22017 3043
rect 21784 3012 22017 3040
rect 21784 3000 21790 3012
rect 22005 3009 22017 3012
rect 22051 3009 22063 3043
rect 22005 3003 22063 3009
rect 23382 3000 23388 3052
rect 23440 3000 23446 3052
rect 20714 2932 20720 2984
rect 20772 2972 20778 2984
rect 22281 2975 22339 2981
rect 22281 2972 22293 2975
rect 20772 2944 22293 2972
rect 20772 2932 20778 2944
rect 22281 2941 22293 2944
rect 22327 2972 22339 2975
rect 24854 2972 24860 2984
rect 22327 2944 24860 2972
rect 22327 2941 22339 2944
rect 22281 2935 22339 2941
rect 24854 2932 24860 2944
rect 24912 2932 24918 2984
rect 25130 2972 25136 2984
rect 25091 2944 25136 2972
rect 25130 2932 25136 2944
rect 25188 2932 25194 2984
rect 24946 2904 24952 2916
rect 12728 2876 13492 2904
rect 20640 2876 22094 2904
rect 13354 2836 13360 2848
rect 11164 2808 13360 2836
rect 13354 2796 13360 2808
rect 13412 2796 13418 2848
rect 13464 2836 13492 2876
rect 14826 2836 14832 2848
rect 13464 2808 14832 2836
rect 14826 2796 14832 2808
rect 14884 2796 14890 2848
rect 17402 2796 17408 2848
rect 17460 2836 17466 2848
rect 18785 2839 18843 2845
rect 18785 2836 18797 2839
rect 17460 2808 18797 2836
rect 17460 2796 17466 2808
rect 18785 2805 18797 2808
rect 18831 2836 18843 2839
rect 20070 2836 20076 2848
rect 18831 2808 20076 2836
rect 18831 2805 18843 2808
rect 18785 2799 18843 2805
rect 20070 2796 20076 2808
rect 20128 2796 20134 2848
rect 20993 2839 21051 2845
rect 20993 2805 21005 2839
rect 21039 2836 21051 2839
rect 21818 2836 21824 2848
rect 21039 2808 21824 2836
rect 21039 2805 21051 2808
rect 20993 2799 21051 2805
rect 21818 2796 21824 2808
rect 21876 2796 21882 2848
rect 22066 2836 22094 2876
rect 23308 2876 24952 2904
rect 23308 2836 23336 2876
rect 24946 2864 24952 2876
rect 25004 2864 25010 2916
rect 22066 2808 23336 2836
rect 25700 2836 25728 3080
rect 25961 3077 25973 3111
rect 26007 3108 26019 3111
rect 26970 3108 26976 3120
rect 26007 3080 26976 3108
rect 26007 3077 26019 3080
rect 25961 3071 26019 3077
rect 26970 3068 26976 3080
rect 27028 3068 27034 3120
rect 27338 3117 27344 3120
rect 27334 3071 27344 3117
rect 27396 3108 27402 3120
rect 27396 3080 27434 3108
rect 27338 3068 27344 3071
rect 27396 3068 27402 3080
rect 27614 3068 27620 3120
rect 27672 3108 27678 3120
rect 27672 3080 29224 3108
rect 27672 3068 27678 3080
rect 28350 3040 28356 3052
rect 28311 3012 28356 3040
rect 28350 3000 28356 3012
rect 28408 3000 28414 3052
rect 28997 3043 29055 3049
rect 28997 3009 29009 3043
rect 29043 3040 29055 3043
rect 29086 3040 29092 3052
rect 29043 3012 29092 3040
rect 29043 3009 29055 3012
rect 28997 3003 29055 3009
rect 29086 3000 29092 3012
rect 29144 3000 29150 3052
rect 25869 2975 25927 2981
rect 25869 2941 25881 2975
rect 25915 2972 25927 2975
rect 26142 2972 26148 2984
rect 25915 2944 26148 2972
rect 25915 2941 25927 2944
rect 25869 2935 25927 2941
rect 26142 2932 26148 2944
rect 26200 2932 26206 2984
rect 27246 2972 27252 2984
rect 27207 2944 27252 2972
rect 27246 2932 27252 2944
rect 27304 2932 27310 2984
rect 27338 2932 27344 2984
rect 27396 2972 27402 2984
rect 27525 2975 27583 2981
rect 27525 2972 27537 2975
rect 27396 2944 27537 2972
rect 27396 2932 27402 2944
rect 27525 2941 27537 2944
rect 27571 2941 27583 2975
rect 28902 2972 28908 2984
rect 27525 2935 27583 2941
rect 27816 2944 28908 2972
rect 26418 2904 26424 2916
rect 26379 2876 26424 2904
rect 26418 2864 26424 2876
rect 26476 2864 26482 2916
rect 26970 2864 26976 2916
rect 27028 2904 27034 2916
rect 27816 2904 27844 2944
rect 28902 2932 28908 2944
rect 28960 2932 28966 2984
rect 29089 2907 29147 2913
rect 29089 2904 29101 2907
rect 27028 2876 27844 2904
rect 27908 2876 29101 2904
rect 27028 2864 27034 2876
rect 27908 2836 27936 2876
rect 29089 2873 29101 2876
rect 29135 2873 29147 2907
rect 29196 2904 29224 3080
rect 30374 3068 30380 3120
rect 30432 3108 30438 3120
rect 33689 3111 33747 3117
rect 33689 3108 33701 3111
rect 30432 3080 33701 3108
rect 30432 3068 30438 3080
rect 33689 3077 33701 3080
rect 33735 3077 33747 3111
rect 33689 3071 33747 3077
rect 29546 3000 29552 3052
rect 29604 3040 29610 3052
rect 29641 3043 29699 3049
rect 29641 3040 29653 3043
rect 29604 3012 29653 3040
rect 29604 3000 29610 3012
rect 29641 3009 29653 3012
rect 29687 3009 29699 3043
rect 29641 3003 29699 3009
rect 29656 2972 29684 3003
rect 29914 3000 29920 3052
rect 29972 3040 29978 3052
rect 30285 3043 30343 3049
rect 30285 3040 30297 3043
rect 29972 3012 30297 3040
rect 29972 3000 29978 3012
rect 30285 3009 30297 3012
rect 30331 3009 30343 3043
rect 30929 3043 30987 3049
rect 30929 3040 30941 3043
rect 30285 3003 30343 3009
rect 30392 3012 30941 3040
rect 30392 2972 30420 3012
rect 30929 3009 30941 3012
rect 30975 3009 30987 3043
rect 31570 3040 31576 3052
rect 31531 3012 31576 3040
rect 30929 3003 30987 3009
rect 31570 3000 31576 3012
rect 31628 3000 31634 3052
rect 31846 3000 31852 3052
rect 31904 3040 31910 3052
rect 32309 3043 32367 3049
rect 32309 3040 32321 3043
rect 31904 3012 32321 3040
rect 31904 3000 31910 3012
rect 32309 3009 32321 3012
rect 32355 3009 32367 3043
rect 32309 3003 32367 3009
rect 32398 3000 32404 3052
rect 32456 3040 32462 3052
rect 32953 3043 33011 3049
rect 32953 3040 32965 3043
rect 32456 3012 32965 3040
rect 32456 3000 32462 3012
rect 32953 3009 32965 3012
rect 32999 3009 33011 3043
rect 32953 3003 33011 3009
rect 33597 3043 33655 3049
rect 33597 3009 33609 3043
rect 33643 3009 33655 3043
rect 33597 3003 33655 3009
rect 29656 2944 30420 2972
rect 30650 2932 30656 2984
rect 30708 2972 30714 2984
rect 30708 2944 32076 2972
rect 30708 2932 30714 2944
rect 31938 2904 31944 2916
rect 29196 2876 31944 2904
rect 29089 2867 29147 2873
rect 31938 2864 31944 2876
rect 31996 2864 32002 2916
rect 32048 2904 32076 2944
rect 33612 2904 33640 3003
rect 35434 3000 35440 3052
rect 35492 3040 35498 3052
rect 35713 3043 35771 3049
rect 35713 3040 35725 3043
rect 35492 3012 35725 3040
rect 35492 3000 35498 3012
rect 35713 3009 35725 3012
rect 35759 3009 35771 3043
rect 35713 3003 35771 3009
rect 36909 3043 36967 3049
rect 36909 3009 36921 3043
rect 36955 3040 36967 3043
rect 37826 3040 37832 3052
rect 36955 3012 37832 3040
rect 36955 3009 36967 3012
rect 36909 3003 36967 3009
rect 37826 3000 37832 3012
rect 37884 3000 37890 3052
rect 37918 3000 37924 3052
rect 37976 3040 37982 3052
rect 38013 3043 38071 3049
rect 38013 3040 38025 3043
rect 37976 3012 38025 3040
rect 37976 3000 37982 3012
rect 38013 3009 38025 3012
rect 38059 3009 38071 3043
rect 38013 3003 38071 3009
rect 32048 2876 33640 2904
rect 34606 2864 34612 2916
rect 34664 2904 34670 2916
rect 35529 2907 35587 2913
rect 35529 2904 35541 2907
rect 34664 2876 35541 2904
rect 34664 2864 34670 2876
rect 35529 2873 35541 2876
rect 35575 2873 35587 2907
rect 35529 2867 35587 2873
rect 28442 2836 28448 2848
rect 25700 2808 27936 2836
rect 28403 2808 28448 2836
rect 28442 2796 28448 2808
rect 28500 2796 28506 2848
rect 29730 2836 29736 2848
rect 29691 2808 29736 2836
rect 29730 2796 29736 2808
rect 29788 2796 29794 2848
rect 30374 2836 30380 2848
rect 30335 2808 30380 2836
rect 30374 2796 30380 2808
rect 30432 2796 30438 2848
rect 30466 2796 30472 2848
rect 30524 2836 30530 2848
rect 31021 2839 31079 2845
rect 31021 2836 31033 2839
rect 30524 2808 31033 2836
rect 30524 2796 30530 2808
rect 31021 2805 31033 2808
rect 31067 2805 31079 2839
rect 31662 2836 31668 2848
rect 31623 2808 31668 2836
rect 31021 2799 31079 2805
rect 31662 2796 31668 2808
rect 31720 2796 31726 2848
rect 38197 2839 38255 2845
rect 38197 2805 38209 2839
rect 38243 2836 38255 2839
rect 38654 2836 38660 2848
rect 38243 2808 38660 2836
rect 38243 2805 38255 2808
rect 38197 2799 38255 2805
rect 38654 2796 38660 2808
rect 38712 2796 38718 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 4982 2592 4988 2644
rect 5040 2632 5046 2644
rect 5997 2635 6055 2641
rect 5997 2632 6009 2635
rect 5040 2604 6009 2632
rect 5040 2592 5046 2604
rect 5997 2601 6009 2604
rect 6043 2632 6055 2635
rect 7466 2632 7472 2644
rect 6043 2604 7472 2632
rect 6043 2601 6055 2604
rect 5997 2595 6055 2601
rect 7466 2592 7472 2604
rect 7524 2592 7530 2644
rect 13725 2635 13783 2641
rect 13725 2632 13737 2635
rect 11072 2604 13737 2632
rect 14 2524 20 2576
rect 72 2564 78 2576
rect 2593 2567 2651 2573
rect 2593 2564 2605 2567
rect 72 2536 2605 2564
rect 72 2524 78 2536
rect 2593 2533 2605 2536
rect 2639 2533 2651 2567
rect 2593 2527 2651 2533
rect 4249 2499 4307 2505
rect 4249 2465 4261 2499
rect 4295 2496 4307 2499
rect 4614 2496 4620 2508
rect 4295 2468 4620 2496
rect 4295 2465 4307 2468
rect 4249 2459 4307 2465
rect 4614 2456 4620 2468
rect 4672 2456 4678 2508
rect 6733 2499 6791 2505
rect 6733 2465 6745 2499
rect 6779 2496 6791 2499
rect 7006 2496 7012 2508
rect 6779 2468 7012 2496
rect 6779 2465 6791 2468
rect 6733 2459 6791 2465
rect 7006 2456 7012 2468
rect 7064 2456 7070 2508
rect 7742 2456 7748 2508
rect 7800 2496 7806 2508
rect 9401 2499 9459 2505
rect 9401 2496 9413 2499
rect 7800 2468 9413 2496
rect 7800 2456 7806 2468
rect 9401 2465 9413 2468
rect 9447 2465 9459 2499
rect 9401 2459 9459 2465
rect 9677 2499 9735 2505
rect 9677 2465 9689 2499
rect 9723 2496 9735 2499
rect 11072 2496 11100 2604
rect 13725 2601 13737 2604
rect 13771 2632 13783 2635
rect 18877 2635 18935 2641
rect 13771 2604 16574 2632
rect 13771 2601 13783 2604
rect 13725 2595 13783 2601
rect 16298 2564 16304 2576
rect 16259 2536 16304 2564
rect 16298 2524 16304 2536
rect 16356 2524 16362 2576
rect 9723 2468 11100 2496
rect 11977 2499 12035 2505
rect 9723 2465 9735 2468
rect 9677 2459 9735 2465
rect 11977 2465 11989 2499
rect 12023 2496 12035 2499
rect 13262 2496 13268 2508
rect 12023 2468 13268 2496
rect 12023 2465 12035 2468
rect 11977 2459 12035 2465
rect 13262 2456 13268 2468
rect 13320 2496 13326 2508
rect 13906 2496 13912 2508
rect 13320 2468 13912 2496
rect 13320 2456 13326 2468
rect 13906 2456 13912 2468
rect 13964 2496 13970 2508
rect 14553 2499 14611 2505
rect 14553 2496 14565 2499
rect 13964 2468 14565 2496
rect 13964 2456 13970 2468
rect 14553 2465 14565 2468
rect 14599 2465 14611 2499
rect 14553 2459 14611 2465
rect 14829 2499 14887 2505
rect 14829 2465 14841 2499
rect 14875 2496 14887 2499
rect 15470 2496 15476 2508
rect 14875 2468 15476 2496
rect 14875 2465 14887 2468
rect 14829 2459 14887 2465
rect 15470 2456 15476 2468
rect 15528 2456 15534 2508
rect 1670 2428 1676 2440
rect 1631 2400 1676 2428
rect 1670 2388 1676 2400
rect 1728 2388 1734 2440
rect 2409 2431 2467 2437
rect 2409 2397 2421 2431
rect 2455 2428 2467 2431
rect 2498 2428 2504 2440
rect 2455 2400 2504 2428
rect 2455 2397 2467 2400
rect 2409 2391 2467 2397
rect 2498 2388 2504 2400
rect 2556 2388 2562 2440
rect 3142 2428 3148 2440
rect 3103 2400 3148 2428
rect 3142 2388 3148 2400
rect 3200 2388 3206 2440
rect 4522 2360 4528 2372
rect 4483 2332 4528 2360
rect 4522 2320 4528 2332
rect 4580 2320 4586 2372
rect 5810 2360 5816 2372
rect 5750 2332 5816 2360
rect 5810 2320 5816 2332
rect 5868 2320 5874 2372
rect 6362 2320 6368 2372
rect 6420 2360 6426 2372
rect 7009 2363 7067 2369
rect 7009 2360 7021 2363
rect 6420 2332 7021 2360
rect 6420 2320 6426 2332
rect 7009 2329 7021 2332
rect 7055 2329 7067 2363
rect 7009 2323 7067 2329
rect 7466 2320 7472 2372
rect 7524 2320 7530 2372
rect 12250 2360 12256 2372
rect 8312 2332 10166 2360
rect 10980 2332 11284 2360
rect 12211 2332 12256 2360
rect 1857 2295 1915 2301
rect 1857 2261 1869 2295
rect 1903 2292 1915 2295
rect 1946 2292 1952 2304
rect 1903 2264 1952 2292
rect 1903 2261 1915 2264
rect 1857 2255 1915 2261
rect 1946 2252 1952 2264
rect 2004 2252 2010 2304
rect 3234 2252 3240 2304
rect 3292 2292 3298 2304
rect 3329 2295 3387 2301
rect 3329 2292 3341 2295
rect 3292 2264 3341 2292
rect 3292 2252 3298 2264
rect 3329 2261 3341 2264
rect 3375 2261 3387 2295
rect 3329 2255 3387 2261
rect 5534 2252 5540 2304
rect 5592 2292 5598 2304
rect 8312 2292 8340 2332
rect 8478 2292 8484 2304
rect 5592 2264 8340 2292
rect 8439 2264 8484 2292
rect 5592 2252 5598 2264
rect 8478 2252 8484 2264
rect 8536 2252 8542 2304
rect 9766 2252 9772 2304
rect 9824 2292 9830 2304
rect 10980 2292 11008 2332
rect 11146 2292 11152 2304
rect 9824 2264 11008 2292
rect 11107 2264 11152 2292
rect 9824 2252 9830 2264
rect 11146 2252 11152 2264
rect 11204 2252 11210 2304
rect 11256 2292 11284 2332
rect 12250 2320 12256 2332
rect 12308 2320 12314 2372
rect 12406 2332 12742 2360
rect 12406 2292 12434 2332
rect 15286 2320 15292 2372
rect 15344 2320 15350 2372
rect 11256 2264 12434 2292
rect 13630 2252 13636 2304
rect 13688 2292 13694 2304
rect 16206 2292 16212 2304
rect 13688 2264 16212 2292
rect 13688 2252 13694 2264
rect 16206 2252 16212 2264
rect 16264 2252 16270 2304
rect 16546 2292 16574 2604
rect 18877 2601 18889 2635
rect 18923 2632 18935 2635
rect 20438 2632 20444 2644
rect 18923 2604 20444 2632
rect 18923 2601 18935 2604
rect 18877 2595 18935 2601
rect 20438 2592 20444 2604
rect 20496 2592 20502 2644
rect 22922 2632 22928 2644
rect 20824 2604 22928 2632
rect 18966 2524 18972 2576
rect 19024 2564 19030 2576
rect 19024 2536 19472 2564
rect 19024 2524 19030 2536
rect 16942 2456 16948 2508
rect 17000 2496 17006 2508
rect 17129 2499 17187 2505
rect 17129 2496 17141 2499
rect 17000 2468 17141 2496
rect 17000 2456 17006 2468
rect 17129 2465 17141 2468
rect 17175 2465 17187 2499
rect 17129 2459 17187 2465
rect 17405 2499 17463 2505
rect 17405 2465 17417 2499
rect 17451 2496 17463 2499
rect 19242 2496 19248 2508
rect 17451 2468 19248 2496
rect 17451 2465 17463 2468
rect 17405 2459 17463 2465
rect 19242 2456 19248 2468
rect 19300 2456 19306 2508
rect 19444 2505 19472 2536
rect 19429 2499 19487 2505
rect 19429 2465 19441 2499
rect 19475 2465 19487 2499
rect 19429 2459 19487 2465
rect 20824 2414 20852 2604
rect 22922 2592 22928 2604
rect 22980 2592 22986 2644
rect 26602 2632 26608 2644
rect 23032 2604 26608 2632
rect 22005 2567 22063 2573
rect 22005 2533 22017 2567
rect 22051 2564 22063 2567
rect 22370 2564 22376 2576
rect 22051 2536 22376 2564
rect 22051 2533 22063 2536
rect 22005 2527 22063 2533
rect 22370 2524 22376 2536
rect 22428 2524 22434 2576
rect 23032 2505 23060 2604
rect 26602 2592 26608 2604
rect 26660 2592 26666 2644
rect 26694 2592 26700 2644
rect 26752 2632 26758 2644
rect 27249 2635 27307 2641
rect 27249 2632 27261 2635
rect 26752 2604 27261 2632
rect 26752 2592 26758 2604
rect 27249 2601 27261 2604
rect 27295 2601 27307 2635
rect 27249 2595 27307 2601
rect 28350 2592 28356 2644
rect 28408 2632 28414 2644
rect 28537 2635 28595 2641
rect 28537 2632 28549 2635
rect 28408 2604 28549 2632
rect 28408 2592 28414 2604
rect 28537 2601 28549 2604
rect 28583 2601 28595 2635
rect 28537 2595 28595 2601
rect 30558 2564 30564 2576
rect 25792 2536 30564 2564
rect 23017 2499 23075 2505
rect 23017 2465 23029 2499
rect 23063 2465 23075 2499
rect 23017 2459 23075 2465
rect 23934 2456 23940 2508
rect 23992 2496 23998 2508
rect 24029 2499 24087 2505
rect 24029 2496 24041 2499
rect 23992 2468 24041 2496
rect 23992 2456 23998 2468
rect 24029 2465 24041 2468
rect 24075 2496 24087 2499
rect 25130 2496 25136 2508
rect 24075 2468 25136 2496
rect 24075 2465 24087 2468
rect 24029 2459 24087 2465
rect 25130 2456 25136 2468
rect 25188 2456 25194 2508
rect 21266 2388 21272 2440
rect 21324 2428 21330 2440
rect 22189 2431 22247 2437
rect 22189 2428 22201 2431
rect 21324 2400 22201 2428
rect 21324 2388 21330 2400
rect 22189 2397 22201 2400
rect 22235 2397 22247 2431
rect 22189 2391 22247 2397
rect 24581 2431 24639 2437
rect 24581 2397 24593 2431
rect 24627 2397 24639 2431
rect 24854 2428 24860 2440
rect 24815 2400 24860 2428
rect 24581 2391 24639 2397
rect 19426 2360 19432 2372
rect 18630 2332 19432 2360
rect 19426 2320 19432 2332
rect 19484 2320 19490 2372
rect 19702 2360 19708 2372
rect 19663 2332 19708 2360
rect 19702 2320 19708 2332
rect 19760 2320 19766 2372
rect 23106 2360 23112 2372
rect 23067 2332 23112 2360
rect 23106 2320 23112 2332
rect 23164 2320 23170 2372
rect 23198 2320 23204 2372
rect 23256 2360 23262 2372
rect 24596 2360 24624 2391
rect 24854 2388 24860 2400
rect 24912 2388 24918 2440
rect 23256 2332 24624 2360
rect 25792 2360 25820 2536
rect 30558 2524 30564 2536
rect 30616 2524 30622 2576
rect 36081 2567 36139 2573
rect 36081 2533 36093 2567
rect 36127 2564 36139 2567
rect 37090 2564 37096 2576
rect 36127 2536 37096 2564
rect 36127 2533 36139 2536
rect 36081 2527 36139 2533
rect 37090 2524 37096 2536
rect 37148 2524 37154 2576
rect 25958 2496 25964 2508
rect 25919 2468 25964 2496
rect 25958 2456 25964 2468
rect 26016 2456 26022 2508
rect 26418 2456 26424 2508
rect 26476 2496 26482 2508
rect 26476 2468 26521 2496
rect 26476 2456 26482 2468
rect 26602 2456 26608 2508
rect 26660 2496 26666 2508
rect 28442 2496 28448 2508
rect 26660 2468 28448 2496
rect 26660 2456 26666 2468
rect 28442 2456 28448 2468
rect 28500 2456 28506 2508
rect 32582 2496 32588 2508
rect 32543 2468 32588 2496
rect 32582 2456 32588 2468
rect 32640 2456 32646 2508
rect 35342 2456 35348 2508
rect 35400 2496 35406 2508
rect 37734 2496 37740 2508
rect 35400 2468 36676 2496
rect 37695 2468 37740 2496
rect 35400 2456 35406 2468
rect 27154 2428 27160 2440
rect 27115 2400 27160 2428
rect 27154 2388 27160 2400
rect 27212 2388 27218 2440
rect 27706 2388 27712 2440
rect 27764 2428 27770 2440
rect 27801 2431 27859 2437
rect 27801 2428 27813 2431
rect 27764 2400 27813 2428
rect 27764 2388 27770 2400
rect 27801 2397 27813 2400
rect 27847 2397 27859 2431
rect 27801 2391 27859 2397
rect 28721 2431 28779 2437
rect 28721 2397 28733 2431
rect 28767 2397 28779 2431
rect 28721 2391 28779 2397
rect 26053 2363 26111 2369
rect 26053 2360 26065 2363
rect 25792 2332 26065 2360
rect 23256 2320 23262 2332
rect 26053 2329 26065 2332
rect 26099 2329 26111 2363
rect 28736 2360 28764 2391
rect 29362 2388 29368 2440
rect 29420 2428 29426 2440
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29420 2400 29745 2428
rect 29420 2388 29426 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 30469 2431 30527 2437
rect 30469 2397 30481 2431
rect 30515 2428 30527 2431
rect 31018 2428 31024 2440
rect 30515 2400 31024 2428
rect 30515 2397 30527 2400
rect 30469 2391 30527 2397
rect 31018 2388 31024 2400
rect 31076 2388 31082 2440
rect 31205 2431 31263 2437
rect 31205 2397 31217 2431
rect 31251 2428 31263 2431
rect 31294 2428 31300 2440
rect 31251 2400 31300 2428
rect 31251 2397 31263 2400
rect 31205 2391 31263 2397
rect 31294 2388 31300 2400
rect 31352 2388 31358 2440
rect 32214 2388 32220 2440
rect 32272 2428 32278 2440
rect 32309 2431 32367 2437
rect 32309 2428 32321 2431
rect 32272 2400 32321 2428
rect 32272 2388 32278 2400
rect 32309 2397 32321 2400
rect 32355 2397 32367 2431
rect 32309 2391 32367 2397
rect 33410 2388 33416 2440
rect 33468 2428 33474 2440
rect 33597 2431 33655 2437
rect 33597 2428 33609 2431
rect 33468 2400 33609 2428
rect 33468 2388 33474 2400
rect 33597 2397 33609 2400
rect 33643 2397 33655 2431
rect 33597 2391 33655 2397
rect 34790 2388 34796 2440
rect 34848 2428 34854 2440
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 34848 2400 34897 2428
rect 34848 2388 34854 2400
rect 34885 2397 34897 2400
rect 34931 2397 34943 2431
rect 34885 2391 34943 2397
rect 35526 2388 35532 2440
rect 35584 2428 35590 2440
rect 36648 2437 36676 2468
rect 37734 2456 37740 2468
rect 37792 2456 37798 2508
rect 35897 2431 35955 2437
rect 35897 2428 35909 2431
rect 35584 2400 35909 2428
rect 35584 2388 35590 2400
rect 35897 2397 35909 2400
rect 35943 2397 35955 2431
rect 35897 2391 35955 2397
rect 36633 2431 36691 2437
rect 36633 2397 36645 2431
rect 36679 2397 36691 2431
rect 36633 2391 36691 2397
rect 37366 2388 37372 2440
rect 37424 2428 37430 2440
rect 37461 2431 37519 2437
rect 37461 2428 37473 2431
rect 37424 2400 37473 2428
rect 37424 2388 37430 2400
rect 37461 2397 37473 2400
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 26053 2323 26111 2329
rect 26160 2332 28764 2360
rect 18690 2292 18696 2304
rect 16546 2264 18696 2292
rect 18690 2252 18696 2264
rect 18748 2252 18754 2304
rect 19150 2252 19156 2304
rect 19208 2292 19214 2304
rect 21174 2292 21180 2304
rect 19208 2264 21180 2292
rect 19208 2252 19214 2264
rect 21174 2252 21180 2264
rect 21232 2252 21238 2304
rect 22554 2252 22560 2304
rect 22612 2292 22618 2304
rect 26160 2292 26188 2332
rect 22612 2264 26188 2292
rect 22612 2252 22618 2264
rect 27706 2252 27712 2304
rect 27764 2292 27770 2304
rect 27985 2295 28043 2301
rect 27985 2292 27997 2295
rect 27764 2264 27997 2292
rect 27764 2252 27770 2264
rect 27985 2261 27997 2264
rect 28031 2261 28043 2295
rect 27985 2255 28043 2261
rect 28994 2252 29000 2304
rect 29052 2292 29058 2304
rect 29917 2295 29975 2301
rect 29917 2292 29929 2295
rect 29052 2264 29929 2292
rect 29052 2252 29058 2264
rect 29917 2261 29929 2264
rect 29963 2261 29975 2295
rect 29917 2255 29975 2261
rect 30282 2252 30288 2304
rect 30340 2292 30346 2304
rect 30653 2295 30711 2301
rect 30653 2292 30665 2295
rect 30340 2264 30665 2292
rect 30340 2252 30346 2264
rect 30653 2261 30665 2264
rect 30699 2261 30711 2295
rect 31294 2292 31300 2304
rect 31255 2264 31300 2292
rect 30653 2255 30711 2261
rect 31294 2252 31300 2264
rect 31352 2252 31358 2304
rect 33502 2252 33508 2304
rect 33560 2292 33566 2304
rect 33781 2295 33839 2301
rect 33781 2292 33793 2295
rect 33560 2264 33793 2292
rect 33560 2252 33566 2264
rect 33781 2261 33793 2264
rect 33827 2261 33839 2295
rect 33781 2255 33839 2261
rect 34146 2252 34152 2304
rect 34204 2292 34210 2304
rect 35069 2295 35127 2301
rect 35069 2292 35081 2295
rect 34204 2264 35081 2292
rect 34204 2252 34210 2264
rect 35069 2261 35081 2264
rect 35115 2261 35127 2295
rect 35069 2255 35127 2261
rect 36722 2252 36728 2304
rect 36780 2292 36786 2304
rect 36817 2295 36875 2301
rect 36817 2292 36829 2295
rect 36780 2264 36829 2292
rect 36780 2252 36786 2264
rect 36817 2261 36829 2264
rect 36863 2261 36875 2295
rect 36817 2255 36875 2261
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 3418 2048 3424 2100
rect 3476 2088 3482 2100
rect 7466 2088 7472 2100
rect 3476 2060 7472 2088
rect 3476 2048 3482 2060
rect 7466 2048 7472 2060
rect 7524 2048 7530 2100
rect 18046 2088 18052 2100
rect 7576 2060 18052 2088
rect 3786 1980 3792 2032
rect 3844 2020 3850 2032
rect 7576 2020 7604 2060
rect 18046 2048 18052 2060
rect 18104 2048 18110 2100
rect 18506 2048 18512 2100
rect 18564 2088 18570 2100
rect 22738 2088 22744 2100
rect 18564 2060 22744 2088
rect 18564 2048 18570 2060
rect 22738 2048 22744 2060
rect 22796 2048 22802 2100
rect 22922 2048 22928 2100
rect 22980 2088 22986 2100
rect 31110 2088 31116 2100
rect 22980 2060 31116 2088
rect 22980 2048 22986 2060
rect 31110 2048 31116 2060
rect 31168 2048 31174 2100
rect 15286 2020 15292 2032
rect 3844 1992 7604 2020
rect 7760 1992 15292 2020
rect 3844 1980 3850 1992
rect 4706 1844 4712 1896
rect 4764 1884 4770 1896
rect 7760 1884 7788 1992
rect 15286 1980 15292 1992
rect 15344 1980 15350 2032
rect 19058 1980 19064 2032
rect 19116 2020 19122 2032
rect 23014 2020 23020 2032
rect 19116 1992 23020 2020
rect 19116 1980 19122 1992
rect 23014 1980 23020 1992
rect 23072 1980 23078 2032
rect 23106 1980 23112 2032
rect 23164 2020 23170 2032
rect 30374 2020 30380 2032
rect 23164 1992 30380 2020
rect 23164 1980 23170 1992
rect 30374 1980 30380 1992
rect 30432 1980 30438 2032
rect 11146 1912 11152 1964
rect 11204 1952 11210 1964
rect 15470 1952 15476 1964
rect 11204 1924 15476 1952
rect 11204 1912 11210 1924
rect 15470 1912 15476 1924
rect 15528 1912 15534 1964
rect 15746 1912 15752 1964
rect 15804 1952 15810 1964
rect 27154 1952 27160 1964
rect 15804 1924 27160 1952
rect 15804 1912 15810 1924
rect 27154 1912 27160 1924
rect 27212 1912 27218 1964
rect 4764 1856 7788 1884
rect 4764 1844 4770 1856
rect 16298 1844 16304 1896
rect 16356 1884 16362 1896
rect 22830 1884 22836 1896
rect 16356 1856 22836 1884
rect 16356 1844 16362 1856
rect 22830 1844 22836 1856
rect 22888 1844 22894 1896
rect 24946 1844 24952 1896
rect 25004 1884 25010 1896
rect 31294 1884 31300 1896
rect 25004 1856 31300 1884
rect 25004 1844 25010 1856
rect 31294 1844 31300 1856
rect 31352 1844 31358 1896
rect 4522 1776 4528 1828
rect 4580 1816 4586 1828
rect 11054 1816 11060 1828
rect 4580 1788 11060 1816
rect 4580 1776 4586 1788
rect 11054 1776 11060 1788
rect 11112 1816 11118 1828
rect 13446 1816 13452 1828
rect 11112 1788 13452 1816
rect 11112 1776 11118 1788
rect 13446 1776 13452 1788
rect 13504 1776 13510 1828
rect 21174 1776 21180 1828
rect 21232 1816 21238 1828
rect 27890 1816 27896 1828
rect 21232 1788 27896 1816
rect 21232 1776 21238 1788
rect 27890 1776 27896 1788
rect 27948 1776 27954 1828
rect 2314 1708 2320 1760
rect 2372 1748 2378 1760
rect 8478 1748 8484 1760
rect 2372 1720 8484 1748
rect 2372 1708 2378 1720
rect 8478 1708 8484 1720
rect 8536 1748 8542 1760
rect 11698 1748 11704 1760
rect 8536 1720 11704 1748
rect 8536 1708 8542 1720
rect 11698 1708 11704 1720
rect 11756 1708 11762 1760
rect 24854 1748 24860 1760
rect 16546 1720 24860 1748
rect 8662 1640 8668 1692
rect 8720 1680 8726 1692
rect 16546 1680 16574 1720
rect 24854 1708 24860 1720
rect 24912 1708 24918 1760
rect 25774 1708 25780 1760
rect 25832 1748 25838 1760
rect 27614 1748 27620 1760
rect 25832 1720 27620 1748
rect 25832 1708 25838 1720
rect 27614 1708 27620 1720
rect 27672 1708 27678 1760
rect 8720 1652 16574 1680
rect 8720 1640 8726 1652
rect 18782 1640 18788 1692
rect 18840 1680 18846 1692
rect 19978 1680 19984 1692
rect 18840 1652 19984 1680
rect 18840 1640 18846 1652
rect 19978 1640 19984 1652
rect 20036 1640 20042 1692
rect 23014 1640 23020 1692
rect 23072 1680 23078 1692
rect 30466 1680 30472 1692
rect 23072 1652 30472 1680
rect 23072 1640 23078 1652
rect 30466 1640 30472 1652
rect 30524 1640 30530 1692
rect 6270 1572 6276 1624
rect 6328 1612 6334 1624
rect 12250 1612 12256 1624
rect 6328 1584 12256 1612
rect 6328 1572 6334 1584
rect 12250 1572 12256 1584
rect 12308 1572 12314 1624
rect 16206 1572 16212 1624
rect 16264 1612 16270 1624
rect 29086 1612 29092 1624
rect 16264 1584 29092 1612
rect 16264 1572 16270 1584
rect 29086 1572 29092 1584
rect 29144 1572 29150 1624
rect 19426 1504 19432 1556
rect 19484 1544 19490 1556
rect 31662 1544 31668 1556
rect 19484 1516 31668 1544
rect 19484 1504 19490 1516
rect 31662 1504 31668 1516
rect 31720 1504 31726 1556
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 20168 37340 20220 37392
rect 36820 37340 36872 37392
rect 39304 37340 39356 37392
rect 1952 37272 2004 37324
rect 3884 37272 3936 37324
rect 8392 37272 8444 37324
rect 22468 37272 22520 37324
rect 22560 37272 22612 37324
rect 29644 37272 29696 37324
rect 2504 37204 2556 37256
rect 5172 37204 5224 37256
rect 5816 37204 5868 37256
rect 7104 37204 7156 37256
rect 8300 37204 8352 37256
rect 10416 37247 10468 37256
rect 10416 37213 10425 37247
rect 10425 37213 10459 37247
rect 10459 37213 10468 37247
rect 10416 37204 10468 37213
rect 11612 37204 11664 37256
rect 12440 37247 12492 37256
rect 12440 37213 12449 37247
rect 12449 37213 12483 37247
rect 12483 37213 12492 37247
rect 12440 37204 12492 37213
rect 13544 37204 13596 37256
rect 15200 37247 15252 37256
rect 15200 37213 15209 37247
rect 15209 37213 15243 37247
rect 15243 37213 15252 37247
rect 15200 37204 15252 37213
rect 16028 37247 16080 37256
rect 16028 37213 16037 37247
rect 16037 37213 16071 37247
rect 16071 37213 16080 37247
rect 16028 37204 16080 37213
rect 16948 37204 17000 37256
rect 18052 37204 18104 37256
rect 20076 37247 20128 37256
rect 20076 37213 20085 37247
rect 20085 37213 20119 37247
rect 20119 37213 20128 37247
rect 20076 37204 20128 37213
rect 21180 37247 21232 37256
rect 21180 37213 21189 37247
rect 21189 37213 21223 37247
rect 21223 37213 21232 37247
rect 21180 37204 21232 37213
rect 22928 37247 22980 37256
rect 22928 37213 22937 37247
rect 22937 37213 22971 37247
rect 22971 37213 22980 37247
rect 22928 37204 22980 37213
rect 24492 37204 24544 37256
rect 25780 37204 25832 37256
rect 27160 37247 27212 37256
rect 27160 37213 27169 37247
rect 27169 37213 27203 37247
rect 27203 37213 27212 37247
rect 27160 37204 27212 37213
rect 27712 37204 27764 37256
rect 29000 37204 29052 37256
rect 38660 37272 38712 37324
rect 31024 37247 31076 37256
rect 31024 37213 31033 37247
rect 31033 37213 31067 37247
rect 31067 37213 31076 37247
rect 31024 37204 31076 37213
rect 32220 37204 32272 37256
rect 10508 37136 10560 37188
rect 25504 37136 25556 37188
rect 33232 37204 33284 37256
rect 35992 37204 36044 37256
rect 37740 37247 37792 37256
rect 37740 37213 37749 37247
rect 37749 37213 37783 37247
rect 37783 37213 37792 37247
rect 37740 37204 37792 37213
rect 6184 37068 6236 37120
rect 6552 37111 6604 37120
rect 6552 37077 6561 37111
rect 6561 37077 6595 37111
rect 6595 37077 6604 37111
rect 6552 37068 6604 37077
rect 7932 37068 7984 37120
rect 10324 37068 10376 37120
rect 11704 37111 11756 37120
rect 11704 37077 11713 37111
rect 11713 37077 11747 37111
rect 11747 37077 11756 37111
rect 11704 37068 11756 37077
rect 15016 37111 15068 37120
rect 15016 37077 15025 37111
rect 15025 37077 15059 37111
rect 15059 37077 15068 37111
rect 15016 37068 15068 37077
rect 16120 37068 16172 37120
rect 16764 37068 16816 37120
rect 17132 37068 17184 37120
rect 19984 37068 20036 37120
rect 21272 37068 21324 37120
rect 24584 37111 24636 37120
rect 24584 37077 24593 37111
rect 24593 37077 24627 37111
rect 24627 37077 24636 37111
rect 24584 37068 24636 37077
rect 25872 37111 25924 37120
rect 25872 37077 25881 37111
rect 25881 37077 25915 37111
rect 25915 37077 25924 37111
rect 25872 37068 25924 37077
rect 26424 37068 26476 37120
rect 27436 37068 27488 37120
rect 29736 37111 29788 37120
rect 29736 37077 29745 37111
rect 29745 37077 29779 37111
rect 29779 37077 29788 37111
rect 29736 37068 29788 37077
rect 30380 37111 30432 37120
rect 30380 37077 30389 37111
rect 30389 37077 30423 37111
rect 30423 37077 30432 37111
rect 30380 37068 30432 37077
rect 30932 37068 30984 37120
rect 31300 37068 31352 37120
rect 33140 37111 33192 37120
rect 33140 37077 33149 37111
rect 33149 37077 33183 37111
rect 33183 37077 33192 37111
rect 33140 37068 33192 37077
rect 34520 37068 34572 37120
rect 36084 37068 36136 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 664 36864 716 36916
rect 2964 36796 3016 36848
rect 2780 36728 2832 36780
rect 6552 36864 6604 36916
rect 9956 36864 10008 36916
rect 10416 36907 10468 36916
rect 10416 36873 10425 36907
rect 10425 36873 10459 36907
rect 10459 36873 10468 36907
rect 10416 36864 10468 36873
rect 19340 36864 19392 36916
rect 23204 36864 23256 36916
rect 27160 36907 27212 36916
rect 27160 36873 27169 36907
rect 27169 36873 27203 36907
rect 27203 36873 27212 36907
rect 27160 36864 27212 36873
rect 27988 36864 28040 36916
rect 31024 36864 31076 36916
rect 36176 36864 36228 36916
rect 36820 36907 36872 36916
rect 36820 36873 36829 36907
rect 36829 36873 36863 36907
rect 36863 36873 36872 36907
rect 36820 36864 36872 36873
rect 37372 36864 37424 36916
rect 9036 36728 9088 36780
rect 10508 36728 10560 36780
rect 19432 36771 19484 36780
rect 19432 36737 19441 36771
rect 19441 36737 19475 36771
rect 19475 36737 19484 36771
rect 19432 36728 19484 36737
rect 23296 36771 23348 36780
rect 23296 36737 23305 36771
rect 23305 36737 23339 36771
rect 23339 36737 23348 36771
rect 23296 36728 23348 36737
rect 35440 36771 35492 36780
rect 35440 36737 35449 36771
rect 35449 36737 35483 36771
rect 35483 36737 35492 36771
rect 35440 36728 35492 36737
rect 35900 36771 35952 36780
rect 35900 36737 35909 36771
rect 35909 36737 35943 36771
rect 35943 36737 35952 36771
rect 36636 36771 36688 36780
rect 35900 36728 35952 36737
rect 36636 36737 36645 36771
rect 36645 36737 36679 36771
rect 36679 36737 36688 36771
rect 36636 36728 36688 36737
rect 37372 36728 37424 36780
rect 27528 36660 27580 36712
rect 37740 36660 37792 36712
rect 1860 36635 1912 36644
rect 1860 36601 1869 36635
rect 1869 36601 1903 36635
rect 1903 36601 1912 36635
rect 1860 36592 1912 36601
rect 3240 36524 3292 36576
rect 6552 36524 6604 36576
rect 9772 36524 9824 36576
rect 32128 36524 32180 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 1768 36363 1820 36372
rect 1768 36329 1777 36363
rect 1777 36329 1811 36363
rect 1811 36329 1820 36363
rect 1768 36320 1820 36329
rect 36636 36363 36688 36372
rect 36636 36329 36645 36363
rect 36645 36329 36679 36363
rect 36679 36329 36688 36363
rect 36636 36320 36688 36329
rect 1584 36159 1636 36168
rect 1584 36125 1593 36159
rect 1593 36125 1627 36159
rect 1627 36125 1636 36159
rect 1584 36116 1636 36125
rect 2872 36116 2924 36168
rect 36820 36159 36872 36168
rect 36820 36125 36829 36159
rect 36829 36125 36863 36159
rect 36863 36125 36872 36159
rect 36820 36116 36872 36125
rect 37188 36116 37240 36168
rect 37832 36116 37884 36168
rect 6460 35980 6512 36032
rect 37280 35980 37332 36032
rect 38200 36023 38252 36032
rect 38200 35989 38209 36023
rect 38209 35989 38243 36023
rect 38243 35989 38252 36023
rect 38200 35980 38252 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 36820 35776 36872 35828
rect 1768 35683 1820 35692
rect 1768 35649 1777 35683
rect 1777 35649 1811 35683
rect 1811 35649 1820 35683
rect 1768 35640 1820 35649
rect 14464 35640 14516 35692
rect 32404 35572 32456 35624
rect 5540 35436 5592 35488
rect 38200 35479 38252 35488
rect 38200 35445 38209 35479
rect 38209 35445 38243 35479
rect 38243 35445 38252 35479
rect 38200 35436 38252 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 16028 35232 16080 35284
rect 13912 35028 13964 35080
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 3056 34552 3108 34604
rect 3240 34552 3292 34604
rect 38016 34595 38068 34604
rect 38016 34561 38025 34595
rect 38025 34561 38059 34595
rect 38059 34561 38068 34595
rect 38016 34552 38068 34561
rect 6736 34484 6788 34536
rect 1768 34391 1820 34400
rect 1768 34357 1777 34391
rect 1777 34357 1811 34391
rect 1811 34357 1820 34391
rect 1768 34348 1820 34357
rect 38200 34391 38252 34400
rect 38200 34357 38209 34391
rect 38209 34357 38243 34391
rect 38243 34357 38252 34391
rect 38200 34348 38252 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 19432 33600 19484 33652
rect 11704 33464 11756 33516
rect 24676 33464 24728 33516
rect 18604 33260 18656 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 35992 33056 36044 33108
rect 2504 32895 2556 32904
rect 1768 32759 1820 32768
rect 1768 32725 1777 32759
rect 1777 32725 1811 32759
rect 1811 32725 1820 32759
rect 1768 32716 1820 32725
rect 2504 32861 2513 32895
rect 2513 32861 2547 32895
rect 2547 32861 2556 32895
rect 2504 32852 2556 32861
rect 31116 32852 31168 32904
rect 37464 32895 37516 32904
rect 37464 32861 37473 32895
rect 37473 32861 37507 32895
rect 37507 32861 37516 32895
rect 37464 32852 37516 32861
rect 38384 32852 38436 32904
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 33232 32512 33284 32564
rect 1860 32376 1912 32428
rect 29644 32376 29696 32428
rect 38292 32419 38344 32428
rect 38292 32385 38301 32419
rect 38301 32385 38335 32419
rect 38335 32385 38344 32419
rect 38292 32376 38344 32385
rect 25688 32240 25740 32292
rect 29736 32240 29788 32292
rect 1768 32215 1820 32224
rect 1768 32181 1777 32215
rect 1777 32181 1811 32215
rect 1811 32181 1820 32215
rect 1768 32172 1820 32181
rect 37648 32172 37700 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 23296 31968 23348 32020
rect 27988 32011 28040 32020
rect 27988 31977 27997 32011
rect 27997 31977 28031 32011
rect 28031 31977 28040 32011
rect 27988 31968 28040 31977
rect 31116 32011 31168 32020
rect 31116 31977 31125 32011
rect 31125 31977 31159 32011
rect 31159 31977 31168 32011
rect 31116 31968 31168 31977
rect 38016 31968 38068 32020
rect 23204 31900 23256 31952
rect 21272 31832 21324 31884
rect 27252 31832 27304 31884
rect 7932 31807 7984 31816
rect 7932 31773 7941 31807
rect 7941 31773 7975 31807
rect 7975 31773 7984 31807
rect 7932 31764 7984 31773
rect 8116 31764 8168 31816
rect 21548 31764 21600 31816
rect 25688 31807 25740 31816
rect 25688 31773 25697 31807
rect 25697 31773 25731 31807
rect 25731 31773 25740 31807
rect 25688 31764 25740 31773
rect 26884 31764 26936 31816
rect 30380 31832 30432 31884
rect 37096 31807 37148 31816
rect 37096 31773 37105 31807
rect 37105 31773 37139 31807
rect 37139 31773 37148 31807
rect 37096 31764 37148 31773
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 35900 31424 35952 31476
rect 6184 31356 6236 31408
rect 6552 31331 6604 31340
rect 6552 31297 6561 31331
rect 6561 31297 6595 31331
rect 6595 31297 6604 31331
rect 6552 31288 6604 31297
rect 17132 31288 17184 31340
rect 30380 31288 30432 31340
rect 6828 31084 6880 31136
rect 7380 31084 7432 31136
rect 15476 31084 15528 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 3056 30880 3108 30932
rect 37096 30880 37148 30932
rect 8484 30676 8536 30728
rect 9956 30676 10008 30728
rect 24584 30744 24636 30796
rect 25872 30676 25924 30728
rect 32128 30676 32180 30728
rect 36176 30719 36228 30728
rect 36176 30685 36185 30719
rect 36185 30685 36219 30719
rect 36219 30685 36228 30719
rect 36176 30676 36228 30685
rect 38292 30719 38344 30728
rect 38292 30685 38301 30719
rect 38301 30685 38335 30719
rect 38335 30685 38344 30719
rect 38292 30676 38344 30685
rect 6276 30608 6328 30660
rect 18420 30608 18472 30660
rect 1768 30583 1820 30592
rect 1768 30549 1777 30583
rect 1777 30549 1811 30583
rect 1811 30549 1820 30583
rect 1768 30540 1820 30549
rect 10232 30540 10284 30592
rect 21916 30583 21968 30592
rect 21916 30549 21925 30583
rect 21925 30549 21959 30583
rect 21959 30549 21968 30583
rect 21916 30540 21968 30549
rect 28080 30583 28132 30592
rect 28080 30549 28089 30583
rect 28089 30549 28123 30583
rect 28123 30549 28132 30583
rect 28080 30540 28132 30549
rect 38016 30540 38068 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 17960 30336 18012 30388
rect 28080 30336 28132 30388
rect 13912 30311 13964 30320
rect 13912 30277 13921 30311
rect 13921 30277 13955 30311
rect 13955 30277 13964 30311
rect 13912 30268 13964 30277
rect 6460 30200 6512 30252
rect 13452 30200 13504 30252
rect 15016 30200 15068 30252
rect 27436 30268 27488 30320
rect 29644 30311 29696 30320
rect 29644 30277 29653 30311
rect 29653 30277 29687 30311
rect 29687 30277 29696 30311
rect 29644 30268 29696 30277
rect 29552 30243 29604 30252
rect 29552 30209 29561 30243
rect 29561 30209 29595 30243
rect 29595 30209 29604 30243
rect 29552 30200 29604 30209
rect 37740 30200 37792 30252
rect 31300 30132 31352 30184
rect 15568 30064 15620 30116
rect 37832 30107 37884 30116
rect 37832 30073 37841 30107
rect 37841 30073 37875 30107
rect 37875 30073 37884 30107
rect 37832 30064 37884 30073
rect 6644 30039 6696 30048
rect 6644 30005 6653 30039
rect 6653 30005 6687 30039
rect 6687 30005 6696 30039
rect 6644 29996 6696 30005
rect 13084 29996 13136 30048
rect 23572 29996 23624 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 21548 29835 21600 29844
rect 21548 29801 21557 29835
rect 21557 29801 21591 29835
rect 21591 29801 21600 29835
rect 21548 29792 21600 29801
rect 30380 29792 30432 29844
rect 1492 29588 1544 29640
rect 9772 29588 9824 29640
rect 15016 29588 15068 29640
rect 27160 29588 27212 29640
rect 38108 29563 38160 29572
rect 38108 29529 38117 29563
rect 38117 29529 38151 29563
rect 38151 29529 38160 29563
rect 38108 29520 38160 29529
rect 1768 29495 1820 29504
rect 1768 29461 1777 29495
rect 1777 29461 1811 29495
rect 1811 29461 1820 29495
rect 1768 29452 1820 29461
rect 11428 29452 11480 29504
rect 38200 29495 38252 29504
rect 38200 29461 38209 29495
rect 38209 29461 38243 29495
rect 38243 29461 38252 29495
rect 38200 29452 38252 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 21180 29248 21232 29300
rect 1768 29155 1820 29164
rect 1768 29121 1777 29155
rect 1777 29121 1811 29155
rect 1811 29121 1820 29155
rect 1768 29112 1820 29121
rect 10508 29112 10560 29164
rect 22100 29112 22152 29164
rect 38292 29155 38344 29164
rect 38292 29121 38301 29155
rect 38301 29121 38335 29155
rect 38335 29121 38344 29155
rect 38292 29112 38344 29121
rect 1952 28976 2004 29028
rect 11336 28976 11388 29028
rect 17592 28976 17644 29028
rect 21916 28976 21968 29028
rect 37924 28976 37976 29028
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 6276 28747 6328 28756
rect 6276 28713 6285 28747
rect 6285 28713 6319 28747
rect 6319 28713 6328 28747
rect 6276 28704 6328 28713
rect 8208 28500 8260 28552
rect 10324 28500 10376 28552
rect 27528 28543 27580 28552
rect 27528 28509 27537 28543
rect 27537 28509 27571 28543
rect 27571 28509 27580 28543
rect 27528 28500 27580 28509
rect 11520 28407 11572 28416
rect 11520 28373 11529 28407
rect 11529 28373 11563 28407
rect 11563 28373 11572 28407
rect 11520 28364 11572 28373
rect 27804 28364 27856 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 10324 28203 10376 28212
rect 10324 28169 10333 28203
rect 10333 28169 10367 28203
rect 10367 28169 10376 28203
rect 10324 28160 10376 28169
rect 5540 28024 5592 28076
rect 11152 28067 11204 28076
rect 11152 28033 11161 28067
rect 11161 28033 11195 28067
rect 11195 28033 11204 28067
rect 11152 28024 11204 28033
rect 11612 27956 11664 28008
rect 11980 28024 12032 28076
rect 12992 28024 13044 28076
rect 12072 27888 12124 27940
rect 9220 27863 9272 27872
rect 9220 27829 9229 27863
rect 9229 27829 9263 27863
rect 9263 27829 9272 27863
rect 9220 27820 9272 27829
rect 11888 27863 11940 27872
rect 11888 27829 11897 27863
rect 11897 27829 11931 27863
rect 11931 27829 11940 27863
rect 11888 27820 11940 27829
rect 12716 27863 12768 27872
rect 12716 27829 12725 27863
rect 12725 27829 12759 27863
rect 12759 27829 12768 27863
rect 12716 27820 12768 27829
rect 13268 27863 13320 27872
rect 13268 27829 13277 27863
rect 13277 27829 13311 27863
rect 13311 27829 13320 27863
rect 13268 27820 13320 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 9220 27616 9272 27668
rect 21824 27616 21876 27668
rect 11152 27548 11204 27600
rect 13452 27591 13504 27600
rect 13452 27557 13461 27591
rect 13461 27557 13495 27591
rect 13495 27557 13504 27591
rect 13452 27548 13504 27557
rect 17684 27548 17736 27600
rect 25504 27548 25556 27600
rect 11888 27523 11940 27532
rect 11888 27489 11897 27523
rect 11897 27489 11931 27523
rect 11931 27489 11940 27523
rect 11888 27480 11940 27489
rect 1584 27455 1636 27464
rect 1584 27421 1593 27455
rect 1593 27421 1627 27455
rect 1627 27421 1636 27455
rect 1584 27412 1636 27421
rect 5540 27412 5592 27464
rect 12532 27480 12584 27532
rect 12716 27480 12768 27532
rect 10968 27344 11020 27396
rect 12440 27412 12492 27464
rect 38200 27480 38252 27532
rect 38292 27455 38344 27464
rect 38292 27421 38301 27455
rect 38301 27421 38335 27455
rect 38335 27421 38344 27455
rect 38292 27412 38344 27421
rect 11152 27276 11204 27328
rect 11980 27276 12032 27328
rect 14740 27319 14792 27328
rect 14740 27285 14749 27319
rect 14749 27285 14783 27319
rect 14783 27285 14792 27319
rect 14740 27276 14792 27285
rect 34612 27276 34664 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 12440 27115 12492 27124
rect 12440 27081 12449 27115
rect 12449 27081 12483 27115
rect 12483 27081 12492 27115
rect 12440 27072 12492 27081
rect 13452 27072 13504 27124
rect 10968 27047 11020 27056
rect 10968 27013 10977 27047
rect 10977 27013 11011 27047
rect 11011 27013 11020 27047
rect 10968 27004 11020 27013
rect 10048 26936 10100 26988
rect 9404 26868 9456 26920
rect 12256 27004 12308 27056
rect 11520 26936 11572 26988
rect 12072 26936 12124 26988
rect 14004 26936 14056 26988
rect 15384 26979 15436 26988
rect 15384 26945 15393 26979
rect 15393 26945 15427 26979
rect 15427 26945 15436 26979
rect 15384 26936 15436 26945
rect 21916 26936 21968 26988
rect 11796 26911 11848 26920
rect 11796 26877 11805 26911
rect 11805 26877 11839 26911
rect 11839 26877 11848 26911
rect 11796 26868 11848 26877
rect 12900 26911 12952 26920
rect 12900 26877 12909 26911
rect 12909 26877 12943 26911
rect 12943 26877 12952 26911
rect 12900 26868 12952 26877
rect 12808 26800 12860 26852
rect 11060 26775 11112 26784
rect 11060 26741 11069 26775
rect 11069 26741 11103 26775
rect 11103 26741 11112 26775
rect 11060 26732 11112 26741
rect 14556 26775 14608 26784
rect 14556 26741 14565 26775
rect 14565 26741 14599 26775
rect 14599 26741 14608 26775
rect 14556 26732 14608 26741
rect 15200 26775 15252 26784
rect 15200 26741 15209 26775
rect 15209 26741 15243 26775
rect 15243 26741 15252 26775
rect 15200 26732 15252 26741
rect 23296 26732 23348 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 9404 26571 9456 26580
rect 9404 26537 9413 26571
rect 9413 26537 9447 26571
rect 9447 26537 9456 26571
rect 9404 26528 9456 26537
rect 10048 26571 10100 26580
rect 10048 26537 10057 26571
rect 10057 26537 10091 26571
rect 10091 26537 10100 26571
rect 10048 26528 10100 26537
rect 10692 26528 10744 26580
rect 12624 26528 12676 26580
rect 15384 26528 15436 26580
rect 20352 26528 20404 26580
rect 33784 26528 33836 26580
rect 34520 26460 34572 26512
rect 6736 26392 6788 26444
rect 12808 26392 12860 26444
rect 2504 26324 2556 26376
rect 10508 26324 10560 26376
rect 10692 26367 10744 26376
rect 10692 26333 10701 26367
rect 10701 26333 10735 26367
rect 10735 26333 10744 26367
rect 10692 26324 10744 26333
rect 11612 26324 11664 26376
rect 12072 26324 12124 26376
rect 1676 26299 1728 26308
rect 1676 26265 1685 26299
rect 1685 26265 1719 26299
rect 1719 26265 1728 26299
rect 1676 26256 1728 26265
rect 8208 26256 8260 26308
rect 12992 26256 13044 26308
rect 14188 26324 14240 26376
rect 15108 26392 15160 26444
rect 20812 26367 20864 26376
rect 20812 26333 20821 26367
rect 20821 26333 20855 26367
rect 20855 26333 20864 26367
rect 20812 26324 20864 26333
rect 12900 26188 12952 26240
rect 13452 26188 13504 26240
rect 17960 26256 18012 26308
rect 18236 26256 18288 26308
rect 21916 26324 21968 26376
rect 38292 26367 38344 26376
rect 38292 26333 38301 26367
rect 38301 26333 38335 26367
rect 38335 26333 38344 26367
rect 38292 26324 38344 26333
rect 15292 26188 15344 26240
rect 22468 26231 22520 26240
rect 22468 26197 22477 26231
rect 22477 26197 22511 26231
rect 22511 26197 22520 26231
rect 22468 26188 22520 26197
rect 23112 26231 23164 26240
rect 23112 26197 23121 26231
rect 23121 26197 23155 26231
rect 23155 26197 23164 26231
rect 23112 26188 23164 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 14004 26027 14056 26036
rect 1768 25916 1820 25968
rect 8484 25916 8536 25968
rect 10784 25916 10836 25968
rect 14004 25993 14013 26027
rect 14013 25993 14047 26027
rect 14047 25993 14056 26027
rect 14004 25984 14056 25993
rect 15292 26027 15344 26036
rect 15292 25993 15301 26027
rect 15301 25993 15335 26027
rect 15335 25993 15344 26027
rect 15292 25984 15344 25993
rect 18420 25959 18472 25968
rect 9956 25848 10008 25900
rect 10508 25891 10560 25900
rect 10508 25857 10517 25891
rect 10517 25857 10551 25891
rect 10551 25857 10560 25891
rect 10508 25848 10560 25857
rect 13176 25848 13228 25900
rect 14188 25891 14240 25900
rect 14188 25857 14197 25891
rect 14197 25857 14231 25891
rect 14231 25857 14240 25891
rect 14188 25848 14240 25857
rect 14740 25848 14792 25900
rect 15200 25848 15252 25900
rect 15752 25848 15804 25900
rect 18420 25925 18429 25959
rect 18429 25925 18463 25959
rect 18463 25925 18472 25959
rect 18420 25916 18472 25925
rect 19524 25916 19576 25968
rect 24216 25916 24268 25968
rect 19340 25848 19392 25900
rect 21824 25848 21876 25900
rect 23112 25891 23164 25900
rect 23112 25857 23121 25891
rect 23121 25857 23155 25891
rect 23155 25857 23164 25891
rect 23112 25848 23164 25857
rect 23296 25891 23348 25900
rect 23296 25857 23305 25891
rect 23305 25857 23339 25891
rect 23339 25857 23348 25891
rect 23296 25848 23348 25857
rect 38108 25848 38160 25900
rect 11796 25780 11848 25832
rect 17960 25780 18012 25832
rect 19248 25823 19300 25832
rect 19248 25789 19257 25823
rect 19257 25789 19291 25823
rect 19291 25789 19300 25823
rect 19248 25780 19300 25789
rect 22192 25823 22244 25832
rect 22192 25789 22201 25823
rect 22201 25789 22235 25823
rect 22235 25789 22244 25823
rect 22192 25780 22244 25789
rect 15200 25712 15252 25764
rect 22928 25712 22980 25764
rect 12164 25644 12216 25696
rect 21272 25644 21324 25696
rect 24400 25644 24452 25696
rect 24768 25644 24820 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 10784 25483 10836 25492
rect 10784 25449 10793 25483
rect 10793 25449 10827 25483
rect 10827 25449 10836 25483
rect 10784 25440 10836 25449
rect 12624 25483 12676 25492
rect 12624 25449 12633 25483
rect 12633 25449 12667 25483
rect 12667 25449 12676 25483
rect 12624 25440 12676 25449
rect 13452 25483 13504 25492
rect 13452 25449 13461 25483
rect 13461 25449 13495 25483
rect 13495 25449 13504 25483
rect 13452 25440 13504 25449
rect 11796 25372 11848 25424
rect 14648 25372 14700 25424
rect 13268 25347 13320 25356
rect 13268 25313 13277 25347
rect 13277 25313 13311 25347
rect 13311 25313 13320 25347
rect 13268 25304 13320 25313
rect 1952 25236 2004 25288
rect 2136 25236 2188 25288
rect 10692 25279 10744 25288
rect 10692 25245 10701 25279
rect 10701 25245 10735 25279
rect 10735 25245 10744 25279
rect 10692 25236 10744 25245
rect 12164 25279 12216 25288
rect 12164 25245 12173 25279
rect 12173 25245 12207 25279
rect 12207 25245 12216 25279
rect 12164 25236 12216 25245
rect 16396 25440 16448 25492
rect 19524 25483 19576 25492
rect 19524 25449 19533 25483
rect 19533 25449 19567 25483
rect 19567 25449 19576 25483
rect 19524 25440 19576 25449
rect 24676 25483 24728 25492
rect 24676 25449 24685 25483
rect 24685 25449 24719 25483
rect 24719 25449 24728 25483
rect 24676 25440 24728 25449
rect 15108 25372 15160 25424
rect 17960 25372 18012 25424
rect 21180 25347 21232 25356
rect 15200 25236 15252 25288
rect 21180 25313 21189 25347
rect 21189 25313 21223 25347
rect 21223 25313 21232 25347
rect 21180 25304 21232 25313
rect 21456 25347 21508 25356
rect 21456 25313 21465 25347
rect 21465 25313 21499 25347
rect 21499 25313 21508 25347
rect 21456 25304 21508 25313
rect 16396 25236 16448 25288
rect 19340 25236 19392 25288
rect 22468 25236 22520 25288
rect 27436 25236 27488 25288
rect 34520 25236 34572 25288
rect 38016 25279 38068 25288
rect 38016 25245 38025 25279
rect 38025 25245 38059 25279
rect 38059 25245 38068 25279
rect 38016 25236 38068 25245
rect 14740 25168 14792 25220
rect 21272 25211 21324 25220
rect 21272 25177 21281 25211
rect 21281 25177 21315 25211
rect 21315 25177 21324 25211
rect 21272 25168 21324 25177
rect 14372 25143 14424 25152
rect 14372 25109 14381 25143
rect 14381 25109 14415 25143
rect 14415 25109 14424 25143
rect 14372 25100 14424 25109
rect 15200 25143 15252 25152
rect 15200 25109 15209 25143
rect 15209 25109 15243 25143
rect 15243 25109 15252 25143
rect 15200 25100 15252 25109
rect 17224 25100 17276 25152
rect 24768 25100 24820 25152
rect 31208 25143 31260 25152
rect 31208 25109 31217 25143
rect 31217 25109 31251 25143
rect 31251 25109 31260 25143
rect 31208 25100 31260 25109
rect 38200 25143 38252 25152
rect 38200 25109 38209 25143
rect 38209 25109 38243 25143
rect 38243 25109 38252 25143
rect 38200 25100 38252 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 14372 24828 14424 24880
rect 19248 24896 19300 24948
rect 22192 24896 22244 24948
rect 4068 24760 4120 24812
rect 8668 24760 8720 24812
rect 10692 24760 10744 24812
rect 11612 24760 11664 24812
rect 12072 24760 12124 24812
rect 12900 24760 12952 24812
rect 12716 24692 12768 24744
rect 13084 24735 13136 24744
rect 13084 24701 13093 24735
rect 13093 24701 13127 24735
rect 13127 24701 13136 24735
rect 13084 24692 13136 24701
rect 13360 24692 13412 24744
rect 15200 24692 15252 24744
rect 16304 24760 16356 24812
rect 22928 24871 22980 24880
rect 22928 24837 22937 24871
rect 22937 24837 22971 24871
rect 22971 24837 22980 24871
rect 22928 24828 22980 24837
rect 19984 24760 20036 24812
rect 21916 24760 21968 24812
rect 24308 24760 24360 24812
rect 25780 24803 25832 24812
rect 25780 24769 25789 24803
rect 25789 24769 25823 24803
rect 25823 24769 25832 24803
rect 25780 24760 25832 24769
rect 26884 24760 26936 24812
rect 37648 24760 37700 24812
rect 15108 24624 15160 24676
rect 18052 24692 18104 24744
rect 20720 24692 20772 24744
rect 1768 24599 1820 24608
rect 1768 24565 1777 24599
rect 1777 24565 1811 24599
rect 1811 24565 1820 24599
rect 1768 24556 1820 24565
rect 10324 24556 10376 24608
rect 12624 24556 12676 24608
rect 31208 24692 31260 24744
rect 27160 24624 27212 24676
rect 27528 24624 27580 24676
rect 22836 24556 22888 24608
rect 22928 24556 22980 24608
rect 30656 24556 30708 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 14648 24352 14700 24404
rect 23112 24352 23164 24404
rect 25780 24352 25832 24404
rect 11888 24284 11940 24336
rect 16856 24284 16908 24336
rect 17684 24327 17736 24336
rect 17684 24293 17693 24327
rect 17693 24293 17727 24327
rect 17727 24293 17736 24327
rect 17684 24284 17736 24293
rect 23296 24284 23348 24336
rect 24860 24284 24912 24336
rect 12532 24259 12584 24268
rect 12532 24225 12541 24259
rect 12541 24225 12575 24259
rect 12575 24225 12584 24259
rect 12532 24216 12584 24225
rect 12900 24216 12952 24268
rect 13268 24216 13320 24268
rect 14556 24259 14608 24268
rect 1584 24191 1636 24200
rect 1584 24157 1593 24191
rect 1593 24157 1627 24191
rect 1627 24157 1636 24191
rect 1584 24148 1636 24157
rect 1860 24191 1912 24200
rect 1860 24157 1869 24191
rect 1869 24157 1903 24191
rect 1903 24157 1912 24191
rect 1860 24148 1912 24157
rect 12624 24123 12676 24132
rect 12624 24089 12633 24123
rect 12633 24089 12667 24123
rect 12667 24089 12676 24123
rect 12624 24080 12676 24089
rect 13728 24080 13780 24132
rect 14556 24225 14565 24259
rect 14565 24225 14599 24259
rect 14599 24225 14608 24259
rect 14556 24216 14608 24225
rect 22100 24216 22152 24268
rect 24584 24259 24636 24268
rect 15200 24148 15252 24200
rect 15292 24148 15344 24200
rect 15844 24080 15896 24132
rect 18328 24191 18380 24200
rect 18328 24157 18337 24191
rect 18337 24157 18371 24191
rect 18371 24157 18380 24191
rect 18328 24148 18380 24157
rect 15660 24055 15712 24064
rect 15660 24021 15669 24055
rect 15669 24021 15703 24055
rect 15703 24021 15712 24055
rect 15660 24012 15712 24021
rect 18788 24012 18840 24064
rect 20076 24055 20128 24064
rect 20076 24021 20085 24055
rect 20085 24021 20119 24055
rect 20119 24021 20128 24055
rect 20076 24012 20128 24021
rect 24584 24225 24593 24259
rect 24593 24225 24627 24259
rect 24627 24225 24636 24259
rect 24584 24216 24636 24225
rect 24768 24259 24820 24268
rect 24768 24225 24777 24259
rect 24777 24225 24811 24259
rect 24811 24225 24820 24259
rect 24768 24216 24820 24225
rect 37740 24259 37792 24268
rect 37740 24225 37749 24259
rect 37749 24225 37783 24259
rect 37783 24225 37792 24259
rect 37740 24216 37792 24225
rect 37464 24191 37516 24200
rect 37464 24157 37473 24191
rect 37473 24157 37507 24191
rect 37507 24157 37516 24191
rect 37464 24148 37516 24157
rect 30472 24080 30524 24132
rect 23480 24012 23532 24064
rect 24308 24012 24360 24064
rect 24768 24012 24820 24064
rect 27988 24012 28040 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 1860 23808 1912 23860
rect 15844 23808 15896 23860
rect 20720 23851 20772 23860
rect 20720 23817 20729 23851
rect 20729 23817 20763 23851
rect 20763 23817 20772 23851
rect 20720 23808 20772 23817
rect 22836 23808 22888 23860
rect 30472 23851 30524 23860
rect 12992 23783 13044 23792
rect 12992 23749 13001 23783
rect 13001 23749 13035 23783
rect 13035 23749 13044 23783
rect 12992 23740 13044 23749
rect 2136 23715 2188 23724
rect 2136 23681 2145 23715
rect 2145 23681 2179 23715
rect 2179 23681 2188 23715
rect 2136 23672 2188 23681
rect 7012 23672 7064 23724
rect 10048 23672 10100 23724
rect 10416 23672 10468 23724
rect 4068 23536 4120 23588
rect 13084 23604 13136 23656
rect 14924 23672 14976 23724
rect 16856 23715 16908 23724
rect 16856 23681 16865 23715
rect 16865 23681 16899 23715
rect 16899 23681 16908 23715
rect 16856 23672 16908 23681
rect 21640 23740 21692 23792
rect 21916 23740 21968 23792
rect 22192 23783 22244 23792
rect 22192 23749 22201 23783
rect 22201 23749 22235 23783
rect 22235 23749 22244 23783
rect 22192 23740 22244 23749
rect 23388 23783 23440 23792
rect 23388 23749 23397 23783
rect 23397 23749 23431 23783
rect 23431 23749 23440 23783
rect 23388 23740 23440 23749
rect 30472 23817 30481 23851
rect 30481 23817 30515 23851
rect 30515 23817 30524 23851
rect 30472 23808 30524 23817
rect 38016 23740 38068 23792
rect 18604 23715 18656 23724
rect 18604 23681 18613 23715
rect 18613 23681 18647 23715
rect 18647 23681 18656 23715
rect 18604 23672 18656 23681
rect 18788 23715 18840 23724
rect 18788 23681 18797 23715
rect 18797 23681 18831 23715
rect 18831 23681 18840 23715
rect 18788 23672 18840 23681
rect 20076 23715 20128 23724
rect 20076 23681 20085 23715
rect 20085 23681 20119 23715
rect 20119 23681 20128 23715
rect 20076 23672 20128 23681
rect 20352 23672 20404 23724
rect 24584 23672 24636 23724
rect 27988 23672 28040 23724
rect 15292 23647 15344 23656
rect 15292 23613 15301 23647
rect 15301 23613 15335 23647
rect 15335 23613 15344 23647
rect 15292 23604 15344 23613
rect 22100 23647 22152 23656
rect 13452 23579 13504 23588
rect 13452 23545 13461 23579
rect 13461 23545 13495 23579
rect 13495 23545 13504 23579
rect 13452 23536 13504 23545
rect 14188 23536 14240 23588
rect 15108 23536 15160 23588
rect 22100 23613 22109 23647
rect 22109 23613 22143 23647
rect 22143 23613 22152 23647
rect 22100 23604 22152 23613
rect 22376 23647 22428 23656
rect 22376 23613 22385 23647
rect 22385 23613 22419 23647
rect 22419 23613 22428 23647
rect 22376 23604 22428 23613
rect 23480 23604 23532 23656
rect 34612 23672 34664 23724
rect 37924 23604 37976 23656
rect 24676 23536 24728 23588
rect 1952 23511 2004 23520
rect 1952 23477 1961 23511
rect 1961 23477 1995 23511
rect 1995 23477 2004 23511
rect 1952 23468 2004 23477
rect 9864 23468 9916 23520
rect 11520 23468 11572 23520
rect 14832 23468 14884 23520
rect 15292 23468 15344 23520
rect 15568 23468 15620 23520
rect 17040 23468 17092 23520
rect 18328 23468 18380 23520
rect 20812 23468 20864 23520
rect 27160 23536 27212 23588
rect 25136 23468 25188 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 23388 23264 23440 23316
rect 29552 23264 29604 23316
rect 10232 23171 10284 23180
rect 10232 23137 10241 23171
rect 10241 23137 10275 23171
rect 10275 23137 10284 23171
rect 10232 23128 10284 23137
rect 13360 23128 13412 23180
rect 13452 23128 13504 23180
rect 17040 23128 17092 23180
rect 18972 23128 19024 23180
rect 24676 23196 24728 23248
rect 23296 23128 23348 23180
rect 11888 23060 11940 23112
rect 13912 23060 13964 23112
rect 15844 23103 15896 23112
rect 15844 23069 15853 23103
rect 15853 23069 15887 23103
rect 15887 23069 15896 23103
rect 15844 23060 15896 23069
rect 16488 23060 16540 23112
rect 10324 23035 10376 23044
rect 10324 23001 10333 23035
rect 10333 23001 10367 23035
rect 10367 23001 10376 23035
rect 10324 22992 10376 23001
rect 9772 22924 9824 22976
rect 12348 22967 12400 22976
rect 12348 22933 12357 22967
rect 12357 22933 12391 22967
rect 12391 22933 12400 22967
rect 12348 22924 12400 22933
rect 14832 23035 14884 23044
rect 14832 23001 14841 23035
rect 14841 23001 14875 23035
rect 14875 23001 14884 23035
rect 14832 22992 14884 23001
rect 15752 22992 15804 23044
rect 16028 22992 16080 23044
rect 15660 22924 15712 22976
rect 19432 22924 19484 22976
rect 20352 22924 20404 22976
rect 21180 23035 21232 23044
rect 21180 23001 21189 23035
rect 21189 23001 21223 23035
rect 21223 23001 21232 23035
rect 21180 22992 21232 23001
rect 21364 22992 21416 23044
rect 25044 22992 25096 23044
rect 21916 22924 21968 22976
rect 22376 22924 22428 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 2044 22720 2096 22772
rect 1768 22627 1820 22636
rect 1768 22593 1777 22627
rect 1777 22593 1811 22627
rect 1811 22593 1820 22627
rect 1768 22584 1820 22593
rect 9772 22695 9824 22704
rect 9772 22661 9781 22695
rect 9781 22661 9815 22695
rect 9815 22661 9824 22695
rect 9772 22652 9824 22661
rect 9864 22695 9916 22704
rect 9864 22661 9873 22695
rect 9873 22661 9907 22695
rect 9907 22661 9916 22695
rect 12992 22720 13044 22772
rect 14648 22720 14700 22772
rect 20352 22763 20404 22772
rect 20352 22729 20361 22763
rect 20361 22729 20395 22763
rect 20395 22729 20404 22763
rect 20352 22720 20404 22729
rect 22192 22720 22244 22772
rect 25044 22763 25096 22772
rect 25044 22729 25053 22763
rect 25053 22729 25087 22763
rect 25087 22729 25096 22763
rect 25044 22720 25096 22729
rect 32404 22720 32456 22772
rect 9864 22652 9916 22661
rect 12440 22652 12492 22704
rect 13360 22652 13412 22704
rect 14372 22652 14424 22704
rect 17224 22695 17276 22704
rect 17224 22661 17233 22695
rect 17233 22661 17267 22695
rect 17267 22661 17276 22695
rect 17224 22652 17276 22661
rect 19432 22652 19484 22704
rect 24860 22652 24912 22704
rect 27252 22695 27304 22704
rect 27252 22661 27261 22695
rect 27261 22661 27295 22695
rect 27295 22661 27304 22695
rect 27252 22652 27304 22661
rect 27344 22695 27396 22704
rect 27344 22661 27353 22695
rect 27353 22661 27387 22695
rect 27387 22661 27396 22695
rect 27344 22652 27396 22661
rect 10876 22627 10928 22636
rect 7564 22516 7616 22568
rect 8576 22448 8628 22500
rect 10876 22593 10885 22627
rect 10885 22593 10919 22627
rect 10919 22593 10928 22627
rect 10876 22584 10928 22593
rect 14740 22627 14792 22636
rect 14740 22593 14749 22627
rect 14749 22593 14783 22627
rect 14783 22593 14792 22627
rect 14740 22584 14792 22593
rect 14924 22584 14976 22636
rect 18604 22627 18656 22636
rect 18604 22593 18613 22627
rect 18613 22593 18647 22627
rect 18647 22593 18656 22627
rect 18604 22584 18656 22593
rect 25044 22584 25096 22636
rect 30932 22627 30984 22636
rect 11612 22516 11664 22568
rect 11704 22448 11756 22500
rect 13728 22516 13780 22568
rect 14556 22559 14608 22568
rect 14556 22525 14565 22559
rect 14565 22525 14599 22559
rect 14599 22525 14608 22559
rect 14556 22516 14608 22525
rect 16212 22516 16264 22568
rect 17960 22559 18012 22568
rect 17960 22525 17969 22559
rect 17969 22525 18003 22559
rect 18003 22525 18012 22559
rect 17960 22516 18012 22525
rect 19248 22516 19300 22568
rect 21364 22516 21416 22568
rect 24768 22516 24820 22568
rect 30932 22593 30941 22627
rect 30941 22593 30975 22627
rect 30975 22593 30984 22627
rect 30932 22584 30984 22593
rect 38016 22627 38068 22636
rect 38016 22593 38025 22627
rect 38025 22593 38059 22627
rect 38059 22593 38068 22627
rect 38016 22584 38068 22593
rect 26884 22516 26936 22568
rect 16120 22448 16172 22500
rect 16488 22448 16540 22500
rect 38200 22491 38252 22500
rect 38200 22457 38209 22491
rect 38209 22457 38243 22491
rect 38243 22457 38252 22491
rect 38200 22448 38252 22457
rect 8300 22380 8352 22432
rect 10140 22380 10192 22432
rect 16580 22380 16632 22432
rect 17960 22380 18012 22432
rect 27068 22380 27120 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 8852 22176 8904 22228
rect 10048 22176 10100 22228
rect 10876 22176 10928 22228
rect 8208 22108 8260 22160
rect 13728 22108 13780 22160
rect 7012 22083 7064 22092
rect 7012 22049 7021 22083
rect 7021 22049 7055 22083
rect 7055 22049 7064 22083
rect 7012 22040 7064 22049
rect 11612 22040 11664 22092
rect 14372 22083 14424 22092
rect 14372 22049 14381 22083
rect 14381 22049 14415 22083
rect 14415 22049 14424 22083
rect 14372 22040 14424 22049
rect 7104 21972 7156 22024
rect 8300 21972 8352 22024
rect 14004 21972 14056 22024
rect 16028 22108 16080 22160
rect 17224 22108 17276 22160
rect 19708 22176 19760 22228
rect 27344 22176 27396 22228
rect 17868 22108 17920 22160
rect 9036 21904 9088 21956
rect 10140 21947 10192 21956
rect 10140 21913 10149 21947
rect 10149 21913 10183 21947
rect 10183 21913 10192 21947
rect 10140 21904 10192 21913
rect 7472 21836 7524 21888
rect 10876 21904 10928 21956
rect 11520 21947 11572 21956
rect 11520 21913 11529 21947
rect 11529 21913 11563 21947
rect 11563 21913 11572 21947
rect 11520 21904 11572 21913
rect 12532 21904 12584 21956
rect 17960 22083 18012 22092
rect 17960 22049 17969 22083
rect 17969 22049 18003 22083
rect 18003 22049 18012 22083
rect 17960 22040 18012 22049
rect 25044 22108 25096 22160
rect 25412 22108 25464 22160
rect 27528 22151 27580 22160
rect 27528 22117 27537 22151
rect 27537 22117 27571 22151
rect 27571 22117 27580 22151
rect 27528 22108 27580 22117
rect 15384 22015 15436 22024
rect 15384 21981 15393 22015
rect 15393 21981 15427 22015
rect 15427 21981 15436 22015
rect 15384 21972 15436 21981
rect 15844 22015 15896 22024
rect 15844 21981 15853 22015
rect 15853 21981 15887 22015
rect 15887 21981 15896 22015
rect 15844 21972 15896 21981
rect 15200 21947 15252 21956
rect 15200 21913 15209 21947
rect 15209 21913 15243 21947
rect 15243 21913 15252 21947
rect 15200 21904 15252 21913
rect 16120 21972 16172 22024
rect 16488 21972 16540 22024
rect 16856 22015 16908 22024
rect 16856 21981 16865 22015
rect 16865 21981 16899 22015
rect 16899 21981 16908 22015
rect 16856 21972 16908 21981
rect 20260 22040 20312 22092
rect 28264 22040 28316 22092
rect 20904 21972 20956 22024
rect 34796 21972 34848 22024
rect 12992 21836 13044 21888
rect 13176 21836 13228 21888
rect 16120 21836 16172 21888
rect 17776 21904 17828 21956
rect 22376 21904 22428 21956
rect 22836 21904 22888 21956
rect 26976 21947 27028 21956
rect 26976 21913 26985 21947
rect 26985 21913 27019 21947
rect 27019 21913 27028 21947
rect 26976 21904 27028 21913
rect 27068 21947 27120 21956
rect 27068 21913 27077 21947
rect 27077 21913 27111 21947
rect 27111 21913 27120 21947
rect 27068 21904 27120 21913
rect 19432 21836 19484 21888
rect 19708 21836 19760 21888
rect 23480 21836 23532 21888
rect 23572 21836 23624 21888
rect 38200 21879 38252 21888
rect 38200 21845 38209 21879
rect 38209 21845 38243 21879
rect 38243 21845 38252 21879
rect 38200 21836 38252 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 8576 21675 8628 21684
rect 8576 21641 8585 21675
rect 8585 21641 8619 21675
rect 8619 21641 8628 21675
rect 8576 21632 8628 21641
rect 8760 21632 8812 21684
rect 6736 21564 6788 21616
rect 7380 21607 7432 21616
rect 7380 21573 7389 21607
rect 7389 21573 7423 21607
rect 7423 21573 7432 21607
rect 7380 21564 7432 21573
rect 7472 21607 7524 21616
rect 7472 21573 7481 21607
rect 7481 21573 7515 21607
rect 7515 21573 7524 21607
rect 7472 21564 7524 21573
rect 1676 21539 1728 21548
rect 1676 21505 1685 21539
rect 1685 21505 1719 21539
rect 1719 21505 1728 21539
rect 1676 21496 1728 21505
rect 7104 21496 7156 21548
rect 10692 21564 10744 21616
rect 12808 21607 12860 21616
rect 12808 21573 12817 21607
rect 12817 21573 12851 21607
rect 12851 21573 12860 21607
rect 12808 21564 12860 21573
rect 11612 21496 11664 21548
rect 15200 21632 15252 21684
rect 14556 21564 14608 21616
rect 16028 21632 16080 21684
rect 15936 21564 15988 21616
rect 17500 21564 17552 21616
rect 17868 21564 17920 21616
rect 5632 21428 5684 21480
rect 6920 21360 6972 21412
rect 8208 21360 8260 21412
rect 8392 21292 8444 21344
rect 9956 21428 10008 21480
rect 9404 21360 9456 21412
rect 12532 21360 12584 21412
rect 13176 21428 13228 21480
rect 13452 21428 13504 21480
rect 15568 21428 15620 21480
rect 13728 21360 13780 21412
rect 16488 21428 16540 21480
rect 18420 21607 18472 21616
rect 18420 21573 18429 21607
rect 18429 21573 18463 21607
rect 18463 21573 18472 21607
rect 18420 21564 18472 21573
rect 18972 21607 19024 21616
rect 18972 21573 18981 21607
rect 18981 21573 19015 21607
rect 19015 21573 19024 21607
rect 18972 21564 19024 21573
rect 19432 21632 19484 21684
rect 19524 21564 19576 21616
rect 28264 21675 28316 21684
rect 23572 21607 23624 21616
rect 23572 21573 23581 21607
rect 23581 21573 23615 21607
rect 23615 21573 23624 21607
rect 23572 21564 23624 21573
rect 20904 21496 20956 21548
rect 21088 21496 21140 21548
rect 28264 21641 28273 21675
rect 28273 21641 28307 21675
rect 28307 21641 28316 21675
rect 28264 21632 28316 21641
rect 18328 21471 18380 21480
rect 18328 21437 18337 21471
rect 18337 21437 18371 21471
rect 18371 21437 18380 21471
rect 18328 21428 18380 21437
rect 18512 21428 18564 21480
rect 19616 21428 19668 21480
rect 15752 21360 15804 21412
rect 14372 21292 14424 21344
rect 17408 21292 17460 21344
rect 17684 21335 17736 21344
rect 17684 21301 17693 21335
rect 17693 21301 17727 21335
rect 17727 21301 17736 21335
rect 17684 21292 17736 21301
rect 17960 21292 18012 21344
rect 20996 21360 21048 21412
rect 23296 21428 23348 21480
rect 37372 21564 37424 21616
rect 37740 21496 37792 21548
rect 20444 21292 20496 21344
rect 22836 21292 22888 21344
rect 24768 21292 24820 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 2228 21088 2280 21140
rect 15936 21088 15988 21140
rect 9036 21020 9088 21072
rect 13544 21020 13596 21072
rect 15384 21020 15436 21072
rect 4804 20995 4856 21004
rect 4804 20961 4813 20995
rect 4813 20961 4847 20995
rect 4847 20961 4856 20995
rect 4804 20952 4856 20961
rect 5632 20995 5684 21004
rect 5632 20961 5641 20995
rect 5641 20961 5675 20995
rect 5675 20961 5684 20995
rect 5632 20952 5684 20961
rect 9956 20952 10008 21004
rect 11336 20952 11388 21004
rect 12256 20995 12308 21004
rect 12256 20961 12265 20995
rect 12265 20961 12299 20995
rect 12299 20961 12308 20995
rect 12256 20952 12308 20961
rect 13268 20995 13320 21004
rect 13268 20961 13277 20995
rect 13277 20961 13311 20995
rect 13311 20961 13320 20995
rect 18052 21088 18104 21140
rect 13268 20952 13320 20961
rect 18144 21020 18196 21072
rect 16948 20995 17000 21004
rect 16948 20961 16957 20995
rect 16957 20961 16991 20995
rect 16991 20961 17000 20995
rect 22744 21088 22796 21140
rect 18604 21020 18656 21072
rect 28540 21088 28592 21140
rect 38016 21088 38068 21140
rect 22928 21020 22980 21072
rect 23572 21020 23624 21072
rect 23756 21063 23808 21072
rect 23756 21029 23765 21063
rect 23765 21029 23799 21063
rect 23799 21029 23808 21063
rect 23756 21020 23808 21029
rect 16948 20952 17000 20961
rect 18972 20952 19024 21004
rect 19616 20995 19668 21004
rect 19616 20961 19625 20995
rect 19625 20961 19659 20995
rect 19659 20961 19668 20995
rect 19616 20952 19668 20961
rect 21272 20952 21324 21004
rect 25780 20952 25832 21004
rect 1584 20927 1636 20936
rect 1584 20893 1593 20927
rect 1593 20893 1627 20927
rect 1627 20893 1636 20927
rect 1584 20884 1636 20893
rect 1860 20927 1912 20936
rect 1860 20893 1869 20927
rect 1869 20893 1903 20927
rect 1903 20893 1912 20927
rect 1860 20884 1912 20893
rect 7472 20884 7524 20936
rect 9312 20884 9364 20936
rect 4528 20859 4580 20868
rect 4528 20825 4537 20859
rect 4537 20825 4571 20859
rect 4571 20825 4580 20859
rect 4528 20816 4580 20825
rect 7748 20816 7800 20868
rect 8668 20816 8720 20868
rect 10140 20859 10192 20868
rect 10140 20825 10149 20859
rect 10149 20825 10183 20859
rect 10183 20825 10192 20859
rect 10140 20816 10192 20825
rect 12348 20859 12400 20868
rect 8484 20791 8536 20800
rect 8484 20757 8493 20791
rect 8493 20757 8527 20791
rect 8527 20757 8536 20791
rect 8484 20748 8536 20757
rect 9220 20791 9272 20800
rect 9220 20757 9229 20791
rect 9229 20757 9263 20791
rect 9263 20757 9272 20791
rect 9220 20748 9272 20757
rect 9956 20748 10008 20800
rect 12348 20825 12357 20859
rect 12357 20825 12391 20859
rect 12391 20825 12400 20859
rect 12348 20816 12400 20825
rect 10692 20748 10744 20800
rect 12624 20816 12676 20868
rect 13728 20884 13780 20936
rect 19524 20884 19576 20936
rect 20076 20884 20128 20936
rect 20996 20927 21048 20936
rect 20996 20893 21005 20927
rect 21005 20893 21039 20927
rect 21039 20893 21048 20927
rect 22468 20927 22520 20936
rect 20996 20884 21048 20893
rect 22468 20893 22477 20927
rect 22477 20893 22511 20927
rect 22511 20893 22520 20927
rect 22468 20884 22520 20893
rect 22560 20927 22612 20936
rect 22560 20893 22569 20927
rect 22569 20893 22603 20927
rect 22603 20893 22612 20927
rect 25228 20927 25280 20936
rect 22560 20884 22612 20893
rect 25228 20893 25237 20927
rect 25237 20893 25271 20927
rect 25271 20893 25280 20927
rect 25228 20884 25280 20893
rect 38384 20884 38436 20936
rect 14648 20859 14700 20868
rect 14648 20825 14657 20859
rect 14657 20825 14691 20859
rect 14691 20825 14700 20859
rect 14648 20816 14700 20825
rect 14740 20859 14792 20868
rect 14740 20825 14749 20859
rect 14749 20825 14783 20859
rect 14783 20825 14792 20859
rect 14740 20816 14792 20825
rect 15936 20816 15988 20868
rect 16580 20748 16632 20800
rect 17776 20816 17828 20868
rect 18328 20859 18380 20868
rect 18328 20825 18337 20859
rect 18337 20825 18371 20859
rect 18371 20825 18380 20859
rect 18328 20816 18380 20825
rect 20444 20859 20496 20868
rect 20444 20825 20453 20859
rect 20453 20825 20487 20859
rect 20487 20825 20496 20859
rect 20444 20816 20496 20825
rect 22928 20816 22980 20868
rect 17684 20748 17736 20800
rect 25044 20791 25096 20800
rect 25044 20757 25053 20791
rect 25053 20757 25087 20791
rect 25087 20757 25096 20791
rect 25044 20748 25096 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 6736 20544 6788 20596
rect 7932 20544 7984 20596
rect 8852 20544 8904 20596
rect 10232 20544 10284 20596
rect 12256 20544 12308 20596
rect 14096 20544 14148 20596
rect 14740 20544 14792 20596
rect 1860 20476 1912 20528
rect 8116 20476 8168 20528
rect 9220 20476 9272 20528
rect 10784 20476 10836 20528
rect 10968 20476 11020 20528
rect 13268 20519 13320 20528
rect 13268 20485 13277 20519
rect 13277 20485 13311 20519
rect 13311 20485 13320 20519
rect 13268 20476 13320 20485
rect 16856 20544 16908 20596
rect 15292 20476 15344 20528
rect 15936 20476 15988 20528
rect 16580 20476 16632 20528
rect 7656 20451 7708 20460
rect 7656 20417 7665 20451
rect 7665 20417 7699 20451
rect 7699 20417 7708 20451
rect 7656 20408 7708 20417
rect 14280 20451 14332 20460
rect 14280 20417 14289 20451
rect 14289 20417 14323 20451
rect 14323 20417 14332 20451
rect 14280 20408 14332 20417
rect 9220 20383 9272 20392
rect 9220 20349 9229 20383
rect 9229 20349 9263 20383
rect 9263 20349 9272 20383
rect 9220 20340 9272 20349
rect 9588 20340 9640 20392
rect 11520 20340 11572 20392
rect 11796 20383 11848 20392
rect 11796 20349 11805 20383
rect 11805 20349 11839 20383
rect 11839 20349 11848 20383
rect 11796 20340 11848 20349
rect 13176 20383 13228 20392
rect 7104 20272 7156 20324
rect 13176 20349 13185 20383
rect 13185 20349 13219 20383
rect 13219 20349 13228 20383
rect 13176 20340 13228 20349
rect 13452 20383 13504 20392
rect 13452 20349 13461 20383
rect 13461 20349 13495 20383
rect 13495 20349 13504 20383
rect 13452 20340 13504 20349
rect 13820 20340 13872 20392
rect 15476 20340 15528 20392
rect 19248 20544 19300 20596
rect 25136 20544 25188 20596
rect 26976 20544 27028 20596
rect 17316 20519 17368 20528
rect 17316 20485 17325 20519
rect 17325 20485 17359 20519
rect 17359 20485 17368 20519
rect 17316 20476 17368 20485
rect 18144 20476 18196 20528
rect 19340 20519 19392 20528
rect 19340 20485 19349 20519
rect 19349 20485 19383 20519
rect 19383 20485 19392 20519
rect 19340 20476 19392 20485
rect 19892 20476 19944 20528
rect 21364 20476 21416 20528
rect 23020 20476 23072 20528
rect 24400 20451 24452 20460
rect 17592 20340 17644 20392
rect 24400 20417 24409 20451
rect 24409 20417 24443 20451
rect 24443 20417 24452 20451
rect 24400 20408 24452 20417
rect 25044 20408 25096 20460
rect 25780 20451 25832 20460
rect 25780 20417 25789 20451
rect 25789 20417 25823 20451
rect 25823 20417 25832 20451
rect 25780 20408 25832 20417
rect 27160 20451 27212 20460
rect 27160 20417 27169 20451
rect 27169 20417 27203 20451
rect 27203 20417 27212 20451
rect 27160 20408 27212 20417
rect 38292 20451 38344 20460
rect 38292 20417 38301 20451
rect 38301 20417 38335 20451
rect 38335 20417 38344 20451
rect 38292 20408 38344 20417
rect 19984 20340 20036 20392
rect 20168 20383 20220 20392
rect 20168 20349 20177 20383
rect 20177 20349 20211 20383
rect 20211 20349 20220 20383
rect 20168 20340 20220 20349
rect 20996 20340 21048 20392
rect 21640 20340 21692 20392
rect 17776 20315 17828 20324
rect 17776 20281 17785 20315
rect 17785 20281 17819 20315
rect 17819 20281 17828 20315
rect 17776 20272 17828 20281
rect 18144 20272 18196 20324
rect 22560 20340 22612 20392
rect 23296 20383 23348 20392
rect 23296 20349 23305 20383
rect 23305 20349 23339 20383
rect 23339 20349 23348 20383
rect 23296 20340 23348 20349
rect 26792 20272 26844 20324
rect 17132 20204 17184 20256
rect 21548 20204 21600 20256
rect 25136 20204 25188 20256
rect 34704 20204 34756 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 9956 20000 10008 20052
rect 10784 20043 10836 20052
rect 10784 20009 10793 20043
rect 10793 20009 10827 20043
rect 10827 20009 10836 20043
rect 10784 20000 10836 20009
rect 11796 20000 11848 20052
rect 17224 20000 17276 20052
rect 7104 19932 7156 19984
rect 7656 19932 7708 19984
rect 11336 19932 11388 19984
rect 22284 20000 22336 20052
rect 23388 20000 23440 20052
rect 25228 20000 25280 20052
rect 8944 19796 8996 19848
rect 9772 19839 9824 19848
rect 9772 19805 9781 19839
rect 9781 19805 9815 19839
rect 9815 19805 9824 19839
rect 9772 19796 9824 19805
rect 10692 19839 10744 19848
rect 10692 19805 10701 19839
rect 10701 19805 10735 19839
rect 10735 19805 10744 19839
rect 10692 19796 10744 19805
rect 11612 19796 11664 19848
rect 14096 19864 14148 19916
rect 19340 19864 19392 19916
rect 3976 19728 4028 19780
rect 5080 19728 5132 19780
rect 6736 19728 6788 19780
rect 8484 19728 8536 19780
rect 8576 19771 8628 19780
rect 8576 19737 8585 19771
rect 8585 19737 8619 19771
rect 8619 19737 8628 19771
rect 8576 19728 8628 19737
rect 10140 19728 10192 19780
rect 11060 19728 11112 19780
rect 12256 19728 12308 19780
rect 12532 19771 12584 19780
rect 12532 19737 12541 19771
rect 12541 19737 12575 19771
rect 12575 19737 12584 19771
rect 13452 19771 13504 19780
rect 12532 19728 12584 19737
rect 13452 19737 13461 19771
rect 13461 19737 13495 19771
rect 13495 19737 13504 19771
rect 13452 19728 13504 19737
rect 14464 19771 14516 19780
rect 14464 19737 14473 19771
rect 14473 19737 14507 19771
rect 14507 19737 14516 19771
rect 14464 19728 14516 19737
rect 16120 19728 16172 19780
rect 8208 19660 8260 19712
rect 10048 19660 10100 19712
rect 10232 19660 10284 19712
rect 10968 19660 11020 19712
rect 12900 19660 12952 19712
rect 13544 19660 13596 19712
rect 17408 19796 17460 19848
rect 22744 19932 22796 19984
rect 19892 19907 19944 19916
rect 19892 19873 19901 19907
rect 19901 19873 19935 19907
rect 19935 19873 19944 19907
rect 21272 19907 21324 19916
rect 19892 19864 19944 19873
rect 21272 19873 21281 19907
rect 21281 19873 21315 19907
rect 21315 19873 21324 19907
rect 21272 19864 21324 19873
rect 22100 19864 22152 19916
rect 22284 19907 22336 19916
rect 22284 19873 22293 19907
rect 22293 19873 22327 19907
rect 22327 19873 22336 19907
rect 22284 19864 22336 19873
rect 24952 19864 25004 19916
rect 17040 19660 17092 19712
rect 17684 19771 17736 19780
rect 17684 19737 17693 19771
rect 17693 19737 17727 19771
rect 17727 19737 17736 19771
rect 18604 19771 18656 19780
rect 17684 19728 17736 19737
rect 18604 19737 18613 19771
rect 18613 19737 18647 19771
rect 18647 19737 18656 19771
rect 18604 19728 18656 19737
rect 19340 19728 19392 19780
rect 20168 19728 20220 19780
rect 21640 19728 21692 19780
rect 24492 19796 24544 19848
rect 24676 19796 24728 19848
rect 25136 19975 25188 19984
rect 25136 19941 25145 19975
rect 25145 19941 25179 19975
rect 25179 19941 25188 19975
rect 25136 19932 25188 19941
rect 27620 19932 27672 19984
rect 25412 19864 25464 19916
rect 26700 19796 26752 19848
rect 28632 19796 28684 19848
rect 25504 19728 25556 19780
rect 37832 19728 37884 19780
rect 21548 19660 21600 19712
rect 25320 19660 25372 19712
rect 26516 19660 26568 19712
rect 29920 19660 29972 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 1492 19456 1544 19508
rect 5080 19499 5132 19508
rect 5080 19465 5089 19499
rect 5089 19465 5123 19499
rect 5123 19465 5132 19499
rect 5080 19456 5132 19465
rect 6736 19456 6788 19508
rect 7840 19388 7892 19440
rect 1860 19320 1912 19372
rect 5632 19363 5684 19372
rect 5632 19329 5641 19363
rect 5641 19329 5675 19363
rect 5675 19329 5684 19363
rect 8116 19456 8168 19508
rect 8392 19431 8444 19440
rect 8392 19397 8401 19431
rect 8401 19397 8435 19431
rect 8435 19397 8444 19431
rect 8392 19388 8444 19397
rect 8576 19388 8628 19440
rect 9404 19388 9456 19440
rect 13268 19456 13320 19508
rect 15108 19456 15160 19508
rect 15292 19499 15344 19508
rect 15292 19465 15301 19499
rect 15301 19465 15335 19499
rect 15335 19465 15344 19499
rect 15292 19456 15344 19465
rect 16212 19456 16264 19508
rect 17408 19456 17460 19508
rect 12532 19388 12584 19440
rect 13084 19431 13136 19440
rect 13084 19397 13093 19431
rect 13093 19397 13127 19431
rect 13127 19397 13136 19431
rect 13084 19388 13136 19397
rect 13452 19388 13504 19440
rect 14372 19388 14424 19440
rect 16120 19388 16172 19440
rect 19432 19456 19484 19508
rect 23020 19499 23072 19508
rect 5632 19320 5684 19329
rect 5816 19252 5868 19304
rect 6920 19252 6972 19304
rect 7104 19295 7156 19304
rect 7104 19261 7113 19295
rect 7113 19261 7147 19295
rect 7147 19261 7156 19295
rect 7104 19252 7156 19261
rect 10876 19320 10928 19372
rect 4804 19184 4856 19236
rect 11244 19252 11296 19304
rect 12992 19295 13044 19304
rect 11060 19184 11112 19236
rect 12072 19184 12124 19236
rect 5724 19159 5776 19168
rect 5724 19125 5733 19159
rect 5733 19125 5767 19159
rect 5767 19125 5776 19159
rect 5724 19116 5776 19125
rect 11428 19116 11480 19168
rect 11796 19116 11848 19168
rect 12256 19116 12308 19168
rect 12992 19261 13001 19295
rect 13001 19261 13035 19295
rect 13035 19261 13044 19295
rect 12992 19252 13044 19261
rect 15752 19320 15804 19372
rect 15936 19363 15988 19372
rect 15936 19329 15945 19363
rect 15945 19329 15979 19363
rect 15979 19329 15988 19363
rect 15936 19320 15988 19329
rect 16488 19252 16540 19304
rect 17960 19320 18012 19372
rect 22560 19388 22612 19440
rect 23020 19465 23029 19499
rect 23029 19465 23063 19499
rect 23063 19465 23072 19499
rect 23020 19456 23072 19465
rect 24676 19499 24728 19508
rect 22928 19388 22980 19440
rect 18512 19320 18564 19372
rect 18236 19252 18288 19304
rect 21088 19320 21140 19372
rect 20628 19252 20680 19304
rect 21364 19363 21416 19372
rect 21364 19329 21373 19363
rect 21373 19329 21407 19363
rect 21407 19329 21416 19363
rect 21364 19320 21416 19329
rect 21732 19320 21784 19372
rect 24676 19465 24685 19499
rect 24685 19465 24719 19499
rect 24719 19465 24728 19499
rect 24676 19456 24728 19465
rect 25780 19456 25832 19508
rect 26976 19456 27028 19508
rect 28632 19499 28684 19508
rect 28632 19465 28641 19499
rect 28641 19465 28675 19499
rect 28675 19465 28684 19499
rect 28632 19456 28684 19465
rect 28724 19456 28776 19508
rect 24492 19320 24544 19372
rect 25504 19320 25556 19372
rect 26608 19320 26660 19372
rect 27160 19320 27212 19372
rect 28908 19320 28960 19372
rect 29092 19320 29144 19372
rect 30104 19363 30156 19372
rect 30104 19329 30113 19363
rect 30113 19329 30147 19363
rect 30147 19329 30156 19363
rect 30104 19320 30156 19329
rect 36912 19320 36964 19372
rect 26056 19295 26108 19304
rect 26056 19261 26065 19295
rect 26065 19261 26099 19295
rect 26099 19261 26108 19295
rect 26056 19252 26108 19261
rect 20444 19184 20496 19236
rect 24584 19184 24636 19236
rect 14372 19116 14424 19168
rect 14556 19116 14608 19168
rect 18144 19116 18196 19168
rect 18604 19116 18656 19168
rect 20536 19116 20588 19168
rect 27068 19116 27120 19168
rect 27528 19116 27580 19168
rect 29368 19159 29420 19168
rect 29368 19125 29377 19159
rect 29377 19125 29411 19159
rect 29411 19125 29420 19159
rect 29368 19116 29420 19125
rect 38200 19159 38252 19168
rect 38200 19125 38209 19159
rect 38209 19125 38243 19159
rect 38243 19125 38252 19159
rect 38200 19116 38252 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 7840 18955 7892 18964
rect 7840 18921 7849 18955
rect 7849 18921 7883 18955
rect 7883 18921 7892 18955
rect 7840 18912 7892 18921
rect 8208 18912 8260 18964
rect 13084 18912 13136 18964
rect 14372 18912 14424 18964
rect 17132 18912 17184 18964
rect 17684 18912 17736 18964
rect 20628 18955 20680 18964
rect 20628 18921 20637 18955
rect 20637 18921 20671 18955
rect 20671 18921 20680 18955
rect 20628 18912 20680 18921
rect 23848 18912 23900 18964
rect 1768 18751 1820 18760
rect 1768 18717 1777 18751
rect 1777 18717 1811 18751
rect 1811 18717 1820 18751
rect 1768 18708 1820 18717
rect 5816 18751 5868 18760
rect 5816 18717 5825 18751
rect 5825 18717 5859 18751
rect 5859 18717 5868 18751
rect 5816 18708 5868 18717
rect 8668 18776 8720 18828
rect 9772 18751 9824 18760
rect 5448 18572 5500 18624
rect 7012 18572 7064 18624
rect 7104 18572 7156 18624
rect 9772 18717 9781 18751
rect 9781 18717 9815 18751
rect 9815 18717 9824 18751
rect 9772 18708 9824 18717
rect 10140 18708 10192 18760
rect 12072 18776 12124 18828
rect 11244 18708 11296 18760
rect 11704 18751 11756 18760
rect 11704 18717 11713 18751
rect 11713 18717 11747 18751
rect 11747 18717 11756 18751
rect 11704 18708 11756 18717
rect 11796 18708 11848 18760
rect 12624 18844 12676 18896
rect 13728 18776 13780 18828
rect 16212 18776 16264 18828
rect 16672 18819 16724 18828
rect 16672 18785 16681 18819
rect 16681 18785 16715 18819
rect 16715 18785 16724 18819
rect 16672 18776 16724 18785
rect 26056 18912 26108 18964
rect 36912 18912 36964 18964
rect 25688 18844 25740 18896
rect 17132 18751 17184 18760
rect 17132 18717 17141 18751
rect 17141 18717 17175 18751
rect 17175 18717 17184 18751
rect 17132 18708 17184 18717
rect 9404 18640 9456 18692
rect 9036 18572 9088 18624
rect 9220 18615 9272 18624
rect 9220 18581 9229 18615
rect 9229 18581 9263 18615
rect 9263 18581 9272 18615
rect 9220 18572 9272 18581
rect 10508 18615 10560 18624
rect 10508 18581 10517 18615
rect 10517 18581 10551 18615
rect 10551 18581 10560 18615
rect 10508 18572 10560 18581
rect 10600 18572 10652 18624
rect 11980 18572 12032 18624
rect 12532 18683 12584 18692
rect 12532 18649 12541 18683
rect 12541 18649 12575 18683
rect 12575 18649 12584 18683
rect 12532 18640 12584 18649
rect 14556 18640 14608 18692
rect 14740 18683 14792 18692
rect 14740 18649 14749 18683
rect 14749 18649 14783 18683
rect 14783 18649 14792 18683
rect 14740 18640 14792 18649
rect 15476 18640 15528 18692
rect 16120 18683 16172 18692
rect 16120 18649 16129 18683
rect 16129 18649 16163 18683
rect 16163 18649 16172 18683
rect 16120 18640 16172 18649
rect 20260 18708 20312 18760
rect 22744 18708 22796 18760
rect 26608 18776 26660 18828
rect 27068 18776 27120 18828
rect 27528 18751 27580 18760
rect 24676 18683 24728 18692
rect 14924 18572 14976 18624
rect 24676 18649 24685 18683
rect 24685 18649 24719 18683
rect 24719 18649 24728 18683
rect 24676 18640 24728 18649
rect 25320 18640 25372 18692
rect 27528 18717 27537 18751
rect 27537 18717 27571 18751
rect 27571 18717 27580 18751
rect 27528 18708 27580 18717
rect 29000 18751 29052 18760
rect 29000 18717 29009 18751
rect 29009 18717 29043 18751
rect 29043 18717 29052 18751
rect 29000 18708 29052 18717
rect 38384 18844 38436 18896
rect 16488 18572 16540 18624
rect 25964 18572 26016 18624
rect 26516 18640 26568 18692
rect 26884 18683 26936 18692
rect 26884 18649 26893 18683
rect 26893 18649 26927 18683
rect 26927 18649 26936 18683
rect 26884 18640 26936 18649
rect 26976 18640 27028 18692
rect 34704 18708 34756 18760
rect 35164 18751 35216 18760
rect 35164 18717 35173 18751
rect 35173 18717 35207 18751
rect 35207 18717 35216 18751
rect 35164 18708 35216 18717
rect 30196 18572 30248 18624
rect 33600 18615 33652 18624
rect 33600 18581 33609 18615
rect 33609 18581 33643 18615
rect 33643 18581 33652 18615
rect 33600 18572 33652 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 8760 18368 8812 18420
rect 4620 18300 4672 18352
rect 4804 18343 4856 18352
rect 4804 18309 4813 18343
rect 4813 18309 4847 18343
rect 4847 18309 4856 18343
rect 4804 18300 4856 18309
rect 5448 18343 5500 18352
rect 5448 18309 5457 18343
rect 5457 18309 5491 18343
rect 5491 18309 5500 18343
rect 5448 18300 5500 18309
rect 6644 18300 6696 18352
rect 7932 18300 7984 18352
rect 8668 18232 8720 18284
rect 11796 18368 11848 18420
rect 11980 18368 12032 18420
rect 12440 18368 12492 18420
rect 13452 18368 13504 18420
rect 14464 18368 14516 18420
rect 10508 18300 10560 18352
rect 9956 18232 10008 18284
rect 10324 18275 10376 18284
rect 10324 18241 10333 18275
rect 10333 18241 10367 18275
rect 10367 18241 10376 18275
rect 10324 18232 10376 18241
rect 11336 18232 11388 18284
rect 14648 18300 14700 18352
rect 17040 18343 17092 18352
rect 17040 18309 17049 18343
rect 17049 18309 17083 18343
rect 17083 18309 17092 18343
rect 17040 18300 17092 18309
rect 18328 18368 18380 18420
rect 18420 18368 18472 18420
rect 20260 18368 20312 18420
rect 20352 18300 20404 18352
rect 22376 18300 22428 18352
rect 23572 18300 23624 18352
rect 27804 18343 27856 18352
rect 27804 18309 27813 18343
rect 27813 18309 27847 18343
rect 27847 18309 27856 18343
rect 27804 18300 27856 18309
rect 29368 18300 29420 18352
rect 30104 18368 30156 18420
rect 35164 18368 35216 18420
rect 35348 18300 35400 18352
rect 14188 18232 14240 18284
rect 18052 18275 18104 18284
rect 18052 18241 18061 18275
rect 18061 18241 18095 18275
rect 18095 18241 18104 18275
rect 18052 18232 18104 18241
rect 18788 18232 18840 18284
rect 20536 18275 20588 18284
rect 20536 18241 20545 18275
rect 20545 18241 20579 18275
rect 20579 18241 20588 18275
rect 20536 18232 20588 18241
rect 23664 18232 23716 18284
rect 24768 18232 24820 18284
rect 28908 18275 28960 18284
rect 28908 18241 28917 18275
rect 28917 18241 28951 18275
rect 28951 18241 28960 18275
rect 28908 18232 28960 18241
rect 29000 18232 29052 18284
rect 30196 18275 30248 18284
rect 30196 18241 30205 18275
rect 30205 18241 30239 18275
rect 30239 18241 30248 18275
rect 30196 18232 30248 18241
rect 1584 18207 1636 18216
rect 1584 18173 1593 18207
rect 1593 18173 1627 18207
rect 1627 18173 1636 18207
rect 1584 18164 1636 18173
rect 5724 18164 5776 18216
rect 6920 18164 6972 18216
rect 8576 18164 8628 18216
rect 10600 18164 10652 18216
rect 11520 18164 11572 18216
rect 12072 18164 12124 18216
rect 13176 18164 13228 18216
rect 13728 18164 13780 18216
rect 15200 18164 15252 18216
rect 15384 18207 15436 18216
rect 15384 18173 15393 18207
rect 15393 18173 15427 18207
rect 15427 18173 15436 18207
rect 15384 18164 15436 18173
rect 15844 18164 15896 18216
rect 16212 18164 16264 18216
rect 9680 18096 9732 18148
rect 9588 18028 9640 18080
rect 12808 18028 12860 18080
rect 16120 18096 16172 18148
rect 14648 18028 14700 18080
rect 14740 18028 14792 18080
rect 23388 18164 23440 18216
rect 24676 18164 24728 18216
rect 25688 18164 25740 18216
rect 27988 18096 28040 18148
rect 21088 18028 21140 18080
rect 26976 18028 27028 18080
rect 28540 18028 28592 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 4620 17824 4672 17876
rect 5172 17824 5224 17876
rect 10232 17756 10284 17808
rect 10324 17756 10376 17808
rect 11980 17756 12032 17808
rect 1860 17688 1912 17740
rect 4252 17663 4304 17672
rect 4252 17629 4261 17663
rect 4261 17629 4295 17663
rect 4295 17629 4304 17663
rect 4252 17620 4304 17629
rect 5448 17620 5500 17672
rect 10784 17688 10836 17740
rect 11428 17688 11480 17740
rect 8668 17620 8720 17672
rect 10324 17620 10376 17672
rect 10600 17663 10652 17672
rect 10600 17629 10609 17663
rect 10609 17629 10643 17663
rect 10643 17629 10652 17663
rect 10600 17620 10652 17629
rect 13728 17824 13780 17876
rect 14096 17688 14148 17740
rect 15200 17731 15252 17740
rect 15200 17697 15209 17731
rect 15209 17697 15243 17731
rect 15243 17697 15252 17731
rect 15200 17688 15252 17697
rect 16764 17731 16816 17740
rect 16764 17697 16773 17731
rect 16773 17697 16807 17731
rect 16807 17697 16816 17731
rect 16764 17688 16816 17697
rect 21088 17824 21140 17876
rect 21180 17824 21232 17876
rect 21916 17867 21968 17876
rect 21916 17833 21925 17867
rect 21925 17833 21959 17867
rect 21959 17833 21968 17867
rect 21916 17824 21968 17833
rect 17960 17688 18012 17740
rect 4252 17484 4304 17536
rect 9864 17484 9916 17536
rect 10508 17484 10560 17536
rect 10692 17527 10744 17536
rect 10692 17493 10701 17527
rect 10701 17493 10735 17527
rect 10735 17493 10744 17527
rect 10692 17484 10744 17493
rect 11520 17552 11572 17604
rect 13820 17620 13872 17672
rect 14832 17620 14884 17672
rect 12992 17552 13044 17604
rect 15292 17595 15344 17604
rect 15292 17561 15301 17595
rect 15301 17561 15335 17595
rect 15335 17561 15344 17595
rect 15844 17595 15896 17604
rect 15292 17552 15344 17561
rect 15844 17561 15853 17595
rect 15853 17561 15887 17595
rect 15887 17561 15896 17595
rect 15844 17552 15896 17561
rect 15660 17484 15712 17536
rect 16488 17595 16540 17604
rect 16488 17561 16497 17595
rect 16497 17561 16531 17595
rect 16531 17561 16540 17595
rect 16488 17552 16540 17561
rect 21364 17756 21416 17808
rect 18420 17688 18472 17740
rect 22468 17688 22520 17740
rect 23296 17688 23348 17740
rect 30564 17756 30616 17808
rect 27804 17688 27856 17740
rect 18236 17620 18288 17672
rect 20168 17620 20220 17672
rect 21640 17620 21692 17672
rect 27620 17620 27672 17672
rect 18880 17484 18932 17536
rect 19984 17484 20036 17536
rect 20260 17484 20312 17536
rect 23848 17552 23900 17604
rect 25964 17595 26016 17604
rect 25964 17561 25973 17595
rect 25973 17561 26007 17595
rect 26007 17561 26016 17595
rect 25964 17552 26016 17561
rect 22192 17484 22244 17536
rect 24768 17484 24820 17536
rect 28172 17484 28224 17536
rect 31300 17484 31352 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 7932 17323 7984 17332
rect 7932 17289 7941 17323
rect 7941 17289 7975 17323
rect 7975 17289 7984 17323
rect 7932 17280 7984 17289
rect 4252 17255 4304 17264
rect 4252 17221 4261 17255
rect 4261 17221 4295 17255
rect 4295 17221 4304 17255
rect 4252 17212 4304 17221
rect 5172 17255 5224 17264
rect 5172 17221 5181 17255
rect 5181 17221 5215 17255
rect 5215 17221 5224 17255
rect 5172 17212 5224 17221
rect 6368 17212 6420 17264
rect 1768 17187 1820 17196
rect 1768 17153 1777 17187
rect 1777 17153 1811 17187
rect 1811 17153 1820 17187
rect 1768 17144 1820 17153
rect 7840 17187 7892 17196
rect 4804 17076 4856 17128
rect 1952 17008 2004 17060
rect 7840 17153 7849 17187
rect 7849 17153 7883 17187
rect 7883 17153 7892 17187
rect 7840 17144 7892 17153
rect 8300 17144 8352 17196
rect 11520 17280 11572 17332
rect 11612 17280 11664 17332
rect 16488 17280 16540 17332
rect 9588 17212 9640 17264
rect 10876 17212 10928 17264
rect 9772 17187 9824 17196
rect 9772 17153 9781 17187
rect 9781 17153 9815 17187
rect 9815 17153 9824 17187
rect 9772 17144 9824 17153
rect 9864 17144 9916 17196
rect 10232 17144 10284 17196
rect 11428 17144 11480 17196
rect 12256 17212 12308 17264
rect 20260 17280 20312 17332
rect 17132 17255 17184 17264
rect 17132 17221 17141 17255
rect 17141 17221 17175 17255
rect 17175 17221 17184 17255
rect 17132 17212 17184 17221
rect 18880 17255 18932 17264
rect 18880 17221 18889 17255
rect 18889 17221 18923 17255
rect 18923 17221 18932 17255
rect 18880 17212 18932 17221
rect 18972 17255 19024 17264
rect 18972 17221 18981 17255
rect 18981 17221 19015 17255
rect 19015 17221 19024 17255
rect 18972 17212 19024 17221
rect 19156 17212 19208 17264
rect 23296 17280 23348 17332
rect 23388 17280 23440 17332
rect 22192 17255 22244 17264
rect 10692 17076 10744 17128
rect 11060 17051 11112 17060
rect 1584 16983 1636 16992
rect 1584 16949 1593 16983
rect 1593 16949 1627 16983
rect 1627 16949 1636 16983
rect 1584 16940 1636 16949
rect 7656 16940 7708 16992
rect 8576 16983 8628 16992
rect 8576 16949 8585 16983
rect 8585 16949 8619 16983
rect 8619 16949 8628 16983
rect 8576 16940 8628 16949
rect 9864 16983 9916 16992
rect 9864 16949 9873 16983
rect 9873 16949 9907 16983
rect 9907 16949 9916 16983
rect 9864 16940 9916 16949
rect 10324 16940 10376 16992
rect 10692 16940 10744 16992
rect 11060 17017 11069 17051
rect 11069 17017 11103 17051
rect 11103 17017 11112 17051
rect 11060 17008 11112 17017
rect 11796 17076 11848 17128
rect 14280 17144 14332 17196
rect 13544 17076 13596 17128
rect 14924 17076 14976 17128
rect 15936 17144 15988 17196
rect 16120 17187 16172 17196
rect 16120 17153 16129 17187
rect 16129 17153 16163 17187
rect 16163 17153 16172 17187
rect 16120 17144 16172 17153
rect 16764 17144 16816 17196
rect 16672 17076 16724 17128
rect 17960 17076 18012 17128
rect 19616 17076 19668 17128
rect 20260 17144 20312 17196
rect 20812 17076 20864 17128
rect 14648 17008 14700 17060
rect 15108 17008 15160 17060
rect 18236 17008 18288 17060
rect 13452 16940 13504 16992
rect 14096 16940 14148 16992
rect 20076 16983 20128 16992
rect 20076 16949 20085 16983
rect 20085 16949 20119 16983
rect 20119 16949 20128 16983
rect 20076 16940 20128 16949
rect 20536 17008 20588 17060
rect 22192 17221 22201 17255
rect 22201 17221 22235 17255
rect 22235 17221 22244 17255
rect 22192 17212 22244 17221
rect 22284 17255 22336 17264
rect 22284 17221 22293 17255
rect 22293 17221 22327 17255
rect 22327 17221 22336 17255
rect 22284 17212 22336 17221
rect 22836 17212 22888 17264
rect 23204 17255 23256 17264
rect 23204 17221 23213 17255
rect 23213 17221 23247 17255
rect 23247 17221 23256 17255
rect 23204 17212 23256 17221
rect 24216 17255 24268 17264
rect 24216 17221 24225 17255
rect 24225 17221 24259 17255
rect 24259 17221 24268 17255
rect 24216 17212 24268 17221
rect 30196 17280 30248 17332
rect 37924 17212 37976 17264
rect 28172 17187 28224 17196
rect 28172 17153 28181 17187
rect 28181 17153 28215 17187
rect 28215 17153 28224 17187
rect 28172 17144 28224 17153
rect 28724 17144 28776 17196
rect 32588 17144 32640 17196
rect 24400 17119 24452 17128
rect 22560 17008 22612 17060
rect 24400 17085 24409 17119
rect 24409 17085 24443 17119
rect 24443 17085 24452 17119
rect 24400 17076 24452 17085
rect 29828 17076 29880 17128
rect 24952 17008 25004 17060
rect 38200 17051 38252 17060
rect 38200 17017 38209 17051
rect 38209 17017 38243 17051
rect 38243 17017 38252 17051
rect 38200 17008 38252 17017
rect 24584 16940 24636 16992
rect 24768 16940 24820 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 3700 16736 3752 16788
rect 9680 16736 9732 16788
rect 9864 16736 9916 16788
rect 14464 16736 14516 16788
rect 16028 16736 16080 16788
rect 16304 16736 16356 16788
rect 17132 16736 17184 16788
rect 18972 16736 19024 16788
rect 6828 16668 6880 16720
rect 1584 16600 1636 16652
rect 7012 16643 7064 16652
rect 7012 16609 7021 16643
rect 7021 16609 7055 16643
rect 7055 16609 7064 16643
rect 7012 16600 7064 16609
rect 8576 16668 8628 16720
rect 14740 16668 14792 16720
rect 14924 16711 14976 16720
rect 14924 16677 14933 16711
rect 14933 16677 14967 16711
rect 14967 16677 14976 16711
rect 14924 16668 14976 16677
rect 10876 16643 10928 16652
rect 10876 16609 10885 16643
rect 10885 16609 10919 16643
rect 10919 16609 10928 16643
rect 10876 16600 10928 16609
rect 11520 16600 11572 16652
rect 12072 16600 12124 16652
rect 15568 16600 15620 16652
rect 16488 16600 16540 16652
rect 24216 16736 24268 16788
rect 24400 16668 24452 16720
rect 9680 16532 9732 16584
rect 10048 16532 10100 16584
rect 11428 16575 11480 16584
rect 11428 16541 11437 16575
rect 11437 16541 11471 16575
rect 11471 16541 11480 16575
rect 11428 16532 11480 16541
rect 11612 16532 11664 16584
rect 15476 16575 15528 16584
rect 15476 16541 15485 16575
rect 15485 16541 15519 16575
rect 15519 16541 15528 16575
rect 15476 16532 15528 16541
rect 7104 16507 7156 16516
rect 7104 16473 7113 16507
rect 7113 16473 7147 16507
rect 7147 16473 7156 16507
rect 8024 16507 8076 16516
rect 7104 16464 7156 16473
rect 8024 16473 8033 16507
rect 8033 16473 8067 16507
rect 8067 16473 8076 16507
rect 8024 16464 8076 16473
rect 9220 16464 9272 16516
rect 10600 16464 10652 16516
rect 12624 16464 12676 16516
rect 12900 16464 12952 16516
rect 14096 16464 14148 16516
rect 8484 16396 8536 16448
rect 14464 16507 14516 16516
rect 14464 16473 14473 16507
rect 14473 16473 14507 16507
rect 14507 16473 14516 16507
rect 14464 16464 14516 16473
rect 15292 16464 15344 16516
rect 16672 16532 16724 16584
rect 16764 16532 16816 16584
rect 17684 16532 17736 16584
rect 20720 16532 20772 16584
rect 23112 16600 23164 16652
rect 22468 16575 22520 16584
rect 15936 16464 15988 16516
rect 19524 16507 19576 16516
rect 14556 16396 14608 16448
rect 19524 16473 19533 16507
rect 19533 16473 19567 16507
rect 19567 16473 19576 16507
rect 19524 16464 19576 16473
rect 19984 16464 20036 16516
rect 20260 16464 20312 16516
rect 22468 16541 22477 16575
rect 22477 16541 22511 16575
rect 22511 16541 22520 16575
rect 22468 16532 22520 16541
rect 22560 16575 22612 16584
rect 22560 16541 22569 16575
rect 22569 16541 22603 16575
rect 22603 16541 22612 16575
rect 23388 16575 23440 16584
rect 22560 16532 22612 16541
rect 23388 16541 23397 16575
rect 23397 16541 23431 16575
rect 23431 16541 23440 16575
rect 23388 16532 23440 16541
rect 22284 16464 22336 16516
rect 27436 16600 27488 16652
rect 29828 16643 29880 16652
rect 29828 16609 29837 16643
rect 29837 16609 29871 16643
rect 29871 16609 29880 16643
rect 29828 16600 29880 16609
rect 26332 16532 26384 16584
rect 28172 16464 28224 16516
rect 28540 16507 28592 16516
rect 28540 16473 28549 16507
rect 28549 16473 28583 16507
rect 28583 16473 28592 16507
rect 29920 16507 29972 16516
rect 28540 16464 28592 16473
rect 29920 16473 29929 16507
rect 29929 16473 29963 16507
rect 29963 16473 29972 16507
rect 29920 16464 29972 16473
rect 21088 16396 21140 16448
rect 24492 16396 24544 16448
rect 38016 16396 38068 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 7564 16192 7616 16244
rect 7380 16124 7432 16176
rect 8208 16124 8260 16176
rect 8484 16167 8536 16176
rect 8484 16133 8493 16167
rect 8493 16133 8527 16167
rect 8527 16133 8536 16167
rect 8484 16124 8536 16133
rect 9496 16124 9548 16176
rect 16120 16192 16172 16244
rect 9772 16167 9824 16176
rect 9772 16133 9781 16167
rect 9781 16133 9815 16167
rect 9815 16133 9824 16167
rect 9772 16124 9824 16133
rect 10784 16124 10836 16176
rect 13452 16167 13504 16176
rect 13452 16133 13461 16167
rect 13461 16133 13495 16167
rect 13495 16133 13504 16167
rect 13452 16124 13504 16133
rect 14372 16167 14424 16176
rect 14372 16133 14381 16167
rect 14381 16133 14415 16167
rect 14415 16133 14424 16167
rect 14372 16124 14424 16133
rect 15016 16124 15068 16176
rect 15660 16167 15712 16176
rect 15660 16133 15669 16167
rect 15669 16133 15703 16167
rect 15703 16133 15712 16167
rect 15660 16124 15712 16133
rect 16672 16124 16724 16176
rect 18512 16167 18564 16176
rect 2504 16099 2556 16108
rect 2504 16065 2513 16099
rect 2513 16065 2547 16099
rect 2547 16065 2556 16099
rect 2504 16056 2556 16065
rect 4068 16099 4120 16108
rect 4068 16065 4077 16099
rect 4077 16065 4111 16099
rect 4111 16065 4120 16099
rect 4068 16056 4120 16065
rect 1492 15988 1544 16040
rect 5632 16056 5684 16108
rect 6736 16056 6788 16108
rect 7288 16056 7340 16108
rect 9220 16056 9272 16108
rect 10968 16056 11020 16108
rect 14832 16099 14884 16108
rect 14832 16065 14841 16099
rect 14841 16065 14875 16099
rect 14875 16065 14884 16099
rect 14832 16056 14884 16065
rect 18512 16133 18521 16167
rect 18521 16133 18555 16167
rect 18555 16133 18564 16167
rect 18512 16124 18564 16133
rect 10600 15920 10652 15972
rect 12348 15988 12400 16040
rect 12808 16031 12860 16040
rect 12808 15997 12817 16031
rect 12817 15997 12851 16031
rect 12851 15997 12860 16031
rect 12808 15988 12860 15997
rect 13452 15988 13504 16040
rect 13728 15988 13780 16040
rect 15292 15988 15344 16040
rect 15568 16031 15620 16040
rect 15568 15997 15577 16031
rect 15577 15997 15611 16031
rect 15611 15997 15620 16031
rect 15568 15988 15620 15997
rect 17132 15988 17184 16040
rect 18420 16031 18472 16040
rect 18420 15997 18429 16031
rect 18429 15997 18463 16031
rect 18463 15997 18472 16031
rect 18420 15988 18472 15997
rect 18696 16031 18748 16040
rect 18696 15997 18705 16031
rect 18705 15997 18739 16031
rect 18739 15997 18748 16031
rect 18696 15988 18748 15997
rect 15200 15920 15252 15972
rect 15844 15920 15896 15972
rect 16120 15963 16172 15972
rect 16120 15929 16129 15963
rect 16129 15929 16163 15963
rect 16163 15929 16172 15963
rect 16120 15920 16172 15929
rect 1768 15895 1820 15904
rect 1768 15861 1777 15895
rect 1777 15861 1811 15895
rect 1811 15861 1820 15895
rect 1768 15852 1820 15861
rect 2596 15852 2648 15904
rect 6552 15852 6604 15904
rect 8576 15852 8628 15904
rect 9220 15852 9272 15904
rect 13544 15852 13596 15904
rect 17316 15920 17368 15972
rect 17592 15852 17644 15904
rect 17868 15852 17920 15904
rect 19984 16192 20036 16244
rect 28172 16235 28224 16244
rect 28172 16201 28181 16235
rect 28181 16201 28215 16235
rect 28215 16201 28224 16235
rect 28172 16192 28224 16201
rect 28264 16192 28316 16244
rect 30656 16192 30708 16244
rect 20076 16167 20128 16176
rect 20076 16133 20085 16167
rect 20085 16133 20119 16167
rect 20119 16133 20128 16167
rect 20076 16124 20128 16133
rect 20352 16124 20404 16176
rect 20720 16124 20772 16176
rect 21088 16099 21140 16108
rect 21088 16065 21097 16099
rect 21097 16065 21131 16099
rect 21131 16065 21140 16099
rect 21088 16056 21140 16065
rect 21916 16056 21968 16108
rect 23664 16056 23716 16108
rect 33600 16124 33652 16176
rect 22100 15988 22152 16040
rect 22928 15988 22980 16040
rect 23112 16031 23164 16040
rect 23112 15997 23121 16031
rect 23121 15997 23155 16031
rect 23155 15997 23164 16031
rect 23112 15988 23164 15997
rect 20076 15920 20128 15972
rect 20536 15963 20588 15972
rect 20536 15929 20545 15963
rect 20545 15929 20579 15963
rect 20579 15929 20588 15963
rect 20536 15920 20588 15929
rect 23204 15920 23256 15972
rect 27160 15988 27212 16040
rect 28540 15988 28592 16040
rect 27436 15920 27488 15972
rect 28356 15920 28408 15972
rect 38016 16099 38068 16108
rect 29276 16031 29328 16040
rect 29276 15997 29285 16031
rect 29285 15997 29319 16031
rect 29319 15997 29328 16031
rect 29276 15988 29328 15997
rect 38016 16065 38025 16099
rect 38025 16065 38059 16099
rect 38059 16065 38068 16099
rect 38016 16056 38068 16065
rect 30196 15920 30248 15972
rect 34796 15920 34848 15972
rect 22100 15895 22152 15904
rect 22100 15861 22109 15895
rect 22109 15861 22143 15895
rect 22143 15861 22152 15895
rect 22100 15852 22152 15861
rect 24216 15852 24268 15904
rect 28264 15852 28316 15904
rect 29920 15852 29972 15904
rect 30748 15895 30800 15904
rect 30748 15861 30757 15895
rect 30757 15861 30791 15895
rect 30791 15861 30800 15895
rect 30748 15852 30800 15861
rect 38200 15895 38252 15904
rect 38200 15861 38209 15895
rect 38209 15861 38243 15895
rect 38243 15861 38252 15895
rect 38200 15852 38252 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 2504 15648 2556 15700
rect 6460 15648 6512 15700
rect 12532 15648 12584 15700
rect 12624 15648 12676 15700
rect 15292 15648 15344 15700
rect 15844 15648 15896 15700
rect 16120 15648 16172 15700
rect 5264 15580 5316 15632
rect 8484 15580 8536 15632
rect 9588 15580 9640 15632
rect 12348 15580 12400 15632
rect 8024 15512 8076 15564
rect 1676 15444 1728 15496
rect 4896 15444 4948 15496
rect 5080 15444 5132 15496
rect 5816 15487 5868 15496
rect 5816 15453 5825 15487
rect 5825 15453 5859 15487
rect 5859 15453 5868 15487
rect 5816 15444 5868 15453
rect 6460 15487 6512 15496
rect 6460 15453 6469 15487
rect 6469 15453 6503 15487
rect 6503 15453 6512 15487
rect 6460 15444 6512 15453
rect 7380 15444 7432 15496
rect 8852 15512 8904 15564
rect 9220 15555 9272 15564
rect 9220 15521 9229 15555
rect 9229 15521 9263 15555
rect 9263 15521 9272 15555
rect 9220 15512 9272 15521
rect 9772 15555 9824 15564
rect 9772 15521 9781 15555
rect 9781 15521 9815 15555
rect 9815 15521 9824 15555
rect 9772 15512 9824 15521
rect 9864 15512 9916 15564
rect 8484 15444 8536 15496
rect 13820 15512 13872 15564
rect 13912 15512 13964 15564
rect 23112 15648 23164 15700
rect 24400 15648 24452 15700
rect 18236 15580 18288 15632
rect 18420 15580 18472 15632
rect 20628 15580 20680 15632
rect 24216 15580 24268 15632
rect 19984 15512 20036 15564
rect 20444 15555 20496 15564
rect 20444 15521 20453 15555
rect 20453 15521 20487 15555
rect 20487 15521 20496 15555
rect 20444 15512 20496 15521
rect 20720 15512 20772 15564
rect 22100 15512 22152 15564
rect 3608 15376 3660 15428
rect 7564 15376 7616 15428
rect 2412 15351 2464 15360
rect 2412 15317 2421 15351
rect 2421 15317 2455 15351
rect 2455 15317 2464 15351
rect 2412 15308 2464 15317
rect 5172 15308 5224 15360
rect 5356 15308 5408 15360
rect 6828 15308 6880 15360
rect 7196 15308 7248 15360
rect 9772 15376 9824 15428
rect 10876 15419 10928 15428
rect 10876 15385 10885 15419
rect 10885 15385 10919 15419
rect 10919 15385 10928 15419
rect 10876 15376 10928 15385
rect 10968 15419 11020 15428
rect 10968 15385 10977 15419
rect 10977 15385 11011 15419
rect 11011 15385 11020 15419
rect 10968 15376 11020 15385
rect 11888 15308 11940 15360
rect 18696 15487 18748 15496
rect 14372 15376 14424 15428
rect 14648 15419 14700 15428
rect 14648 15385 14657 15419
rect 14657 15385 14691 15419
rect 14691 15385 14700 15419
rect 14648 15376 14700 15385
rect 15568 15376 15620 15428
rect 17132 15376 17184 15428
rect 18696 15453 18705 15487
rect 18705 15453 18739 15487
rect 18739 15453 18748 15487
rect 18696 15444 18748 15453
rect 19340 15444 19392 15496
rect 22008 15444 22060 15496
rect 22376 15444 22428 15496
rect 26148 15580 26200 15632
rect 28172 15648 28224 15700
rect 28540 15691 28592 15700
rect 28540 15657 28549 15691
rect 28549 15657 28583 15691
rect 28583 15657 28592 15691
rect 28540 15648 28592 15657
rect 30196 15580 30248 15632
rect 26424 15512 26476 15564
rect 30748 15512 30800 15564
rect 26056 15444 26108 15496
rect 26516 15487 26568 15496
rect 26516 15453 26525 15487
rect 26525 15453 26559 15487
rect 26559 15453 26568 15487
rect 26516 15444 26568 15453
rect 27436 15444 27488 15496
rect 28356 15444 28408 15496
rect 29920 15487 29972 15496
rect 29920 15453 29929 15487
rect 29929 15453 29963 15487
rect 29963 15453 29972 15487
rect 29920 15444 29972 15453
rect 13084 15308 13136 15360
rect 13452 15308 13504 15360
rect 15016 15308 15068 15360
rect 17960 15376 18012 15428
rect 20076 15376 20128 15428
rect 19524 15308 19576 15360
rect 23664 15376 23716 15428
rect 24400 15376 24452 15428
rect 38108 15419 38160 15428
rect 38108 15385 38117 15419
rect 38117 15385 38151 15419
rect 38151 15385 38160 15419
rect 38108 15376 38160 15385
rect 21180 15308 21232 15360
rect 23296 15308 23348 15360
rect 24676 15308 24728 15360
rect 24768 15308 24820 15360
rect 26240 15308 26292 15360
rect 29000 15308 29052 15360
rect 38200 15351 38252 15360
rect 38200 15317 38209 15351
rect 38209 15317 38243 15351
rect 38243 15317 38252 15351
rect 38200 15308 38252 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 1676 14968 1728 15020
rect 2412 15011 2464 15020
rect 2412 14977 2421 15011
rect 2421 14977 2455 15011
rect 2455 14977 2464 15011
rect 2412 14968 2464 14977
rect 2596 15011 2648 15020
rect 2596 14977 2605 15011
rect 2605 14977 2639 15011
rect 2639 14977 2648 15011
rect 2596 14968 2648 14977
rect 5080 15036 5132 15088
rect 10600 15079 10652 15088
rect 10600 15045 10609 15079
rect 10609 15045 10643 15079
rect 10643 15045 10652 15079
rect 10600 15036 10652 15045
rect 4988 14968 5040 15020
rect 5816 15011 5868 15020
rect 5816 14977 5825 15011
rect 5825 14977 5859 15011
rect 5859 14977 5868 15011
rect 5816 14968 5868 14977
rect 6000 14968 6052 15020
rect 7472 14968 7524 15020
rect 8024 15011 8076 15020
rect 8024 14977 8033 15011
rect 8033 14977 8067 15011
rect 8067 14977 8076 15011
rect 8024 14968 8076 14977
rect 12532 15036 12584 15088
rect 13084 15036 13136 15088
rect 14556 15036 14608 15088
rect 11612 14968 11664 15020
rect 14924 15011 14976 15020
rect 7564 14900 7616 14952
rect 8392 14900 8444 14952
rect 9128 14943 9180 14952
rect 9128 14909 9137 14943
rect 9137 14909 9171 14943
rect 9171 14909 9180 14943
rect 9128 14900 9180 14909
rect 9680 14900 9732 14952
rect 10232 14900 10284 14952
rect 11336 14900 11388 14952
rect 11704 14900 11756 14952
rect 14924 14977 14933 15011
rect 14933 14977 14967 15011
rect 14967 14977 14976 15011
rect 14924 14968 14976 14977
rect 15384 14968 15436 15020
rect 12624 14900 12676 14952
rect 14372 14943 14424 14952
rect 14372 14909 14381 14943
rect 14381 14909 14415 14943
rect 14415 14909 14424 14943
rect 14372 14900 14424 14909
rect 15200 14943 15252 14952
rect 15200 14909 15209 14943
rect 15209 14909 15243 14943
rect 15243 14909 15252 14943
rect 15200 14900 15252 14909
rect 17776 15104 17828 15156
rect 19524 15104 19576 15156
rect 20076 15104 20128 15156
rect 22836 15104 22888 15156
rect 23204 15104 23256 15156
rect 26056 15147 26108 15156
rect 17592 15079 17644 15088
rect 17592 15045 17601 15079
rect 17601 15045 17635 15079
rect 17635 15045 17644 15079
rect 17592 15036 17644 15045
rect 20536 15036 20588 15088
rect 18972 15011 19024 15020
rect 18972 14977 18981 15011
rect 18981 14977 19015 15011
rect 19015 14977 19024 15011
rect 18972 14968 19024 14977
rect 5632 14832 5684 14884
rect 10784 14832 10836 14884
rect 10968 14832 11020 14884
rect 16304 14900 16356 14952
rect 18144 14943 18196 14952
rect 18144 14909 18153 14943
rect 18153 14909 18187 14943
rect 18187 14909 18196 14943
rect 18144 14900 18196 14909
rect 19984 14900 20036 14952
rect 20076 14943 20128 14952
rect 20076 14909 20085 14943
rect 20085 14909 20119 14943
rect 20119 14909 20128 14943
rect 20076 14900 20128 14909
rect 20536 14900 20588 14952
rect 24676 15079 24728 15088
rect 24676 15045 24685 15079
rect 24685 15045 24719 15079
rect 24719 15045 24728 15079
rect 24676 15036 24728 15045
rect 26056 15113 26065 15147
rect 26065 15113 26099 15147
rect 26099 15113 26108 15147
rect 26056 15104 26108 15113
rect 26240 15011 26292 15020
rect 26240 14977 26249 15011
rect 26249 14977 26283 15011
rect 26283 14977 26292 15011
rect 26240 14968 26292 14977
rect 29000 14968 29052 15020
rect 29092 14968 29144 15020
rect 30472 14968 30524 15020
rect 31300 14968 31352 15020
rect 21456 14900 21508 14952
rect 21916 14900 21968 14952
rect 23112 14943 23164 14952
rect 23112 14909 23121 14943
rect 23121 14909 23155 14943
rect 23155 14909 23164 14943
rect 23112 14900 23164 14909
rect 24768 14900 24820 14952
rect 27344 14943 27396 14952
rect 27344 14909 27353 14943
rect 27353 14909 27387 14943
rect 27387 14909 27396 14943
rect 27344 14900 27396 14909
rect 29276 14900 29328 14952
rect 2688 14764 2740 14816
rect 3056 14807 3108 14816
rect 3056 14773 3065 14807
rect 3065 14773 3099 14807
rect 3099 14773 3108 14807
rect 3056 14764 3108 14773
rect 3792 14764 3844 14816
rect 5908 14807 5960 14816
rect 5908 14773 5917 14807
rect 5917 14773 5951 14807
rect 5951 14773 5960 14807
rect 5908 14764 5960 14773
rect 15016 14764 15068 14816
rect 15108 14764 15160 14816
rect 25228 14832 25280 14884
rect 16672 14764 16724 14816
rect 17960 14764 18012 14816
rect 19432 14764 19484 14816
rect 20444 14764 20496 14816
rect 21088 14764 21140 14816
rect 22744 14764 22796 14816
rect 23112 14764 23164 14816
rect 26884 14764 26936 14816
rect 28816 14807 28868 14816
rect 28816 14773 28825 14807
rect 28825 14773 28859 14807
rect 28859 14773 28868 14807
rect 28816 14764 28868 14773
rect 29920 14764 29972 14816
rect 31484 14764 31536 14816
rect 34428 14764 34480 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 1860 14560 1912 14612
rect 3056 14603 3108 14612
rect 3056 14569 3065 14603
rect 3065 14569 3099 14603
rect 3099 14569 3108 14603
rect 3056 14560 3108 14569
rect 10600 14560 10652 14612
rect 2688 14467 2740 14476
rect 2688 14433 2697 14467
rect 2697 14433 2731 14467
rect 2731 14433 2740 14467
rect 2688 14424 2740 14433
rect 1768 14399 1820 14408
rect 1768 14365 1777 14399
rect 1777 14365 1811 14399
rect 1811 14365 1820 14399
rect 1768 14356 1820 14365
rect 2504 14399 2556 14408
rect 2504 14365 2513 14399
rect 2513 14365 2547 14399
rect 2547 14365 2556 14399
rect 2504 14356 2556 14365
rect 4712 14356 4764 14408
rect 4896 14399 4948 14408
rect 4896 14365 4905 14399
rect 4905 14365 4939 14399
rect 4939 14365 4948 14399
rect 4896 14356 4948 14365
rect 5632 14356 5684 14408
rect 8392 14492 8444 14544
rect 8484 14492 8536 14544
rect 9588 14492 9640 14544
rect 15752 14560 15804 14612
rect 16856 14560 16908 14612
rect 17040 14560 17092 14612
rect 19432 14560 19484 14612
rect 20536 14603 20588 14612
rect 20536 14569 20545 14603
rect 20545 14569 20579 14603
rect 20579 14569 20588 14603
rect 20536 14560 20588 14569
rect 7840 14467 7892 14476
rect 7840 14433 7849 14467
rect 7849 14433 7883 14467
rect 7883 14433 7892 14467
rect 7840 14424 7892 14433
rect 6276 14356 6328 14408
rect 6460 14356 6512 14408
rect 7380 14356 7432 14408
rect 7104 14288 7156 14340
rect 7564 14331 7616 14340
rect 7564 14297 7573 14331
rect 7573 14297 7607 14331
rect 7607 14297 7616 14331
rect 7564 14288 7616 14297
rect 7656 14331 7708 14340
rect 7656 14297 7665 14331
rect 7665 14297 7699 14331
rect 7699 14297 7708 14331
rect 7656 14288 7708 14297
rect 4712 14220 4764 14272
rect 5632 14263 5684 14272
rect 5632 14229 5641 14263
rect 5641 14229 5675 14263
rect 5675 14229 5684 14263
rect 5632 14220 5684 14229
rect 6920 14220 6972 14272
rect 12348 14424 12400 14476
rect 14280 14492 14332 14544
rect 14464 14492 14516 14544
rect 22008 14560 22060 14612
rect 23204 14535 23256 14544
rect 23204 14501 23213 14535
rect 23213 14501 23247 14535
rect 23247 14501 23256 14535
rect 23204 14492 23256 14501
rect 16120 14424 16172 14476
rect 18236 14424 18288 14476
rect 21824 14424 21876 14476
rect 25412 14424 25464 14476
rect 10232 14356 10284 14408
rect 11060 14399 11112 14408
rect 11060 14365 11069 14399
rect 11069 14365 11103 14399
rect 11103 14365 11112 14399
rect 11060 14356 11112 14365
rect 12624 14356 12676 14408
rect 14924 14356 14976 14408
rect 15292 14399 15344 14408
rect 15292 14365 15301 14399
rect 15301 14365 15335 14399
rect 15335 14365 15344 14399
rect 15292 14356 15344 14365
rect 16948 14356 17000 14408
rect 18972 14356 19024 14408
rect 20444 14399 20496 14408
rect 20444 14365 20453 14399
rect 20453 14365 20487 14399
rect 20487 14365 20496 14399
rect 20444 14356 20496 14365
rect 23572 14356 23624 14408
rect 24308 14356 24360 14408
rect 25688 14467 25740 14476
rect 25688 14433 25697 14467
rect 25697 14433 25731 14467
rect 25731 14433 25740 14467
rect 25688 14424 25740 14433
rect 38200 14424 38252 14476
rect 9220 14288 9272 14340
rect 11336 14331 11388 14340
rect 11336 14297 11345 14331
rect 11345 14297 11379 14331
rect 11379 14297 11388 14331
rect 11336 14288 11388 14297
rect 8760 14220 8812 14272
rect 14372 14288 14424 14340
rect 13084 14220 13136 14272
rect 17040 14331 17092 14340
rect 17040 14297 17049 14331
rect 17049 14297 17083 14331
rect 17083 14297 17092 14331
rect 17040 14288 17092 14297
rect 17776 14288 17828 14340
rect 21272 14288 21324 14340
rect 21548 14331 21600 14340
rect 21548 14297 21557 14331
rect 21557 14297 21591 14331
rect 21591 14297 21600 14331
rect 22652 14331 22704 14340
rect 21548 14288 21600 14297
rect 22652 14297 22661 14331
rect 22661 14297 22695 14331
rect 22695 14297 22704 14331
rect 22652 14288 22704 14297
rect 17316 14220 17368 14272
rect 17592 14220 17644 14272
rect 18328 14220 18380 14272
rect 19156 14220 19208 14272
rect 19984 14220 20036 14272
rect 25780 14331 25832 14340
rect 25780 14297 25789 14331
rect 25789 14297 25823 14331
rect 25823 14297 25832 14331
rect 25780 14288 25832 14297
rect 24308 14220 24360 14272
rect 24676 14263 24728 14272
rect 24676 14229 24685 14263
rect 24685 14229 24719 14263
rect 24719 14229 24728 14263
rect 24676 14220 24728 14229
rect 24768 14220 24820 14272
rect 27252 14331 27304 14340
rect 27252 14297 27261 14331
rect 27261 14297 27295 14331
rect 27295 14297 27304 14331
rect 27252 14288 27304 14297
rect 28264 14331 28316 14340
rect 26332 14220 26384 14272
rect 28264 14297 28273 14331
rect 28273 14297 28307 14331
rect 28307 14297 28316 14331
rect 28264 14288 28316 14297
rect 28816 14356 28868 14408
rect 32588 14288 32640 14340
rect 38016 14220 38068 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 3516 14016 3568 14068
rect 4068 14016 4120 14068
rect 3056 13948 3108 14000
rect 1584 13923 1636 13932
rect 1584 13889 1593 13923
rect 1593 13889 1627 13923
rect 1627 13889 1636 13923
rect 1584 13880 1636 13889
rect 5540 14016 5592 14068
rect 6920 14059 6972 14068
rect 6920 14025 6929 14059
rect 6929 14025 6963 14059
rect 6963 14025 6972 14059
rect 6920 14016 6972 14025
rect 7472 14016 7524 14068
rect 7380 13948 7432 14000
rect 7748 13991 7800 14000
rect 7748 13957 7757 13991
rect 7757 13957 7791 13991
rect 7791 13957 7800 13991
rect 7748 13948 7800 13957
rect 8300 13948 8352 14000
rect 4620 13880 4672 13932
rect 5448 13812 5500 13864
rect 1768 13719 1820 13728
rect 1768 13685 1777 13719
rect 1777 13685 1811 13719
rect 1811 13685 1820 13719
rect 1768 13676 1820 13685
rect 6092 13880 6144 13932
rect 6920 13880 6972 13932
rect 7380 13812 7432 13864
rect 7840 13812 7892 13864
rect 9772 13948 9824 14000
rect 10232 13923 10284 13932
rect 10232 13889 10241 13923
rect 10241 13889 10275 13923
rect 10275 13889 10284 13923
rect 13084 13948 13136 14000
rect 13820 13948 13872 14000
rect 19984 14016 20036 14068
rect 20076 14016 20128 14068
rect 20352 14016 20404 14068
rect 21548 14016 21600 14068
rect 21916 14016 21968 14068
rect 15384 13948 15436 14000
rect 11888 13923 11940 13932
rect 10232 13880 10284 13889
rect 11888 13889 11897 13923
rect 11897 13889 11931 13923
rect 11931 13889 11940 13923
rect 11888 13880 11940 13889
rect 10508 13812 10560 13864
rect 11060 13855 11112 13864
rect 11060 13821 11069 13855
rect 11069 13821 11103 13855
rect 11103 13821 11112 13855
rect 11060 13812 11112 13821
rect 14004 13812 14056 13864
rect 16120 13812 16172 13864
rect 17776 13812 17828 13864
rect 19340 13948 19392 14000
rect 21824 13948 21876 14000
rect 25780 14016 25832 14068
rect 26332 14059 26384 14068
rect 26332 14025 26341 14059
rect 26341 14025 26375 14059
rect 26375 14025 26384 14059
rect 26332 14016 26384 14025
rect 27252 14016 27304 14068
rect 28264 14016 28316 14068
rect 36176 14016 36228 14068
rect 24032 13991 24084 14000
rect 24032 13957 24041 13991
rect 24041 13957 24075 13991
rect 24075 13957 24084 13991
rect 24032 13948 24084 13957
rect 24584 13948 24636 14000
rect 24768 13948 24820 14000
rect 9220 13744 9272 13796
rect 9772 13744 9824 13796
rect 11244 13744 11296 13796
rect 6184 13676 6236 13728
rect 6736 13676 6788 13728
rect 6920 13676 6972 13728
rect 7196 13676 7248 13728
rect 7748 13676 7800 13728
rect 8208 13676 8260 13728
rect 8484 13676 8536 13728
rect 12348 13676 12400 13728
rect 16580 13744 16632 13796
rect 18420 13744 18472 13796
rect 20536 13812 20588 13864
rect 22100 13880 22152 13932
rect 25596 13923 25648 13932
rect 25596 13889 25605 13923
rect 25605 13889 25639 13923
rect 25639 13889 25648 13923
rect 25596 13880 25648 13889
rect 25872 13880 25924 13932
rect 27160 13923 27212 13932
rect 27160 13889 27169 13923
rect 27169 13889 27203 13923
rect 27203 13889 27212 13923
rect 27160 13880 27212 13889
rect 27344 13880 27396 13932
rect 31484 13923 31536 13932
rect 31484 13889 31493 13923
rect 31493 13889 31527 13923
rect 31527 13889 31536 13923
rect 31484 13880 31536 13889
rect 38016 13923 38068 13932
rect 38016 13889 38025 13923
rect 38025 13889 38059 13923
rect 38059 13889 38068 13923
rect 38016 13880 38068 13889
rect 14096 13676 14148 13728
rect 14464 13676 14516 13728
rect 17224 13676 17276 13728
rect 20996 13744 21048 13796
rect 21916 13744 21968 13796
rect 22928 13744 22980 13796
rect 23388 13812 23440 13864
rect 29736 13812 29788 13864
rect 25964 13744 26016 13796
rect 20352 13676 20404 13728
rect 21456 13676 21508 13728
rect 27620 13676 27672 13728
rect 28448 13676 28500 13728
rect 31300 13719 31352 13728
rect 31300 13685 31309 13719
rect 31309 13685 31343 13719
rect 31343 13685 31352 13719
rect 31300 13676 31352 13685
rect 38200 13719 38252 13728
rect 38200 13685 38209 13719
rect 38209 13685 38243 13719
rect 38243 13685 38252 13719
rect 38200 13676 38252 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 5908 13472 5960 13524
rect 8300 13472 8352 13524
rect 9128 13472 9180 13524
rect 4620 13336 4672 13388
rect 5264 13336 5316 13388
rect 6736 13336 6788 13388
rect 7840 13336 7892 13388
rect 8300 13336 8352 13388
rect 9128 13379 9180 13388
rect 9128 13345 9137 13379
rect 9137 13345 9171 13379
rect 9171 13345 9180 13379
rect 9128 13336 9180 13345
rect 9772 13336 9824 13388
rect 4712 13311 4764 13320
rect 4712 13277 4721 13311
rect 4721 13277 4755 13311
rect 4755 13277 4764 13311
rect 4712 13268 4764 13277
rect 5816 13311 5868 13320
rect 5816 13277 5825 13311
rect 5825 13277 5859 13311
rect 5859 13277 5868 13311
rect 5816 13268 5868 13277
rect 4620 13132 4672 13184
rect 4712 13132 4764 13184
rect 4896 13132 4948 13184
rect 7012 13200 7064 13252
rect 7196 13200 7248 13252
rect 7472 13132 7524 13184
rect 8484 13132 8536 13184
rect 9312 13200 9364 13252
rect 12532 13472 12584 13524
rect 15200 13472 15252 13524
rect 17040 13472 17092 13524
rect 17500 13472 17552 13524
rect 18236 13472 18288 13524
rect 19708 13472 19760 13524
rect 21824 13515 21876 13524
rect 21824 13481 21833 13515
rect 21833 13481 21867 13515
rect 21867 13481 21876 13515
rect 21824 13472 21876 13481
rect 13636 13447 13688 13456
rect 13636 13413 13645 13447
rect 13645 13413 13679 13447
rect 13679 13413 13688 13447
rect 13636 13404 13688 13413
rect 12164 13379 12216 13388
rect 12164 13345 12173 13379
rect 12173 13345 12207 13379
rect 12207 13345 12216 13379
rect 12164 13336 12216 13345
rect 12716 13336 12768 13388
rect 13728 13336 13780 13388
rect 14556 13379 14608 13388
rect 14556 13345 14565 13379
rect 14565 13345 14599 13379
rect 14599 13345 14608 13379
rect 14556 13336 14608 13345
rect 14924 13336 14976 13388
rect 11888 13311 11940 13320
rect 11888 13277 11897 13311
rect 11897 13277 11931 13311
rect 11931 13277 11940 13311
rect 11888 13268 11940 13277
rect 14004 13268 14056 13320
rect 15016 13200 15068 13252
rect 14096 13132 14148 13184
rect 21088 13336 21140 13388
rect 16580 13311 16632 13320
rect 16580 13277 16589 13311
rect 16589 13277 16623 13311
rect 16623 13277 16632 13311
rect 16580 13268 16632 13277
rect 19340 13268 19392 13320
rect 21640 13268 21692 13320
rect 16856 13243 16908 13252
rect 16856 13209 16865 13243
rect 16865 13209 16899 13243
rect 16899 13209 16908 13243
rect 16856 13200 16908 13209
rect 17316 13200 17368 13252
rect 19708 13243 19760 13252
rect 19708 13209 19717 13243
rect 19717 13209 19751 13243
rect 19751 13209 19760 13243
rect 19708 13200 19760 13209
rect 21824 13200 21876 13252
rect 16304 13132 16356 13184
rect 26700 13472 26752 13524
rect 27620 13472 27672 13524
rect 29736 13515 29788 13524
rect 29736 13481 29745 13515
rect 29745 13481 29779 13515
rect 29779 13481 29788 13515
rect 29736 13472 29788 13481
rect 22836 13404 22888 13456
rect 23296 13336 23348 13388
rect 24400 13404 24452 13456
rect 24676 13379 24728 13388
rect 24676 13345 24685 13379
rect 24685 13345 24719 13379
rect 24719 13345 24728 13379
rect 24676 13336 24728 13345
rect 27436 13404 27488 13456
rect 30840 13336 30892 13388
rect 22928 13268 22980 13320
rect 27620 13268 27672 13320
rect 24492 13200 24544 13252
rect 29184 13268 29236 13320
rect 29920 13311 29972 13320
rect 29920 13277 29929 13311
rect 29929 13277 29963 13311
rect 29963 13277 29972 13311
rect 29920 13268 29972 13277
rect 23940 13132 23992 13184
rect 29092 13200 29144 13252
rect 29368 13132 29420 13184
rect 30656 13132 30708 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 3976 12928 4028 12980
rect 8760 12928 8812 12980
rect 9036 12928 9088 12980
rect 9312 12928 9364 12980
rect 3240 12860 3292 12912
rect 7380 12860 7432 12912
rect 11612 12928 11664 12980
rect 11980 12928 12032 12980
rect 14004 12928 14056 12980
rect 14740 12928 14792 12980
rect 15016 12928 15068 12980
rect 15384 12928 15436 12980
rect 16212 12971 16264 12980
rect 1860 12792 1912 12844
rect 5080 12792 5132 12844
rect 5908 12792 5960 12844
rect 6184 12792 6236 12844
rect 6828 12792 6880 12844
rect 7196 12792 7248 12844
rect 7748 12835 7800 12844
rect 7472 12724 7524 12776
rect 7748 12801 7757 12835
rect 7757 12801 7791 12835
rect 7791 12801 7800 12835
rect 7748 12792 7800 12801
rect 7656 12724 7708 12776
rect 9772 12724 9824 12776
rect 10324 12767 10376 12776
rect 10324 12733 10333 12767
rect 10333 12733 10367 12767
rect 10367 12733 10376 12767
rect 10324 12724 10376 12733
rect 6920 12656 6972 12708
rect 1768 12631 1820 12640
rect 1768 12597 1777 12631
rect 1777 12597 1811 12631
rect 1811 12597 1820 12631
rect 1768 12588 1820 12597
rect 3608 12588 3660 12640
rect 3976 12588 4028 12640
rect 4712 12588 4764 12640
rect 7380 12656 7432 12708
rect 9036 12656 9088 12708
rect 9220 12656 9272 12708
rect 13820 12860 13872 12912
rect 16212 12937 16221 12971
rect 16221 12937 16255 12971
rect 16255 12937 16264 12971
rect 16212 12928 16264 12937
rect 19524 12928 19576 12980
rect 19984 12928 20036 12980
rect 17224 12860 17276 12912
rect 22652 12928 22704 12980
rect 23848 12860 23900 12912
rect 11980 12792 12032 12844
rect 14004 12792 14056 12844
rect 19340 12792 19392 12844
rect 22008 12792 22060 12844
rect 22468 12792 22520 12844
rect 26240 12928 26292 12980
rect 26424 12928 26476 12980
rect 26700 12928 26752 12980
rect 29184 12971 29236 12980
rect 29184 12937 29193 12971
rect 29193 12937 29227 12971
rect 29227 12937 29236 12971
rect 29184 12928 29236 12937
rect 24308 12903 24360 12912
rect 24308 12869 24317 12903
rect 24317 12869 24351 12903
rect 24351 12869 24360 12903
rect 24308 12860 24360 12869
rect 25688 12835 25740 12844
rect 25688 12801 25697 12835
rect 25697 12801 25731 12835
rect 25731 12801 25740 12835
rect 25688 12792 25740 12801
rect 11704 12724 11756 12776
rect 14096 12724 14148 12776
rect 15384 12724 15436 12776
rect 15752 12724 15804 12776
rect 16304 12724 16356 12776
rect 16580 12724 16632 12776
rect 20352 12724 20404 12776
rect 20720 12724 20772 12776
rect 23940 12724 23992 12776
rect 24676 12724 24728 12776
rect 26424 12724 26476 12776
rect 8208 12588 8260 12640
rect 8576 12588 8628 12640
rect 11428 12656 11480 12708
rect 9680 12588 9732 12640
rect 14188 12588 14240 12640
rect 14464 12588 14516 12640
rect 17500 12588 17552 12640
rect 21272 12656 21324 12708
rect 21732 12656 21784 12708
rect 21640 12588 21692 12640
rect 22376 12656 22428 12708
rect 22836 12656 22888 12708
rect 30472 12792 30524 12844
rect 30656 12835 30708 12844
rect 30656 12801 30665 12835
rect 30665 12801 30699 12835
rect 30699 12801 30708 12835
rect 30656 12792 30708 12801
rect 31300 12792 31352 12844
rect 34428 12792 34480 12844
rect 27988 12767 28040 12776
rect 27988 12733 27997 12767
rect 27997 12733 28031 12767
rect 28031 12733 28040 12767
rect 27988 12724 28040 12733
rect 28172 12767 28224 12776
rect 28172 12733 28181 12767
rect 28181 12733 28215 12767
rect 28215 12733 28224 12767
rect 28172 12724 28224 12733
rect 29368 12656 29420 12708
rect 29000 12588 29052 12640
rect 38200 12631 38252 12640
rect 38200 12597 38209 12631
rect 38209 12597 38243 12631
rect 38243 12597 38252 12631
rect 38200 12588 38252 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 5448 12384 5500 12436
rect 9220 12384 9272 12436
rect 9864 12427 9916 12436
rect 9864 12393 9873 12427
rect 9873 12393 9907 12427
rect 9907 12393 9916 12427
rect 9864 12384 9916 12393
rect 10048 12384 10100 12436
rect 11428 12384 11480 12436
rect 13268 12384 13320 12436
rect 13820 12384 13872 12436
rect 15752 12384 15804 12436
rect 18512 12427 18564 12436
rect 2964 12316 3016 12368
rect 5908 12316 5960 12368
rect 6736 12291 6788 12300
rect 6736 12257 6745 12291
rect 6745 12257 6779 12291
rect 6779 12257 6788 12291
rect 6736 12248 6788 12257
rect 9680 12248 9732 12300
rect 9128 12223 9180 12232
rect 9128 12189 9137 12223
rect 9137 12189 9171 12223
rect 9171 12189 9180 12223
rect 9128 12180 9180 12189
rect 10416 12316 10468 12368
rect 11244 12248 11296 12300
rect 10416 12223 10468 12232
rect 10416 12189 10425 12223
rect 10425 12189 10459 12223
rect 10459 12189 10468 12223
rect 10416 12180 10468 12189
rect 7104 12112 7156 12164
rect 2596 12044 2648 12096
rect 8484 12087 8536 12096
rect 8484 12053 8493 12087
rect 8493 12053 8527 12087
rect 8527 12053 8536 12087
rect 8484 12044 8536 12053
rect 10784 12044 10836 12096
rect 10968 12112 11020 12164
rect 12256 12248 12308 12300
rect 12716 12248 12768 12300
rect 15568 12248 15620 12300
rect 16580 12248 16632 12300
rect 18512 12393 18521 12427
rect 18521 12393 18555 12427
rect 18555 12393 18564 12427
rect 18512 12384 18564 12393
rect 18236 12316 18288 12368
rect 20904 12384 20956 12436
rect 21732 12384 21784 12436
rect 22100 12384 22152 12436
rect 23204 12384 23256 12436
rect 21456 12316 21508 12368
rect 24584 12384 24636 12436
rect 26424 12427 26476 12436
rect 26424 12393 26433 12427
rect 26433 12393 26467 12427
rect 26467 12393 26476 12427
rect 26424 12384 26476 12393
rect 28172 12384 28224 12436
rect 33784 12384 33836 12436
rect 34520 12384 34572 12436
rect 19432 12248 19484 12300
rect 21548 12248 21600 12300
rect 21916 12248 21968 12300
rect 22100 12248 22152 12300
rect 23388 12248 23440 12300
rect 12808 12180 12860 12232
rect 13728 12180 13780 12232
rect 15476 12180 15528 12232
rect 18420 12223 18472 12232
rect 18420 12189 18429 12223
rect 18429 12189 18463 12223
rect 18463 12189 18472 12223
rect 18420 12180 18472 12189
rect 21640 12180 21692 12232
rect 14832 12112 14884 12164
rect 16488 12112 16540 12164
rect 16672 12112 16724 12164
rect 12716 12044 12768 12096
rect 19984 12112 20036 12164
rect 19340 12044 19392 12096
rect 19524 12044 19576 12096
rect 22100 12044 22152 12096
rect 22376 12112 22428 12164
rect 23296 12112 23348 12164
rect 23572 12044 23624 12096
rect 24768 12223 24820 12232
rect 24768 12189 24777 12223
rect 24777 12189 24811 12223
rect 24811 12189 24820 12223
rect 24768 12180 24820 12189
rect 26332 12223 26384 12232
rect 26332 12189 26341 12223
rect 26341 12189 26375 12223
rect 26375 12189 26384 12223
rect 26332 12180 26384 12189
rect 28356 12223 28408 12232
rect 28356 12189 28365 12223
rect 28365 12189 28399 12223
rect 28399 12189 28408 12223
rect 28356 12180 28408 12189
rect 30472 12180 30524 12232
rect 25136 12112 25188 12164
rect 24492 12044 24544 12096
rect 28264 12112 28316 12164
rect 25320 12044 25372 12096
rect 29460 12044 29512 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 10416 11840 10468 11892
rect 10784 11840 10836 11892
rect 8208 11772 8260 11824
rect 11520 11772 11572 11824
rect 11888 11772 11940 11824
rect 12440 11772 12492 11824
rect 10324 11704 10376 11756
rect 10692 11704 10744 11756
rect 11060 11704 11112 11756
rect 10416 11636 10468 11688
rect 11152 11636 11204 11688
rect 14556 11840 14608 11892
rect 15752 11840 15804 11892
rect 16488 11840 16540 11892
rect 18236 11840 18288 11892
rect 19340 11840 19392 11892
rect 22376 11883 22428 11892
rect 17408 11815 17460 11824
rect 17408 11781 17417 11815
rect 17417 11781 17451 11815
rect 17451 11781 17460 11815
rect 17408 11772 17460 11781
rect 17868 11772 17920 11824
rect 18972 11772 19024 11824
rect 21180 11772 21232 11824
rect 22376 11849 22385 11883
rect 22385 11849 22419 11883
rect 22419 11849 22428 11883
rect 22376 11840 22428 11849
rect 24768 11883 24820 11892
rect 23296 11815 23348 11824
rect 23296 11781 23305 11815
rect 23305 11781 23339 11815
rect 23339 11781 23348 11815
rect 23296 11772 23348 11781
rect 23388 11772 23440 11824
rect 24768 11849 24777 11883
rect 24777 11849 24811 11883
rect 24811 11849 24820 11883
rect 24768 11840 24820 11849
rect 26332 11840 26384 11892
rect 30472 11883 30524 11892
rect 30472 11849 30481 11883
rect 30481 11849 30515 11883
rect 30515 11849 30524 11883
rect 30472 11840 30524 11849
rect 30840 11840 30892 11892
rect 25504 11815 25556 11824
rect 16580 11704 16632 11756
rect 19432 11747 19484 11756
rect 19432 11713 19441 11747
rect 19441 11713 19475 11747
rect 19475 11713 19484 11747
rect 19432 11704 19484 11713
rect 14004 11679 14056 11688
rect 14004 11645 14013 11679
rect 14013 11645 14047 11679
rect 14047 11645 14056 11679
rect 14004 11636 14056 11645
rect 16672 11636 16724 11688
rect 21088 11704 21140 11756
rect 9220 11568 9272 11620
rect 9864 11568 9916 11620
rect 18880 11568 18932 11620
rect 5632 11500 5684 11552
rect 10968 11500 11020 11552
rect 11244 11500 11296 11552
rect 13360 11500 13412 11552
rect 17132 11500 17184 11552
rect 18972 11500 19024 11552
rect 25504 11781 25513 11815
rect 25513 11781 25547 11815
rect 25547 11781 25556 11815
rect 25504 11772 25556 11781
rect 26792 11772 26844 11824
rect 27896 11772 27948 11824
rect 29368 11815 29420 11824
rect 29368 11781 29377 11815
rect 29377 11781 29411 11815
rect 29411 11781 29420 11815
rect 29368 11772 29420 11781
rect 29460 11815 29512 11824
rect 29460 11781 29469 11815
rect 29469 11781 29503 11815
rect 29503 11781 29512 11815
rect 29460 11772 29512 11781
rect 30656 11747 30708 11756
rect 30656 11713 30665 11747
rect 30665 11713 30699 11747
rect 30699 11713 30708 11747
rect 30656 11704 30708 11713
rect 34060 11704 34112 11756
rect 22284 11568 22336 11620
rect 23664 11636 23716 11688
rect 24216 11679 24268 11688
rect 24216 11645 24225 11679
rect 24225 11645 24259 11679
rect 24259 11645 24268 11679
rect 24216 11636 24268 11645
rect 24676 11568 24728 11620
rect 26240 11636 26292 11688
rect 27620 11679 27672 11688
rect 27620 11645 27629 11679
rect 27629 11645 27663 11679
rect 27663 11645 27672 11679
rect 27620 11636 27672 11645
rect 28356 11500 28408 11552
rect 29920 11500 29972 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 1768 11135 1820 11144
rect 1768 11101 1777 11135
rect 1777 11101 1811 11135
rect 1811 11101 1820 11135
rect 1768 11092 1820 11101
rect 5724 11296 5776 11348
rect 6460 11228 6512 11280
rect 8484 11296 8536 11348
rect 11152 11296 11204 11348
rect 8668 11228 8720 11280
rect 9496 11228 9548 11280
rect 12992 11228 13044 11280
rect 13360 11228 13412 11280
rect 22100 11296 22152 11348
rect 23204 11339 23256 11348
rect 14096 11228 14148 11280
rect 18880 11228 18932 11280
rect 22284 11228 22336 11280
rect 23204 11305 23213 11339
rect 23213 11305 23247 11339
rect 23247 11305 23256 11339
rect 23204 11296 23256 11305
rect 23848 11339 23900 11348
rect 23848 11305 23857 11339
rect 23857 11305 23891 11339
rect 23891 11305 23900 11339
rect 23848 11296 23900 11305
rect 27896 11339 27948 11348
rect 27896 11305 27905 11339
rect 27905 11305 27939 11339
rect 27939 11305 27948 11339
rect 27896 11296 27948 11305
rect 23572 11228 23624 11280
rect 25136 11228 25188 11280
rect 27804 11228 27856 11280
rect 38200 11271 38252 11280
rect 38200 11237 38209 11271
rect 38209 11237 38243 11271
rect 38243 11237 38252 11271
rect 38200 11228 38252 11237
rect 6736 11160 6788 11212
rect 6000 11024 6052 11076
rect 6552 11024 6604 11076
rect 2320 10999 2372 11008
rect 2320 10965 2329 10999
rect 2329 10965 2363 10999
rect 2363 10965 2372 10999
rect 2320 10956 2372 10965
rect 8944 11024 8996 11076
rect 10784 11160 10836 11212
rect 11704 11203 11756 11212
rect 11704 11169 11713 11203
rect 11713 11169 11747 11203
rect 11747 11169 11756 11203
rect 11704 11160 11756 11169
rect 12532 11160 12584 11212
rect 16580 11160 16632 11212
rect 16672 11160 16724 11212
rect 18052 11160 18104 11212
rect 18236 11160 18288 11212
rect 18512 11203 18564 11212
rect 18512 11169 18521 11203
rect 18521 11169 18555 11203
rect 18555 11169 18564 11203
rect 18512 11160 18564 11169
rect 18788 11160 18840 11212
rect 19248 11160 19300 11212
rect 19432 11160 19484 11212
rect 21548 11160 21600 11212
rect 26240 11203 26292 11212
rect 9496 11135 9548 11144
rect 9496 11101 9505 11135
rect 9505 11101 9539 11135
rect 9539 11101 9548 11135
rect 9496 11092 9548 11101
rect 10876 11092 10928 11144
rect 18604 11092 18656 11144
rect 23020 11092 23072 11144
rect 7380 10956 7432 11008
rect 8116 10956 8168 11008
rect 9680 11024 9732 11076
rect 11980 11024 12032 11076
rect 13360 11024 13412 11076
rect 14004 11024 14056 11076
rect 14556 11067 14608 11076
rect 14556 11033 14565 11067
rect 14565 11033 14599 11067
rect 14599 11033 14608 11067
rect 14556 11024 14608 11033
rect 14832 11024 14884 11076
rect 16304 11067 16356 11076
rect 16304 11033 16313 11067
rect 16313 11033 16347 11067
rect 16347 11033 16356 11067
rect 16304 11024 16356 11033
rect 17040 11024 17092 11076
rect 18328 11024 18380 11076
rect 19432 11067 19484 11076
rect 11520 10956 11572 11008
rect 19432 11033 19441 11067
rect 19441 11033 19475 11067
rect 19475 11033 19484 11067
rect 19432 11024 19484 11033
rect 22008 11024 22060 11076
rect 24216 11092 24268 11144
rect 26240 11169 26249 11203
rect 26249 11169 26283 11203
rect 26283 11169 26292 11203
rect 26240 11160 26292 11169
rect 28448 11203 28500 11212
rect 28448 11169 28457 11203
rect 28457 11169 28491 11203
rect 28491 11169 28500 11203
rect 28448 11160 28500 11169
rect 30656 11160 30708 11212
rect 29276 11092 29328 11144
rect 29920 11135 29972 11144
rect 29920 11101 29929 11135
rect 29929 11101 29963 11135
rect 29963 11101 29972 11135
rect 29920 11092 29972 11101
rect 37372 11135 37424 11144
rect 37372 11101 37381 11135
rect 37381 11101 37415 11135
rect 37415 11101 37424 11135
rect 37372 11092 37424 11101
rect 25136 11067 25188 11076
rect 25136 11033 25145 11067
rect 25145 11033 25179 11067
rect 25179 11033 25188 11067
rect 25136 11024 25188 11033
rect 25320 11024 25372 11076
rect 25412 11024 25464 11076
rect 25872 11024 25924 11076
rect 29092 11067 29144 11076
rect 29092 11033 29101 11067
rect 29101 11033 29135 11067
rect 29135 11033 29144 11067
rect 29092 11024 29144 11033
rect 36912 11024 36964 11076
rect 29000 10956 29052 11008
rect 29460 10956 29512 11008
rect 37464 10999 37516 11008
rect 37464 10965 37473 10999
rect 37473 10965 37507 10999
rect 37507 10965 37516 10999
rect 37464 10956 37516 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 1952 10752 2004 10804
rect 4804 10752 4856 10804
rect 7380 10752 7432 10804
rect 7932 10752 7984 10804
rect 10876 10752 10928 10804
rect 12348 10752 12400 10804
rect 12624 10752 12676 10804
rect 7472 10684 7524 10736
rect 1768 10659 1820 10668
rect 1768 10625 1777 10659
rect 1777 10625 1811 10659
rect 1811 10625 1820 10659
rect 1768 10616 1820 10625
rect 2780 10616 2832 10668
rect 1952 10548 2004 10600
rect 4804 10616 4856 10668
rect 6828 10548 6880 10600
rect 10324 10684 10376 10736
rect 10508 10684 10560 10736
rect 10692 10684 10744 10736
rect 15200 10752 15252 10804
rect 16028 10752 16080 10804
rect 10232 10616 10284 10668
rect 10784 10659 10836 10668
rect 10784 10625 10793 10659
rect 10793 10625 10827 10659
rect 10827 10625 10836 10659
rect 10784 10616 10836 10625
rect 11980 10616 12032 10668
rect 15292 10684 15344 10736
rect 17960 10684 18012 10736
rect 18604 10752 18656 10804
rect 19340 10752 19392 10804
rect 20260 10752 20312 10804
rect 20444 10752 20496 10804
rect 12532 10616 12584 10668
rect 13360 10659 13412 10668
rect 11428 10548 11480 10600
rect 11704 10548 11756 10600
rect 13360 10625 13369 10659
rect 13369 10625 13403 10659
rect 13403 10625 13412 10659
rect 13360 10616 13412 10625
rect 15844 10616 15896 10668
rect 16120 10616 16172 10668
rect 8576 10480 8628 10532
rect 9864 10412 9916 10464
rect 10324 10412 10376 10464
rect 12716 10412 12768 10464
rect 16948 10591 17000 10600
rect 13728 10412 13780 10464
rect 16948 10557 16957 10591
rect 16957 10557 16991 10591
rect 16991 10557 17000 10591
rect 16948 10548 17000 10557
rect 17868 10548 17920 10600
rect 19984 10684 20036 10736
rect 19248 10659 19300 10668
rect 19248 10625 19257 10659
rect 19257 10625 19291 10659
rect 19291 10625 19300 10659
rect 19248 10616 19300 10625
rect 18788 10548 18840 10600
rect 19616 10548 19668 10600
rect 21824 10548 21876 10600
rect 18236 10480 18288 10532
rect 25504 10752 25556 10804
rect 29276 10795 29328 10804
rect 29276 10761 29285 10795
rect 29285 10761 29319 10795
rect 29319 10761 29328 10795
rect 29276 10752 29328 10761
rect 36912 10752 36964 10804
rect 23756 10727 23808 10736
rect 23756 10693 23765 10727
rect 23765 10693 23799 10727
rect 23799 10693 23808 10727
rect 23756 10684 23808 10693
rect 25964 10684 26016 10736
rect 31760 10684 31812 10736
rect 22560 10659 22612 10668
rect 22560 10625 22569 10659
rect 22569 10625 22603 10659
rect 22603 10625 22612 10659
rect 22560 10616 22612 10625
rect 29460 10659 29512 10668
rect 23480 10548 23532 10600
rect 23848 10548 23900 10600
rect 16120 10412 16172 10464
rect 17684 10412 17736 10464
rect 24952 10480 25004 10532
rect 21916 10412 21968 10464
rect 22836 10412 22888 10464
rect 29460 10625 29469 10659
rect 29469 10625 29503 10659
rect 29503 10625 29512 10659
rect 29460 10616 29512 10625
rect 34520 10659 34572 10668
rect 34520 10625 34529 10659
rect 34529 10625 34563 10659
rect 34563 10625 34572 10659
rect 34520 10616 34572 10625
rect 38016 10659 38068 10668
rect 33140 10548 33192 10600
rect 38016 10625 38025 10659
rect 38025 10625 38059 10659
rect 38059 10625 38068 10659
rect 38016 10616 38068 10625
rect 35532 10412 35584 10464
rect 38200 10455 38252 10464
rect 38200 10421 38209 10455
rect 38209 10421 38243 10455
rect 38243 10421 38252 10455
rect 38200 10412 38252 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 6460 10140 6512 10192
rect 9036 10208 9088 10260
rect 11336 10208 11388 10260
rect 11704 10208 11756 10260
rect 16028 10208 16080 10260
rect 11520 10140 11572 10192
rect 13636 10183 13688 10192
rect 13636 10149 13645 10183
rect 13645 10149 13679 10183
rect 13679 10149 13688 10183
rect 13636 10140 13688 10149
rect 13728 10140 13780 10192
rect 17316 10140 17368 10192
rect 5540 10072 5592 10124
rect 2780 10004 2832 10056
rect 4804 10004 4856 10056
rect 4988 10004 5040 10056
rect 5448 10004 5500 10056
rect 5816 10004 5868 10056
rect 6552 10004 6604 10056
rect 6828 10047 6880 10056
rect 6828 10013 6837 10047
rect 6837 10013 6871 10047
rect 6871 10013 6880 10047
rect 6828 10004 6880 10013
rect 8576 10004 8628 10056
rect 9496 10004 9548 10056
rect 11888 10047 11940 10056
rect 11888 10013 11897 10047
rect 11897 10013 11931 10047
rect 11931 10013 11940 10047
rect 11888 10004 11940 10013
rect 3884 9936 3936 9988
rect 5724 9936 5776 9988
rect 6092 9936 6144 9988
rect 7012 9936 7064 9988
rect 9956 9979 10008 9988
rect 9956 9945 9965 9979
rect 9965 9945 9999 9979
rect 9999 9945 10008 9979
rect 9956 9936 10008 9945
rect 10232 9936 10284 9988
rect 4988 9868 5040 9920
rect 5356 9868 5408 9920
rect 9772 9868 9824 9920
rect 12624 9936 12676 9988
rect 15108 10072 15160 10124
rect 16304 10072 16356 10124
rect 16856 10072 16908 10124
rect 15476 10004 15528 10056
rect 17868 10072 17920 10124
rect 18236 10140 18288 10192
rect 19616 10140 19668 10192
rect 23296 10208 23348 10260
rect 38016 10208 38068 10260
rect 24032 10140 24084 10192
rect 15200 9936 15252 9988
rect 13912 9868 13964 9920
rect 15292 9868 15344 9920
rect 17592 9936 17644 9988
rect 18972 10072 19024 10124
rect 20168 10072 20220 10124
rect 20536 10072 20588 10124
rect 21824 10072 21876 10124
rect 24676 10115 24728 10124
rect 19340 10004 19392 10056
rect 24676 10081 24685 10115
rect 24685 10081 24719 10115
rect 24719 10081 24728 10115
rect 24676 10072 24728 10081
rect 37464 10004 37516 10056
rect 19984 9936 20036 9988
rect 20168 9936 20220 9988
rect 22744 9936 22796 9988
rect 24768 9979 24820 9988
rect 24768 9945 24777 9979
rect 24777 9945 24811 9979
rect 24811 9945 24820 9979
rect 24768 9936 24820 9945
rect 25964 9936 26016 9988
rect 18972 9868 19024 9920
rect 27160 9868 27212 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 4528 9707 4580 9716
rect 4528 9673 4537 9707
rect 4537 9673 4571 9707
rect 4571 9673 4580 9707
rect 4528 9664 4580 9673
rect 4804 9664 4856 9716
rect 2228 9596 2280 9648
rect 5540 9664 5592 9716
rect 9036 9664 9088 9716
rect 9588 9664 9640 9716
rect 12532 9664 12584 9716
rect 2136 9528 2188 9580
rect 2596 9528 2648 9580
rect 3240 9571 3292 9580
rect 3240 9537 3249 9571
rect 3249 9537 3283 9571
rect 3283 9537 3292 9571
rect 3240 9528 3292 9537
rect 3884 9571 3936 9580
rect 3884 9537 3893 9571
rect 3893 9537 3927 9571
rect 3927 9537 3936 9571
rect 3884 9528 3936 9537
rect 4252 9528 4304 9580
rect 9496 9596 9548 9648
rect 13636 9664 13688 9716
rect 15384 9664 15436 9716
rect 22560 9664 22612 9716
rect 10140 9528 10192 9580
rect 3792 9460 3844 9512
rect 4160 9460 4212 9512
rect 6828 9460 6880 9512
rect 13084 9596 13136 9648
rect 14372 9596 14424 9648
rect 14740 9596 14792 9648
rect 15476 9639 15528 9648
rect 15476 9605 15485 9639
rect 15485 9605 15519 9639
rect 15519 9605 15528 9639
rect 15476 9596 15528 9605
rect 12256 9528 12308 9580
rect 14648 9571 14700 9580
rect 14648 9537 14657 9571
rect 14657 9537 14691 9571
rect 14691 9537 14700 9571
rect 14648 9528 14700 9537
rect 15016 9528 15068 9580
rect 17776 9596 17828 9648
rect 19156 9596 19208 9648
rect 23664 9596 23716 9648
rect 33140 9596 33192 9648
rect 16028 9571 16080 9580
rect 16028 9537 16037 9571
rect 16037 9537 16071 9571
rect 16071 9537 16080 9571
rect 16028 9528 16080 9537
rect 16948 9528 17000 9580
rect 11888 9460 11940 9512
rect 12348 9503 12400 9512
rect 12348 9469 12357 9503
rect 12357 9469 12391 9503
rect 12391 9469 12400 9503
rect 12348 9460 12400 9469
rect 16212 9460 16264 9512
rect 18512 9460 18564 9512
rect 18972 9503 19024 9512
rect 18972 9469 18981 9503
rect 18981 9469 19015 9503
rect 19015 9469 19024 9503
rect 18972 9460 19024 9469
rect 19340 9460 19392 9512
rect 20720 9460 20772 9512
rect 21088 9460 21140 9512
rect 3332 9435 3384 9444
rect 3332 9401 3341 9435
rect 3341 9401 3375 9435
rect 3375 9401 3384 9435
rect 3332 9392 3384 9401
rect 5632 9392 5684 9444
rect 5816 9324 5868 9376
rect 6920 9324 6972 9376
rect 9312 9324 9364 9376
rect 15108 9392 15160 9444
rect 30380 9528 30432 9580
rect 30840 9528 30892 9580
rect 23940 9460 23992 9512
rect 24032 9503 24084 9512
rect 24032 9469 24041 9503
rect 24041 9469 24075 9503
rect 24075 9469 24084 9503
rect 24032 9460 24084 9469
rect 29276 9460 29328 9512
rect 25780 9392 25832 9444
rect 14096 9367 14148 9376
rect 14096 9333 14105 9367
rect 14105 9333 14139 9367
rect 14139 9333 14148 9367
rect 14096 9324 14148 9333
rect 15016 9324 15068 9376
rect 19248 9324 19300 9376
rect 20904 9324 20956 9376
rect 29460 9324 29512 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 2320 9120 2372 9172
rect 2596 9052 2648 9104
rect 2964 8916 3016 8968
rect 3240 8959 3292 8968
rect 3240 8925 3249 8959
rect 3249 8925 3283 8959
rect 3283 8925 3292 8959
rect 3240 8916 3292 8925
rect 4528 9120 4580 9172
rect 6920 9120 6972 9172
rect 7840 9120 7892 9172
rect 8392 9052 8444 9104
rect 8852 9052 8904 9104
rect 10600 9120 10652 9172
rect 14096 9120 14148 9172
rect 14280 9120 14332 9172
rect 1768 8823 1820 8832
rect 1768 8789 1777 8823
rect 1777 8789 1811 8823
rect 1811 8789 1820 8823
rect 1768 8780 1820 8789
rect 2872 8780 2924 8832
rect 4620 8848 4672 8900
rect 4804 8823 4856 8832
rect 4804 8789 4813 8823
rect 4813 8789 4847 8823
rect 4847 8789 4856 8823
rect 13912 9052 13964 9104
rect 16488 9120 16540 9172
rect 21364 9120 21416 9172
rect 22744 9120 22796 9172
rect 23664 9163 23716 9172
rect 23664 9129 23673 9163
rect 23673 9129 23707 9163
rect 23707 9129 23716 9163
rect 23664 9120 23716 9129
rect 9404 9027 9456 9036
rect 9404 8993 9413 9027
rect 9413 8993 9447 9027
rect 9447 8993 9456 9027
rect 9404 8984 9456 8993
rect 9496 8984 9548 9036
rect 11244 8984 11296 9036
rect 12348 8984 12400 9036
rect 12900 8984 12952 9036
rect 15384 8984 15436 9036
rect 16856 8984 16908 9036
rect 19340 8984 19392 9036
rect 20904 9052 20956 9104
rect 25688 9052 25740 9104
rect 20260 8984 20312 9036
rect 20352 8984 20404 9036
rect 5172 8916 5224 8968
rect 6828 8959 6880 8968
rect 5264 8848 5316 8900
rect 6276 8891 6328 8900
rect 4804 8780 4856 8789
rect 5172 8780 5224 8832
rect 6276 8857 6285 8891
rect 6285 8857 6319 8891
rect 6319 8857 6328 8891
rect 6276 8848 6328 8857
rect 6828 8925 6837 8959
rect 6837 8925 6871 8959
rect 6871 8925 6880 8959
rect 6828 8916 6880 8925
rect 8484 8916 8536 8968
rect 8852 8916 8904 8968
rect 12716 8916 12768 8968
rect 16580 8959 16632 8968
rect 16580 8925 16589 8959
rect 16589 8925 16623 8959
rect 16623 8925 16632 8959
rect 16580 8916 16632 8925
rect 19248 8916 19300 8968
rect 7196 8780 7248 8832
rect 7748 8780 7800 8832
rect 9312 8848 9364 8900
rect 9404 8848 9456 8900
rect 9588 8780 9640 8832
rect 9772 8780 9824 8832
rect 10876 8780 10928 8832
rect 14188 8848 14240 8900
rect 15108 8848 15160 8900
rect 17960 8891 18012 8900
rect 17960 8857 17969 8891
rect 17969 8857 18003 8891
rect 18003 8857 18012 8891
rect 17960 8848 18012 8857
rect 19432 8848 19484 8900
rect 21732 8916 21784 8968
rect 21180 8848 21232 8900
rect 12992 8780 13044 8832
rect 13176 8780 13228 8832
rect 16672 8823 16724 8832
rect 16672 8789 16681 8823
rect 16681 8789 16715 8823
rect 16715 8789 16724 8823
rect 16672 8780 16724 8789
rect 20628 8780 20680 8832
rect 20720 8780 20772 8832
rect 21824 8780 21876 8832
rect 23020 8916 23072 8968
rect 23480 8916 23532 8968
rect 29092 8916 29144 8968
rect 30840 8959 30892 8968
rect 24952 8891 25004 8900
rect 24952 8857 24961 8891
rect 24961 8857 24995 8891
rect 24995 8857 25004 8891
rect 24952 8848 25004 8857
rect 25044 8891 25096 8900
rect 25044 8857 25053 8891
rect 25053 8857 25087 8891
rect 25087 8857 25096 8891
rect 25964 8891 26016 8900
rect 25044 8848 25096 8857
rect 25964 8857 25973 8891
rect 25973 8857 26007 8891
rect 26007 8857 26016 8891
rect 25964 8848 26016 8857
rect 26700 8848 26752 8900
rect 30840 8925 30849 8959
rect 30849 8925 30883 8959
rect 30883 8925 30892 8959
rect 30840 8916 30892 8925
rect 38292 8959 38344 8968
rect 38292 8925 38301 8959
rect 38301 8925 38335 8959
rect 38335 8925 38344 8959
rect 38292 8916 38344 8925
rect 25596 8780 25648 8832
rect 25688 8780 25740 8832
rect 30196 8780 30248 8832
rect 30380 8823 30432 8832
rect 30380 8789 30389 8823
rect 30389 8789 30423 8823
rect 30423 8789 30432 8823
rect 30380 8780 30432 8789
rect 38108 8823 38160 8832
rect 38108 8789 38117 8823
rect 38117 8789 38151 8823
rect 38151 8789 38160 8823
rect 38108 8780 38160 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 1860 8576 1912 8628
rect 2228 8619 2280 8628
rect 2228 8585 2237 8619
rect 2237 8585 2271 8619
rect 2271 8585 2280 8619
rect 2228 8576 2280 8585
rect 1400 8440 1452 8492
rect 1860 8440 1912 8492
rect 3056 8483 3108 8492
rect 3056 8449 3065 8483
rect 3065 8449 3099 8483
rect 3099 8449 3108 8483
rect 3056 8440 3108 8449
rect 3884 8440 3936 8492
rect 6828 8576 6880 8628
rect 4528 8551 4580 8560
rect 4528 8517 4537 8551
rect 4537 8517 4571 8551
rect 4571 8517 4580 8551
rect 4528 8508 4580 8517
rect 5540 8508 5592 8560
rect 6644 8551 6696 8560
rect 6644 8517 6653 8551
rect 6653 8517 6687 8551
rect 6687 8517 6696 8551
rect 6644 8508 6696 8517
rect 10140 8576 10192 8628
rect 13360 8576 13412 8628
rect 14648 8576 14700 8628
rect 7196 8483 7248 8492
rect 7196 8449 7205 8483
rect 7205 8449 7239 8483
rect 7239 8449 7248 8483
rect 9312 8508 9364 8560
rect 12348 8551 12400 8560
rect 12348 8517 12357 8551
rect 12357 8517 12391 8551
rect 12391 8517 12400 8551
rect 12348 8508 12400 8517
rect 13176 8551 13228 8560
rect 13176 8517 13185 8551
rect 13185 8517 13219 8551
rect 13219 8517 13228 8551
rect 13176 8508 13228 8517
rect 13636 8508 13688 8560
rect 15108 8508 15160 8560
rect 17960 8576 18012 8628
rect 17132 8551 17184 8560
rect 17132 8517 17141 8551
rect 17141 8517 17175 8551
rect 17175 8517 17184 8551
rect 17132 8508 17184 8517
rect 7196 8440 7248 8449
rect 10232 8440 10284 8492
rect 10508 8440 10560 8492
rect 10968 8483 11020 8492
rect 10968 8449 10977 8483
rect 10977 8449 11011 8483
rect 11011 8449 11020 8483
rect 10968 8440 11020 8449
rect 12256 8483 12308 8492
rect 12256 8449 12265 8483
rect 12265 8449 12299 8483
rect 12299 8449 12308 8483
rect 12256 8440 12308 8449
rect 12900 8483 12952 8492
rect 12900 8449 12909 8483
rect 12909 8449 12943 8483
rect 12943 8449 12952 8483
rect 12900 8440 12952 8449
rect 16856 8483 16908 8492
rect 16856 8449 16865 8483
rect 16865 8449 16899 8483
rect 16899 8449 16908 8483
rect 16856 8440 16908 8449
rect 19340 8508 19392 8560
rect 20996 8508 21048 8560
rect 21180 8576 21232 8628
rect 23572 8576 23624 8628
rect 24032 8576 24084 8628
rect 25044 8619 25096 8628
rect 25044 8585 25053 8619
rect 25053 8585 25087 8619
rect 25087 8585 25096 8619
rect 25044 8576 25096 8585
rect 26608 8576 26660 8628
rect 30380 8576 30432 8628
rect 24124 8508 24176 8560
rect 7104 8372 7156 8424
rect 7564 8372 7616 8424
rect 8576 8415 8628 8424
rect 8576 8381 8585 8415
rect 8585 8381 8619 8415
rect 8619 8381 8628 8415
rect 8576 8372 8628 8381
rect 8852 8415 8904 8424
rect 8852 8381 8861 8415
rect 8861 8381 8895 8415
rect 8895 8381 8904 8415
rect 8852 8372 8904 8381
rect 8944 8372 8996 8424
rect 12440 8372 12492 8424
rect 16120 8415 16172 8424
rect 16120 8381 16129 8415
rect 16129 8381 16163 8415
rect 16163 8381 16172 8415
rect 16120 8372 16172 8381
rect 20076 8372 20128 8424
rect 21364 8440 21416 8492
rect 23664 8483 23716 8492
rect 23664 8449 23673 8483
rect 23673 8449 23707 8483
rect 23707 8449 23716 8483
rect 23664 8440 23716 8449
rect 24216 8440 24268 8492
rect 8484 8304 8536 8356
rect 10140 8304 10192 8356
rect 12900 8304 12952 8356
rect 3976 8236 4028 8288
rect 6828 8236 6880 8288
rect 8024 8236 8076 8288
rect 8944 8236 8996 8288
rect 10048 8236 10100 8288
rect 10600 8236 10652 8288
rect 14556 8236 14608 8288
rect 15844 8236 15896 8288
rect 20444 8304 20496 8356
rect 23388 8372 23440 8424
rect 20352 8236 20404 8288
rect 21272 8304 21324 8356
rect 25964 8440 26016 8492
rect 27344 8483 27396 8492
rect 27344 8449 27353 8483
rect 27353 8449 27387 8483
rect 27387 8449 27396 8483
rect 27344 8440 27396 8449
rect 28448 8483 28500 8492
rect 28448 8449 28457 8483
rect 28457 8449 28491 8483
rect 28491 8449 28500 8483
rect 28448 8440 28500 8449
rect 29276 8483 29328 8492
rect 29276 8449 29285 8483
rect 29285 8449 29319 8483
rect 29319 8449 29328 8483
rect 29276 8440 29328 8449
rect 29460 8483 29512 8492
rect 29460 8449 29469 8483
rect 29469 8449 29503 8483
rect 29503 8449 29512 8483
rect 29460 8440 29512 8449
rect 38108 8440 38160 8492
rect 27712 8304 27764 8356
rect 28632 8347 28684 8356
rect 28632 8313 28641 8347
rect 28641 8313 28675 8347
rect 28675 8313 28684 8347
rect 28632 8304 28684 8313
rect 30472 8347 30524 8356
rect 30472 8313 30481 8347
rect 30481 8313 30515 8347
rect 30515 8313 30524 8347
rect 30472 8304 30524 8313
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 1952 8075 2004 8084
rect 1952 8041 1961 8075
rect 1961 8041 1995 8075
rect 1995 8041 2004 8075
rect 1952 8032 2004 8041
rect 5540 8032 5592 8084
rect 7380 8032 7432 8084
rect 4068 8007 4120 8016
rect 4068 7973 4077 8007
rect 4077 7973 4111 8007
rect 4111 7973 4120 8007
rect 4068 7964 4120 7973
rect 5908 7964 5960 8016
rect 1584 7828 1636 7880
rect 3608 7896 3660 7948
rect 6276 7896 6328 7948
rect 6736 7939 6788 7948
rect 6736 7905 6745 7939
rect 6745 7905 6779 7939
rect 6779 7905 6788 7939
rect 6736 7896 6788 7905
rect 8668 7964 8720 8016
rect 10600 7964 10652 8016
rect 16764 8032 16816 8084
rect 19064 8032 19116 8084
rect 20996 8032 21048 8084
rect 23756 8032 23808 8084
rect 14556 7964 14608 8016
rect 3976 7871 4028 7880
rect 3976 7837 3985 7871
rect 3985 7837 4019 7871
rect 4019 7837 4028 7871
rect 3976 7828 4028 7837
rect 4620 7760 4672 7812
rect 5080 7828 5132 7880
rect 6552 7828 6604 7880
rect 8576 7896 8628 7948
rect 14096 7896 14148 7948
rect 14188 7896 14240 7948
rect 16120 7896 16172 7948
rect 16856 7896 16908 7948
rect 18696 7964 18748 8016
rect 21548 7964 21600 8016
rect 21824 7964 21876 8016
rect 24768 8032 24820 8084
rect 25964 8032 26016 8084
rect 8760 7828 8812 7880
rect 10968 7828 11020 7880
rect 3148 7692 3200 7744
rect 3424 7692 3476 7744
rect 6920 7760 6972 7812
rect 7104 7760 7156 7812
rect 7472 7760 7524 7812
rect 8300 7760 8352 7812
rect 12900 7828 12952 7880
rect 13360 7828 13412 7880
rect 19984 7871 20036 7880
rect 19984 7837 19993 7871
rect 19993 7837 20027 7871
rect 20027 7837 20036 7871
rect 19984 7828 20036 7837
rect 22376 7828 22428 7880
rect 23664 7828 23716 7880
rect 29000 7964 29052 8016
rect 31668 7964 31720 8016
rect 24216 7896 24268 7948
rect 24768 7896 24820 7948
rect 27252 7939 27304 7948
rect 24492 7828 24544 7880
rect 5356 7692 5408 7744
rect 6092 7735 6144 7744
rect 6092 7701 6101 7735
rect 6101 7701 6135 7735
rect 6135 7701 6144 7735
rect 6092 7692 6144 7701
rect 7656 7692 7708 7744
rect 16672 7760 16724 7812
rect 16304 7692 16356 7744
rect 22008 7760 22060 7812
rect 22928 7760 22980 7812
rect 21272 7692 21324 7744
rect 21548 7692 21600 7744
rect 24952 7828 25004 7880
rect 27252 7905 27261 7939
rect 27261 7905 27295 7939
rect 27295 7905 27304 7939
rect 27252 7896 27304 7905
rect 37464 7871 37516 7880
rect 37464 7837 37473 7871
rect 37473 7837 37507 7871
rect 37507 7837 37516 7871
rect 37464 7828 37516 7837
rect 26240 7803 26292 7812
rect 26240 7769 26249 7803
rect 26249 7769 26283 7803
rect 26283 7769 26292 7803
rect 26240 7760 26292 7769
rect 27436 7692 27488 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 2504 7488 2556 7540
rect 2688 7488 2740 7540
rect 4712 7420 4764 7472
rect 3700 7352 3752 7404
rect 5356 7420 5408 7472
rect 1952 7327 2004 7336
rect 1952 7293 1961 7327
rect 1961 7293 1995 7327
rect 1995 7293 2004 7327
rect 1952 7284 2004 7293
rect 2136 7327 2188 7336
rect 2136 7293 2145 7327
rect 2145 7293 2179 7327
rect 2179 7293 2188 7327
rect 2136 7284 2188 7293
rect 2228 7284 2280 7336
rect 2596 7284 2648 7336
rect 5080 7352 5132 7404
rect 8024 7488 8076 7540
rect 8760 7488 8812 7540
rect 7840 7420 7892 7472
rect 13176 7488 13228 7540
rect 14280 7488 14332 7540
rect 15844 7488 15896 7540
rect 6736 7352 6788 7404
rect 7380 7327 7432 7336
rect 7380 7293 7389 7327
rect 7389 7293 7423 7327
rect 7423 7293 7432 7327
rect 7380 7284 7432 7293
rect 7932 7284 7984 7336
rect 4528 7216 4580 7268
rect 5080 7216 5132 7268
rect 2780 7148 2832 7200
rect 5448 7148 5500 7200
rect 7104 7148 7156 7200
rect 15200 7420 15252 7472
rect 14188 7395 14240 7404
rect 14188 7361 14197 7395
rect 14197 7361 14231 7395
rect 14231 7361 14240 7395
rect 14188 7352 14240 7361
rect 16488 7352 16540 7404
rect 17224 7352 17276 7404
rect 17776 7463 17828 7472
rect 17776 7429 17785 7463
rect 17785 7429 17819 7463
rect 17819 7429 17828 7463
rect 17776 7420 17828 7429
rect 19984 7488 20036 7540
rect 21364 7420 21416 7472
rect 23388 7488 23440 7540
rect 25780 7531 25832 7540
rect 25780 7497 25789 7531
rect 25789 7497 25823 7531
rect 25823 7497 25832 7531
rect 25780 7488 25832 7497
rect 26240 7488 26292 7540
rect 34060 7488 34112 7540
rect 23112 7420 23164 7472
rect 18880 7352 18932 7404
rect 19708 7395 19760 7404
rect 19708 7361 19717 7395
rect 19717 7361 19751 7395
rect 19751 7361 19760 7395
rect 19708 7352 19760 7361
rect 9312 7327 9364 7336
rect 9312 7293 9321 7327
rect 9321 7293 9355 7327
rect 9355 7293 9364 7327
rect 9312 7284 9364 7293
rect 9680 7284 9732 7336
rect 11612 7284 11664 7336
rect 12164 7327 12216 7336
rect 10968 7148 11020 7200
rect 12164 7293 12173 7327
rect 12173 7293 12207 7327
rect 12207 7293 12216 7327
rect 12164 7284 12216 7293
rect 16212 7284 16264 7336
rect 17776 7284 17828 7336
rect 19616 7284 19668 7336
rect 20352 7284 20404 7336
rect 20628 7284 20680 7336
rect 24768 7352 24820 7404
rect 26240 7352 26292 7404
rect 26516 7352 26568 7404
rect 27896 7352 27948 7404
rect 24216 7327 24268 7336
rect 24216 7293 24225 7327
rect 24225 7293 24259 7327
rect 24259 7293 24268 7327
rect 24216 7284 24268 7293
rect 14188 7216 14240 7268
rect 14096 7148 14148 7200
rect 17500 7216 17552 7268
rect 20996 7216 21048 7268
rect 18144 7148 18196 7200
rect 20168 7148 20220 7200
rect 21088 7148 21140 7200
rect 21916 7216 21968 7268
rect 24952 7284 25004 7336
rect 25780 7284 25832 7336
rect 38292 7395 38344 7404
rect 38292 7361 38301 7395
rect 38301 7361 38335 7395
rect 38335 7361 38344 7395
rect 38292 7352 38344 7361
rect 24492 7216 24544 7268
rect 29552 7216 29604 7268
rect 26240 7148 26292 7200
rect 26332 7148 26384 7200
rect 35808 7148 35860 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 2688 6987 2740 6996
rect 2688 6953 2697 6987
rect 2697 6953 2731 6987
rect 2731 6953 2740 6987
rect 2688 6944 2740 6953
rect 1952 6876 2004 6928
rect 5448 6876 5500 6928
rect 2872 6808 2924 6860
rect 7472 6944 7524 6996
rect 7564 6944 7616 6996
rect 10968 6944 11020 6996
rect 12072 6944 12124 6996
rect 12164 6944 12216 6996
rect 6184 6876 6236 6928
rect 6552 6876 6604 6928
rect 6736 6808 6788 6860
rect 13268 6876 13320 6928
rect 13728 6876 13780 6928
rect 18880 6944 18932 6996
rect 26240 6944 26292 6996
rect 1768 6783 1820 6792
rect 1768 6749 1777 6783
rect 1777 6749 1811 6783
rect 1811 6749 1820 6783
rect 1768 6740 1820 6749
rect 2228 6783 2280 6792
rect 2228 6749 2237 6783
rect 2237 6749 2271 6783
rect 2271 6749 2280 6783
rect 2228 6740 2280 6749
rect 3332 6740 3384 6792
rect 4344 6783 4396 6792
rect 4344 6749 4353 6783
rect 4353 6749 4387 6783
rect 4387 6749 4396 6783
rect 4344 6740 4396 6749
rect 2964 6672 3016 6724
rect 3700 6672 3752 6724
rect 5080 6740 5132 6792
rect 5540 6783 5592 6792
rect 5540 6749 5549 6783
rect 5549 6749 5583 6783
rect 5583 6749 5592 6783
rect 5540 6740 5592 6749
rect 5724 6740 5776 6792
rect 7012 6672 7064 6724
rect 1492 6604 1544 6656
rect 6828 6604 6880 6656
rect 7564 6672 7616 6724
rect 12072 6808 12124 6860
rect 12348 6808 12400 6860
rect 8668 6740 8720 6792
rect 10140 6740 10192 6792
rect 11704 6783 11756 6792
rect 11704 6749 11713 6783
rect 11713 6749 11747 6783
rect 11747 6749 11756 6783
rect 11704 6740 11756 6749
rect 8484 6604 8536 6656
rect 9404 6604 9456 6656
rect 9772 6647 9824 6656
rect 9772 6613 9781 6647
rect 9781 6613 9815 6647
rect 9815 6613 9824 6647
rect 9772 6604 9824 6613
rect 11980 6672 12032 6724
rect 12072 6604 12124 6656
rect 12440 6672 12492 6724
rect 14188 6808 14240 6860
rect 16028 6808 16080 6860
rect 17224 6808 17276 6860
rect 17500 6808 17552 6860
rect 19432 6808 19484 6860
rect 19708 6851 19760 6860
rect 19708 6817 19717 6851
rect 19717 6817 19751 6851
rect 19751 6817 19760 6851
rect 19708 6808 19760 6817
rect 21548 6876 21600 6928
rect 21180 6808 21232 6860
rect 22008 6851 22060 6860
rect 22008 6817 22017 6851
rect 22017 6817 22051 6851
rect 22051 6817 22060 6851
rect 22008 6808 22060 6817
rect 25964 6876 26016 6928
rect 25228 6851 25280 6860
rect 19616 6740 19668 6792
rect 21272 6740 21324 6792
rect 18144 6672 18196 6724
rect 19984 6715 20036 6724
rect 19984 6681 19993 6715
rect 19993 6681 20027 6715
rect 20027 6681 20036 6715
rect 19984 6672 20036 6681
rect 21548 6672 21600 6724
rect 22376 6740 22428 6792
rect 23020 6740 23072 6792
rect 25228 6817 25237 6851
rect 25237 6817 25271 6851
rect 25271 6817 25280 6851
rect 25228 6808 25280 6817
rect 26148 6808 26200 6860
rect 26700 6808 26752 6860
rect 26976 6876 27028 6928
rect 30472 6808 30524 6860
rect 26332 6740 26384 6792
rect 27988 6783 28040 6792
rect 27988 6749 27997 6783
rect 27997 6749 28031 6783
rect 28031 6749 28040 6783
rect 27988 6740 28040 6749
rect 28448 6740 28500 6792
rect 24952 6715 25004 6724
rect 17408 6604 17460 6656
rect 22008 6604 22060 6656
rect 22192 6604 22244 6656
rect 23112 6604 23164 6656
rect 24952 6681 24961 6715
rect 24961 6681 24995 6715
rect 24995 6681 25004 6715
rect 24952 6672 25004 6681
rect 28724 6647 28776 6656
rect 28724 6613 28733 6647
rect 28733 6613 28767 6647
rect 28767 6613 28776 6647
rect 28724 6604 28776 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 5908 6443 5960 6452
rect 5908 6409 5917 6443
rect 5917 6409 5951 6443
rect 5951 6409 5960 6443
rect 5908 6400 5960 6409
rect 2964 6375 3016 6384
rect 2964 6341 2973 6375
rect 2973 6341 3007 6375
rect 3007 6341 3016 6375
rect 2964 6332 3016 6341
rect 4068 6332 4120 6384
rect 9956 6400 10008 6452
rect 7104 6332 7156 6384
rect 8116 6375 8168 6384
rect 8116 6341 8125 6375
rect 8125 6341 8159 6375
rect 8159 6341 8168 6375
rect 8116 6332 8168 6341
rect 2228 6196 2280 6248
rect 5540 6264 5592 6316
rect 5724 6264 5776 6316
rect 7104 6196 7156 6248
rect 8024 6307 8076 6316
rect 8024 6273 8033 6307
rect 8033 6273 8067 6307
rect 8067 6273 8076 6307
rect 8024 6264 8076 6273
rect 8576 6264 8628 6316
rect 9220 6332 9272 6384
rect 9404 6332 9456 6384
rect 12716 6400 12768 6452
rect 10324 6332 10376 6384
rect 12440 6332 12492 6384
rect 10784 6264 10836 6316
rect 8484 6128 8536 6180
rect 8668 6128 8720 6180
rect 6552 6060 6604 6112
rect 9956 6128 10008 6180
rect 11520 6196 11572 6248
rect 11704 6239 11756 6248
rect 11704 6205 11713 6239
rect 11713 6205 11747 6239
rect 11747 6205 11756 6239
rect 11704 6196 11756 6205
rect 15200 6400 15252 6452
rect 16764 6400 16816 6452
rect 14188 6332 14240 6384
rect 14372 6332 14424 6384
rect 15292 6332 15344 6384
rect 19064 6400 19116 6452
rect 19340 6400 19392 6452
rect 20260 6400 20312 6452
rect 23388 6400 23440 6452
rect 22008 6332 22060 6384
rect 23020 6332 23072 6384
rect 24032 6332 24084 6384
rect 25320 6375 25372 6384
rect 25320 6341 25329 6375
rect 25329 6341 25363 6375
rect 25363 6341 25372 6375
rect 25320 6332 25372 6341
rect 27528 6332 27580 6384
rect 27804 6400 27856 6452
rect 31484 6332 31536 6384
rect 17224 6307 17276 6316
rect 17224 6273 17233 6307
rect 17233 6273 17267 6307
rect 17267 6273 17276 6307
rect 17224 6264 17276 6273
rect 19340 6264 19392 6316
rect 19432 6264 19484 6316
rect 22100 6264 22152 6316
rect 27160 6307 27212 6316
rect 27160 6273 27169 6307
rect 27169 6273 27203 6307
rect 27203 6273 27212 6307
rect 27160 6264 27212 6273
rect 27252 6264 27304 6316
rect 30196 6307 30248 6316
rect 22836 6196 22888 6248
rect 23664 6239 23716 6248
rect 23664 6205 23673 6239
rect 23673 6205 23707 6239
rect 23707 6205 23716 6239
rect 23664 6196 23716 6205
rect 23756 6196 23808 6248
rect 24952 6196 25004 6248
rect 26516 6196 26568 6248
rect 30196 6273 30205 6307
rect 30205 6273 30239 6307
rect 30239 6273 30248 6307
rect 30196 6264 30248 6273
rect 35808 6264 35860 6316
rect 34612 6196 34664 6248
rect 9588 6060 9640 6112
rect 13176 6060 13228 6112
rect 13636 6060 13688 6112
rect 19708 6128 19760 6180
rect 21640 6128 21692 6180
rect 22284 6128 22336 6180
rect 23848 6128 23900 6180
rect 25320 6128 25372 6180
rect 19340 6060 19392 6112
rect 21916 6060 21968 6112
rect 23020 6060 23072 6112
rect 23204 6060 23256 6112
rect 25964 6060 26016 6112
rect 26332 6060 26384 6112
rect 28264 6060 28316 6112
rect 33416 6060 33468 6112
rect 38016 6060 38068 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 2228 5856 2280 5908
rect 6000 5856 6052 5908
rect 6276 5899 6328 5908
rect 6276 5865 6285 5899
rect 6285 5865 6319 5899
rect 6319 5865 6328 5899
rect 6276 5856 6328 5865
rect 3240 5788 3292 5840
rect 7748 5856 7800 5908
rect 8116 5856 8168 5908
rect 8484 5831 8536 5840
rect 2228 5652 2280 5704
rect 2412 5652 2464 5704
rect 3332 5652 3384 5704
rect 4528 5695 4580 5704
rect 4528 5661 4537 5695
rect 4537 5661 4571 5695
rect 4571 5661 4580 5695
rect 4528 5652 4580 5661
rect 5264 5584 5316 5636
rect 8484 5797 8493 5831
rect 8493 5797 8527 5831
rect 8527 5797 8536 5831
rect 8484 5788 8536 5797
rect 11336 5788 11388 5840
rect 11980 5788 12032 5840
rect 14372 5856 14424 5908
rect 22284 5856 22336 5908
rect 22468 5856 22520 5908
rect 26332 5856 26384 5908
rect 26608 5856 26660 5908
rect 27528 5899 27580 5908
rect 27528 5865 27537 5899
rect 27537 5865 27571 5899
rect 27571 5865 27580 5899
rect 27528 5856 27580 5865
rect 6552 5720 6604 5772
rect 6736 5763 6788 5772
rect 6736 5729 6745 5763
rect 6745 5729 6779 5763
rect 6779 5729 6788 5763
rect 6736 5720 6788 5729
rect 7012 5720 7064 5772
rect 8300 5720 8352 5772
rect 9312 5763 9364 5772
rect 9312 5729 9321 5763
rect 9321 5729 9355 5763
rect 9355 5729 9364 5763
rect 9312 5720 9364 5729
rect 13728 5763 13780 5772
rect 13728 5729 13737 5763
rect 13737 5729 13771 5763
rect 13771 5729 13780 5763
rect 13728 5720 13780 5729
rect 14188 5720 14240 5772
rect 16212 5720 16264 5772
rect 17132 5763 17184 5772
rect 17132 5729 17141 5763
rect 17141 5729 17175 5763
rect 17175 5729 17184 5763
rect 17132 5720 17184 5729
rect 18972 5720 19024 5772
rect 19432 5720 19484 5772
rect 31852 5788 31904 5840
rect 21916 5720 21968 5772
rect 23020 5763 23072 5772
rect 23020 5729 23029 5763
rect 23029 5729 23063 5763
rect 23063 5729 23072 5763
rect 23020 5720 23072 5729
rect 23664 5720 23716 5772
rect 28724 5720 28776 5772
rect 28816 5720 28868 5772
rect 11796 5652 11848 5704
rect 21456 5652 21508 5704
rect 22192 5652 22244 5704
rect 25596 5652 25648 5704
rect 26240 5695 26292 5704
rect 26240 5661 26249 5695
rect 26249 5661 26283 5695
rect 26283 5661 26292 5695
rect 26240 5652 26292 5661
rect 26424 5652 26476 5704
rect 27160 5652 27212 5704
rect 27436 5695 27488 5704
rect 27436 5661 27445 5695
rect 27445 5661 27479 5695
rect 27479 5661 27488 5695
rect 27436 5652 27488 5661
rect 27988 5652 28040 5704
rect 29736 5695 29788 5704
rect 29736 5661 29745 5695
rect 29745 5661 29779 5695
rect 29779 5661 29788 5695
rect 29736 5652 29788 5661
rect 6644 5584 6696 5636
rect 7196 5516 7248 5568
rect 9036 5516 9088 5568
rect 12716 5584 12768 5636
rect 11152 5516 11204 5568
rect 14372 5516 14424 5568
rect 15108 5584 15160 5636
rect 17408 5627 17460 5636
rect 17408 5593 17417 5627
rect 17417 5593 17451 5627
rect 17451 5593 17460 5627
rect 17408 5584 17460 5593
rect 15936 5516 15988 5568
rect 18052 5516 18104 5568
rect 18972 5516 19024 5568
rect 20352 5584 20404 5636
rect 23020 5584 23072 5636
rect 23112 5627 23164 5636
rect 23112 5593 23121 5627
rect 23121 5593 23155 5627
rect 23155 5593 23164 5627
rect 23112 5584 23164 5593
rect 24308 5584 24360 5636
rect 25688 5627 25740 5636
rect 21548 5559 21600 5568
rect 21548 5525 21557 5559
rect 21557 5525 21591 5559
rect 21591 5525 21600 5559
rect 21548 5516 21600 5525
rect 22468 5516 22520 5568
rect 24400 5516 24452 5568
rect 25688 5593 25697 5627
rect 25697 5593 25731 5627
rect 25731 5593 25740 5627
rect 25688 5584 25740 5593
rect 26240 5516 26292 5568
rect 27988 5516 28040 5568
rect 28172 5559 28224 5568
rect 28172 5525 28181 5559
rect 28181 5525 28215 5559
rect 28215 5525 28224 5559
rect 28172 5516 28224 5525
rect 28724 5559 28776 5568
rect 28724 5525 28733 5559
rect 28733 5525 28767 5559
rect 28767 5525 28776 5559
rect 28724 5516 28776 5525
rect 29828 5559 29880 5568
rect 29828 5525 29837 5559
rect 29837 5525 29871 5559
rect 29871 5525 29880 5559
rect 29828 5516 29880 5525
rect 38200 5559 38252 5568
rect 38200 5525 38209 5559
rect 38209 5525 38243 5559
rect 38243 5525 38252 5559
rect 38200 5516 38252 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 2136 5312 2188 5364
rect 2964 5312 3016 5364
rect 2228 5244 2280 5296
rect 2320 5219 2372 5228
rect 2320 5185 2329 5219
rect 2329 5185 2363 5219
rect 2363 5185 2372 5219
rect 2320 5176 2372 5185
rect 3332 5176 3384 5228
rect 3608 5219 3660 5228
rect 3608 5185 3617 5219
rect 3617 5185 3651 5219
rect 3651 5185 3660 5219
rect 3608 5176 3660 5185
rect 4620 5244 4672 5296
rect 6092 5244 6144 5296
rect 6000 5176 6052 5228
rect 7196 5244 7248 5296
rect 7472 5287 7524 5296
rect 7472 5253 7481 5287
rect 7481 5253 7515 5287
rect 7515 5253 7524 5287
rect 7472 5244 7524 5253
rect 7564 5244 7616 5296
rect 4528 5151 4580 5160
rect 4528 5117 4537 5151
rect 4537 5117 4571 5151
rect 4571 5117 4580 5151
rect 7196 5151 7248 5160
rect 4528 5108 4580 5117
rect 7196 5117 7205 5151
rect 7205 5117 7239 5151
rect 7239 5117 7248 5151
rect 7196 5108 7248 5117
rect 14556 5312 14608 5364
rect 14648 5312 14700 5364
rect 15936 5355 15988 5364
rect 9956 5244 10008 5296
rect 13452 5244 13504 5296
rect 13820 5244 13872 5296
rect 15936 5321 15945 5355
rect 15945 5321 15979 5355
rect 15979 5321 15988 5355
rect 15936 5312 15988 5321
rect 16120 5312 16172 5364
rect 20076 5312 20128 5364
rect 21916 5312 21968 5364
rect 21640 5244 21692 5296
rect 21732 5244 21784 5296
rect 9312 5176 9364 5228
rect 13544 5176 13596 5228
rect 10048 5108 10100 5160
rect 11152 5151 11204 5160
rect 11152 5117 11161 5151
rect 11161 5117 11195 5151
rect 11195 5117 11204 5151
rect 11152 5108 11204 5117
rect 11704 5151 11756 5160
rect 11704 5117 11713 5151
rect 11713 5117 11747 5151
rect 11747 5117 11756 5151
rect 11704 5108 11756 5117
rect 14188 5151 14240 5160
rect 2872 4972 2924 5024
rect 5540 5040 5592 5092
rect 6828 5040 6880 5092
rect 5908 4972 5960 5024
rect 9128 4972 9180 5024
rect 13820 4972 13872 5024
rect 14188 5117 14197 5151
rect 14197 5117 14231 5151
rect 14231 5117 14240 5151
rect 14188 5108 14240 5117
rect 14464 5151 14516 5160
rect 14464 5117 14473 5151
rect 14473 5117 14507 5151
rect 14507 5117 14516 5151
rect 14464 5108 14516 5117
rect 14556 5108 14608 5160
rect 15660 5108 15712 5160
rect 16120 5108 16172 5160
rect 16948 5151 17000 5160
rect 16948 5117 16957 5151
rect 16957 5117 16991 5151
rect 16991 5117 17000 5151
rect 16948 5108 17000 5117
rect 18880 5176 18932 5228
rect 19432 5176 19484 5228
rect 22560 5244 22612 5296
rect 24584 5176 24636 5228
rect 28172 5244 28224 5296
rect 28632 5244 28684 5296
rect 19340 5108 19392 5160
rect 21272 5108 21324 5160
rect 22928 5108 22980 5160
rect 23204 5151 23256 5160
rect 23204 5117 23213 5151
rect 23213 5117 23247 5151
rect 23247 5117 23256 5151
rect 23204 5108 23256 5117
rect 24032 5151 24084 5160
rect 24032 5117 24041 5151
rect 24041 5117 24075 5151
rect 24075 5117 24084 5151
rect 24032 5108 24084 5117
rect 16304 4972 16356 5024
rect 19524 5040 19576 5092
rect 18788 4972 18840 5024
rect 21916 5040 21968 5092
rect 22008 5040 22060 5092
rect 26792 5176 26844 5228
rect 25688 5108 25740 5160
rect 28356 5176 28408 5228
rect 29000 5176 29052 5228
rect 29184 5176 29236 5228
rect 30380 5219 30432 5228
rect 30380 5185 30389 5219
rect 30389 5185 30423 5219
rect 30423 5185 30432 5219
rect 30380 5176 30432 5185
rect 32956 5108 33008 5160
rect 28264 5040 28316 5092
rect 30012 5040 30064 5092
rect 20904 4972 20956 5024
rect 22376 4972 22428 5024
rect 23296 4972 23348 5024
rect 23388 4972 23440 5024
rect 26792 4972 26844 5024
rect 27528 4972 27580 5024
rect 29276 4972 29328 5024
rect 30564 4972 30616 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 1584 4607 1636 4616
rect 1584 4573 1593 4607
rect 1593 4573 1627 4607
rect 1627 4573 1636 4607
rect 1584 4564 1636 4573
rect 3792 4700 3844 4752
rect 7564 4768 7616 4820
rect 8300 4768 8352 4820
rect 9956 4768 10008 4820
rect 10508 4768 10560 4820
rect 18788 4768 18840 4820
rect 5908 4700 5960 4752
rect 4896 4632 4948 4684
rect 6736 4675 6788 4684
rect 6736 4641 6745 4675
rect 6745 4641 6779 4675
rect 6779 4641 6788 4675
rect 6736 4632 6788 4641
rect 8208 4700 8260 4752
rect 9496 4700 9548 4752
rect 7380 4632 7432 4684
rect 9588 4675 9640 4684
rect 9588 4641 9597 4675
rect 9597 4641 9631 4675
rect 9631 4641 9640 4675
rect 9588 4632 9640 4641
rect 11152 4632 11204 4684
rect 11796 4675 11848 4684
rect 11796 4641 11805 4675
rect 11805 4641 11839 4675
rect 11839 4641 11848 4675
rect 11796 4632 11848 4641
rect 14464 4700 14516 4752
rect 16304 4743 16356 4752
rect 16304 4709 16313 4743
rect 16313 4709 16347 4743
rect 16347 4709 16356 4743
rect 16304 4700 16356 4709
rect 21272 4743 21324 4752
rect 21272 4709 21281 4743
rect 21281 4709 21315 4743
rect 21315 4709 21324 4743
rect 21272 4700 21324 4709
rect 13268 4632 13320 4684
rect 17316 4632 17368 4684
rect 19248 4632 19300 4684
rect 22008 4768 22060 4820
rect 25688 4700 25740 4752
rect 26700 4700 26752 4752
rect 26884 4700 26936 4752
rect 3240 4607 3292 4616
rect 3240 4573 3249 4607
rect 3249 4573 3283 4607
rect 3283 4573 3292 4607
rect 3240 4564 3292 4573
rect 4528 4607 4580 4616
rect 4528 4573 4537 4607
rect 4537 4573 4571 4607
rect 4571 4573 4580 4607
rect 4528 4564 4580 4573
rect 14280 4564 14332 4616
rect 16948 4564 17000 4616
rect 19156 4564 19208 4616
rect 24124 4632 24176 4684
rect 24952 4675 25004 4684
rect 24952 4641 24961 4675
rect 24961 4641 24995 4675
rect 24995 4641 25004 4675
rect 24952 4632 25004 4641
rect 25780 4675 25832 4684
rect 25780 4641 25789 4675
rect 25789 4641 25823 4675
rect 25823 4641 25832 4675
rect 25780 4632 25832 4641
rect 26240 4632 26292 4684
rect 26792 4632 26844 4684
rect 28816 4743 28868 4752
rect 28816 4709 28825 4743
rect 28825 4709 28859 4743
rect 28859 4709 28868 4743
rect 28816 4700 28868 4709
rect 27804 4632 27856 4684
rect 29276 4632 29328 4684
rect 21732 4607 21784 4616
rect 21732 4573 21741 4607
rect 21741 4573 21775 4607
rect 21775 4573 21784 4607
rect 21732 4564 21784 4573
rect 26424 4564 26476 4616
rect 28172 4564 28224 4616
rect 28356 4564 28408 4616
rect 30012 4768 30064 4820
rect 31760 4811 31812 4820
rect 31760 4777 31769 4811
rect 31769 4777 31803 4811
rect 31803 4777 31812 4811
rect 31760 4768 31812 4777
rect 37832 4768 37884 4820
rect 5816 4496 5868 4548
rect 1768 4471 1820 4480
rect 1768 4437 1777 4471
rect 1777 4437 1811 4471
rect 1811 4437 1820 4471
rect 1768 4428 1820 4437
rect 6920 4496 6972 4548
rect 8392 4428 8444 4480
rect 11796 4496 11848 4548
rect 12072 4539 12124 4548
rect 12072 4505 12081 4539
rect 12081 4505 12115 4539
rect 12115 4505 12124 4539
rect 12072 4496 12124 4505
rect 10048 4428 10100 4480
rect 12256 4428 12308 4480
rect 13544 4471 13596 4480
rect 13544 4437 13553 4471
rect 13553 4437 13587 4471
rect 13587 4437 13596 4471
rect 13544 4428 13596 4437
rect 14832 4539 14884 4548
rect 14832 4505 14841 4539
rect 14841 4505 14875 4539
rect 14875 4505 14884 4539
rect 14832 4496 14884 4505
rect 15108 4496 15160 4548
rect 17224 4496 17276 4548
rect 16580 4428 16632 4480
rect 18696 4428 18748 4480
rect 18880 4428 18932 4480
rect 19984 4428 20036 4480
rect 21180 4496 21232 4548
rect 21548 4496 21600 4548
rect 24768 4496 24820 4548
rect 25504 4496 25556 4548
rect 27804 4496 27856 4548
rect 28264 4496 28316 4548
rect 30380 4607 30432 4616
rect 30380 4573 30389 4607
rect 30389 4573 30423 4607
rect 30423 4573 30432 4607
rect 30380 4564 30432 4573
rect 31668 4607 31720 4616
rect 31668 4573 31677 4607
rect 31677 4573 31711 4607
rect 31711 4573 31720 4607
rect 31668 4564 31720 4573
rect 34704 4564 34756 4616
rect 33048 4496 33100 4548
rect 38108 4539 38160 4548
rect 38108 4505 38117 4539
rect 38117 4505 38151 4539
rect 38151 4505 38160 4539
rect 38108 4496 38160 4505
rect 20720 4428 20772 4480
rect 20812 4428 20864 4480
rect 21916 4428 21968 4480
rect 22284 4428 22336 4480
rect 26240 4428 26292 4480
rect 28908 4428 28960 4480
rect 31024 4471 31076 4480
rect 31024 4437 31033 4471
rect 31033 4437 31067 4471
rect 31067 4437 31076 4471
rect 31024 4428 31076 4437
rect 33508 4428 33560 4480
rect 33600 4471 33652 4480
rect 33600 4437 33609 4471
rect 33609 4437 33643 4471
rect 33643 4437 33652 4471
rect 33600 4428 33652 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 4068 4224 4120 4276
rect 8024 4224 8076 4276
rect 8116 4224 8168 4276
rect 12256 4224 12308 4276
rect 3240 4156 3292 4208
rect 3700 4156 3752 4208
rect 3516 4088 3568 4140
rect 4160 4131 4212 4140
rect 4160 4097 4169 4131
rect 4169 4097 4203 4131
rect 4203 4097 4212 4131
rect 4160 4088 4212 4097
rect 3240 4020 3292 4072
rect 4712 4088 4764 4140
rect 5816 4156 5868 4208
rect 6460 4156 6512 4208
rect 7932 4156 7984 4208
rect 7104 4131 7156 4140
rect 7104 4097 7113 4131
rect 7113 4097 7147 4131
rect 7147 4097 7156 4131
rect 7104 4088 7156 4097
rect 7012 4020 7064 4072
rect 7932 4020 7984 4072
rect 8024 4020 8076 4072
rect 9128 4131 9180 4140
rect 9128 4097 9137 4131
rect 9137 4097 9171 4131
rect 9171 4097 9180 4131
rect 9128 4088 9180 4097
rect 10140 4156 10192 4208
rect 12624 4224 12676 4276
rect 13268 4224 13320 4276
rect 12532 4156 12584 4208
rect 17316 4224 17368 4276
rect 22744 4224 22796 4276
rect 11704 4088 11756 4140
rect 2964 3884 3016 3936
rect 3792 3884 3844 3936
rect 5080 3884 5132 3936
rect 5172 3884 5224 3936
rect 8392 3952 8444 4004
rect 9220 3952 9272 4004
rect 9680 3952 9732 4004
rect 10048 4020 10100 4072
rect 11060 4020 11112 4072
rect 12624 4020 12676 4072
rect 17224 4156 17276 4208
rect 18880 4156 18932 4208
rect 24768 4224 24820 4276
rect 25780 4224 25832 4276
rect 26884 4224 26936 4276
rect 26976 4224 27028 4276
rect 23296 4199 23348 4208
rect 23296 4165 23305 4199
rect 23305 4165 23339 4199
rect 23339 4165 23348 4199
rect 23296 4156 23348 4165
rect 25044 4156 25096 4208
rect 27528 4156 27580 4208
rect 27988 4156 28040 4208
rect 29000 4224 29052 4276
rect 30656 4224 30708 4276
rect 33600 4156 33652 4208
rect 14280 4020 14332 4072
rect 18052 4088 18104 4140
rect 20536 4088 20588 4140
rect 20720 4131 20772 4140
rect 20720 4097 20729 4131
rect 20729 4097 20763 4131
rect 20763 4097 20772 4131
rect 20720 4088 20772 4097
rect 21088 4088 21140 4140
rect 21364 4131 21416 4140
rect 21364 4097 21373 4131
rect 21373 4097 21407 4131
rect 21407 4097 21416 4131
rect 21364 4088 21416 4097
rect 21916 4088 21968 4140
rect 22560 4131 22612 4140
rect 22560 4097 22569 4131
rect 22569 4097 22603 4131
rect 22603 4097 22612 4131
rect 27160 4131 27212 4140
rect 22560 4088 22612 4097
rect 27160 4097 27169 4131
rect 27169 4097 27203 4131
rect 27203 4097 27212 4131
rect 27160 4088 27212 4097
rect 27896 4088 27948 4140
rect 28172 4088 28224 4140
rect 28356 4088 28408 4140
rect 29000 4088 29052 4140
rect 29736 4131 29788 4140
rect 29736 4097 29745 4131
rect 29745 4097 29779 4131
rect 29779 4097 29788 4131
rect 29736 4088 29788 4097
rect 30012 4088 30064 4140
rect 30472 4131 30524 4140
rect 30472 4097 30481 4131
rect 30481 4097 30515 4131
rect 30515 4097 30524 4131
rect 30472 4088 30524 4097
rect 30656 4088 30708 4140
rect 31576 4088 31628 4140
rect 32496 4131 32548 4140
rect 32496 4097 32505 4131
rect 32505 4097 32539 4131
rect 32539 4097 32548 4131
rect 32496 4088 32548 4097
rect 33508 4088 33560 4140
rect 16580 4020 16632 4072
rect 16948 4020 17000 4072
rect 11336 3952 11388 4004
rect 13360 3884 13412 3936
rect 13452 3884 13504 3936
rect 14556 3884 14608 3936
rect 16764 3884 16816 3936
rect 18236 3952 18288 4004
rect 18696 4020 18748 4072
rect 20812 4020 20864 4072
rect 23204 4063 23256 4072
rect 23204 4029 23213 4063
rect 23213 4029 23247 4063
rect 23247 4029 23256 4063
rect 23204 4020 23256 4029
rect 24124 4063 24176 4072
rect 24124 4029 24133 4063
rect 24133 4029 24167 4063
rect 24167 4029 24176 4063
rect 24124 4020 24176 4029
rect 24400 4020 24452 4072
rect 24860 4020 24912 4072
rect 26056 4020 26108 4072
rect 27620 4020 27672 4072
rect 21088 3952 21140 4004
rect 23756 3952 23808 4004
rect 25596 3952 25648 4004
rect 26424 3952 26476 4004
rect 19156 3884 19208 3936
rect 19984 3884 20036 3936
rect 22652 3884 22704 3936
rect 25320 3884 25372 3936
rect 25964 3884 26016 3936
rect 30932 3952 30984 4004
rect 33784 3952 33836 4004
rect 26792 3884 26844 3936
rect 27988 3884 28040 3936
rect 30012 3884 30064 3936
rect 30288 3884 30340 3936
rect 32312 3927 32364 3936
rect 32312 3893 32321 3927
rect 32321 3893 32355 3927
rect 32355 3893 32364 3927
rect 32312 3884 32364 3893
rect 34796 3884 34848 3936
rect 37188 3884 37240 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 4068 3723 4120 3732
rect 4068 3689 4077 3723
rect 4077 3689 4111 3723
rect 4111 3689 4120 3723
rect 4068 3680 4120 3689
rect 4528 3680 4580 3732
rect 6920 3680 6972 3732
rect 2228 3587 2280 3596
rect 2228 3553 2237 3587
rect 2237 3553 2271 3587
rect 2271 3553 2280 3587
rect 2228 3544 2280 3553
rect 4528 3544 4580 3596
rect 4620 3587 4672 3596
rect 4620 3553 4629 3587
rect 4629 3553 4663 3587
rect 4663 3553 4672 3587
rect 4620 3544 4672 3553
rect 6552 3612 6604 3664
rect 8208 3612 8260 3664
rect 9496 3680 9548 3732
rect 6736 3544 6788 3596
rect 7196 3544 7248 3596
rect 9128 3612 9180 3664
rect 9956 3612 10008 3664
rect 10692 3680 10744 3732
rect 11888 3680 11940 3732
rect 12900 3680 12952 3732
rect 16028 3723 16080 3732
rect 14188 3612 14240 3664
rect 16028 3689 16037 3723
rect 16037 3689 16071 3723
rect 16071 3689 16080 3723
rect 16028 3680 16080 3689
rect 22192 3680 22244 3732
rect 23848 3723 23900 3732
rect 12532 3544 12584 3596
rect 2596 3519 2648 3528
rect 2596 3485 2605 3519
rect 2605 3485 2639 3519
rect 2639 3485 2648 3519
rect 2596 3476 2648 3485
rect 3700 3476 3752 3528
rect 3976 3519 4028 3528
rect 3976 3485 3985 3519
rect 3985 3485 4019 3519
rect 4019 3485 4028 3519
rect 3976 3476 4028 3485
rect 9588 3476 9640 3528
rect 10048 3519 10100 3528
rect 10048 3485 10057 3519
rect 10057 3485 10091 3519
rect 10091 3485 10100 3519
rect 10048 3476 10100 3485
rect 13268 3544 13320 3596
rect 16948 3544 17000 3596
rect 18420 3544 18472 3596
rect 19156 3544 19208 3596
rect 20904 3612 20956 3664
rect 23848 3689 23857 3723
rect 23857 3689 23891 3723
rect 23891 3689 23900 3723
rect 23848 3680 23900 3689
rect 24492 3680 24544 3732
rect 26700 3612 26752 3664
rect 22652 3587 22704 3596
rect 14280 3519 14332 3528
rect 14280 3485 14289 3519
rect 14289 3485 14323 3519
rect 14323 3485 14332 3519
rect 14280 3476 14332 3485
rect 4804 3408 4856 3460
rect 4988 3408 5040 3460
rect 5632 3408 5684 3460
rect 1768 3383 1820 3392
rect 1768 3349 1777 3383
rect 1777 3349 1811 3383
rect 1811 3349 1820 3383
rect 1768 3340 1820 3349
rect 2964 3340 3016 3392
rect 8760 3408 8812 3460
rect 9404 3451 9456 3460
rect 9404 3417 9413 3451
rect 9413 3417 9447 3451
rect 9447 3417 9456 3451
rect 9404 3408 9456 3417
rect 9864 3408 9916 3460
rect 12624 3408 12676 3460
rect 13176 3408 13228 3460
rect 13912 3408 13964 3460
rect 14464 3408 14516 3460
rect 6920 3340 6972 3392
rect 12348 3340 12400 3392
rect 13360 3340 13412 3392
rect 18512 3476 18564 3528
rect 22652 3553 22661 3587
rect 22661 3553 22695 3587
rect 22695 3553 22704 3587
rect 22652 3544 22704 3553
rect 22744 3544 22796 3596
rect 26792 3544 26844 3596
rect 27068 3587 27120 3596
rect 27068 3553 27077 3587
rect 27077 3553 27111 3587
rect 27111 3553 27120 3587
rect 27068 3544 27120 3553
rect 27528 3680 27580 3732
rect 29276 3680 29328 3732
rect 29460 3680 29512 3732
rect 30748 3680 30800 3732
rect 32956 3723 33008 3732
rect 27252 3612 27304 3664
rect 29828 3612 29880 3664
rect 32956 3689 32965 3723
rect 32965 3689 32999 3723
rect 32999 3689 33008 3723
rect 32956 3680 33008 3689
rect 21916 3519 21968 3528
rect 21916 3485 21925 3519
rect 21925 3485 21959 3519
rect 21959 3485 21968 3519
rect 21916 3476 21968 3485
rect 22284 3476 22336 3528
rect 23296 3519 23348 3528
rect 23296 3485 23305 3519
rect 23305 3485 23339 3519
rect 23339 3485 23348 3519
rect 23756 3519 23808 3528
rect 23296 3476 23348 3485
rect 23756 3485 23765 3519
rect 23765 3485 23799 3519
rect 23799 3485 23808 3519
rect 23756 3476 23808 3485
rect 25320 3519 25372 3528
rect 25320 3485 25329 3519
rect 25329 3485 25363 3519
rect 25363 3485 25372 3519
rect 25320 3476 25372 3485
rect 17408 3451 17460 3460
rect 17408 3417 17417 3451
rect 17417 3417 17451 3451
rect 17451 3417 17460 3451
rect 17408 3408 17460 3417
rect 21456 3451 21508 3460
rect 21456 3417 21465 3451
rect 21465 3417 21499 3451
rect 21499 3417 21508 3451
rect 21456 3408 21508 3417
rect 22744 3451 22796 3460
rect 22744 3417 22753 3451
rect 22753 3417 22787 3451
rect 22787 3417 22796 3451
rect 22744 3408 22796 3417
rect 24676 3451 24728 3460
rect 24676 3417 24685 3451
rect 24685 3417 24719 3451
rect 24719 3417 24728 3451
rect 24676 3408 24728 3417
rect 25872 3451 25924 3460
rect 18788 3340 18840 3392
rect 19340 3340 19392 3392
rect 25872 3417 25881 3451
rect 25881 3417 25915 3451
rect 25915 3417 25924 3451
rect 25872 3408 25924 3417
rect 25964 3451 26016 3460
rect 25964 3417 25973 3451
rect 25973 3417 26007 3451
rect 26007 3417 26016 3451
rect 25964 3408 26016 3417
rect 26240 3408 26292 3460
rect 27068 3408 27120 3460
rect 27344 3408 27396 3460
rect 28080 3451 28132 3460
rect 28080 3417 28089 3451
rect 28089 3417 28123 3451
rect 28123 3417 28132 3451
rect 28080 3408 28132 3417
rect 28448 3544 28500 3596
rect 28356 3476 28408 3528
rect 28816 3476 28868 3528
rect 29000 3476 29052 3528
rect 32312 3544 32364 3596
rect 30748 3476 30800 3528
rect 31300 3476 31352 3528
rect 31944 3476 31996 3528
rect 33784 3519 33836 3528
rect 33784 3485 33793 3519
rect 33793 3485 33827 3519
rect 33827 3485 33836 3519
rect 33784 3476 33836 3485
rect 38016 3519 38068 3528
rect 38016 3485 38025 3519
rect 38025 3485 38059 3519
rect 38059 3485 38068 3519
rect 38016 3476 38068 3485
rect 24860 3340 24912 3392
rect 27988 3340 28040 3392
rect 28540 3340 28592 3392
rect 28816 3340 28868 3392
rect 29460 3340 29512 3392
rect 29644 3340 29696 3392
rect 30472 3383 30524 3392
rect 30472 3349 30481 3383
rect 30481 3349 30515 3383
rect 30515 3349 30524 3383
rect 30472 3340 30524 3349
rect 31116 3383 31168 3392
rect 31116 3349 31125 3383
rect 31125 3349 31159 3383
rect 31159 3349 31168 3383
rect 31116 3340 31168 3349
rect 31484 3340 31536 3392
rect 31760 3340 31812 3392
rect 38200 3383 38252 3392
rect 38200 3349 38209 3383
rect 38209 3349 38243 3383
rect 38243 3349 38252 3383
rect 38200 3340 38252 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 2780 3136 2832 3188
rect 3148 3136 3200 3188
rect 3792 3136 3844 3188
rect 5540 3136 5592 3188
rect 6368 3136 6420 3188
rect 2412 3111 2464 3120
rect 2412 3077 2421 3111
rect 2421 3077 2455 3111
rect 2455 3077 2464 3111
rect 2412 3068 2464 3077
rect 2872 3000 2924 3052
rect 3240 3000 3292 3052
rect 3792 3043 3844 3052
rect 3792 3009 3801 3043
rect 3801 3009 3835 3043
rect 3835 3009 3844 3043
rect 3792 3000 3844 3009
rect 4620 3068 4672 3120
rect 4804 3068 4856 3120
rect 11888 3136 11940 3188
rect 8116 3111 8168 3120
rect 8116 3077 8125 3111
rect 8125 3077 8159 3111
rect 8159 3077 8168 3111
rect 8116 3068 8168 3077
rect 8576 3068 8628 3120
rect 11152 3068 11204 3120
rect 23204 3136 23256 3188
rect 24032 3136 24084 3188
rect 7196 3000 7248 3052
rect 7748 3000 7800 3052
rect 4528 2975 4580 2984
rect 4528 2941 4537 2975
rect 4537 2941 4571 2975
rect 4571 2941 4580 2975
rect 4528 2932 4580 2941
rect 5080 2932 5132 2984
rect 10232 3000 10284 3052
rect 10508 3000 10560 3052
rect 10876 3000 10928 3052
rect 12900 3043 12952 3052
rect 664 2796 716 2848
rect 6460 2796 6512 2848
rect 7104 2796 7156 2848
rect 7656 2796 7708 2848
rect 9128 2864 9180 2916
rect 10600 2932 10652 2984
rect 11152 2932 11204 2984
rect 11980 2907 12032 2916
rect 11980 2873 11989 2907
rect 11989 2873 12023 2907
rect 12023 2873 12032 2907
rect 11980 2864 12032 2873
rect 12900 3009 12909 3043
rect 12909 3009 12943 3043
rect 12943 3009 12952 3043
rect 12900 3000 12952 3009
rect 13544 3068 13596 3120
rect 15016 3068 15068 3120
rect 16304 3111 16356 3120
rect 16304 3077 16313 3111
rect 16313 3077 16347 3111
rect 16347 3077 16356 3111
rect 16304 3068 16356 3077
rect 19064 3068 19116 3120
rect 19156 3068 19208 3120
rect 26240 3136 26292 3188
rect 27436 3136 27488 3188
rect 33048 3179 33100 3188
rect 33048 3145 33057 3179
rect 33057 3145 33091 3179
rect 33091 3145 33100 3179
rect 33048 3136 33100 3145
rect 34704 3136 34756 3188
rect 13268 3000 13320 3052
rect 16120 3043 16172 3052
rect 16120 3009 16129 3043
rect 16129 3009 16163 3043
rect 16163 3009 16172 3043
rect 16120 3000 16172 3009
rect 16948 3000 17000 3052
rect 18972 3000 19024 3052
rect 14832 2932 14884 2984
rect 14924 2932 14976 2984
rect 19156 2932 19208 2984
rect 19524 2975 19576 2984
rect 19524 2941 19533 2975
rect 19533 2941 19567 2975
rect 19567 2941 19576 2975
rect 19524 2932 19576 2941
rect 20536 2932 20588 2984
rect 21732 3000 21784 3052
rect 23388 3000 23440 3052
rect 20720 2932 20772 2984
rect 24860 2932 24912 2984
rect 25136 2975 25188 2984
rect 25136 2941 25145 2975
rect 25145 2941 25179 2975
rect 25179 2941 25188 2975
rect 25136 2932 25188 2941
rect 13360 2796 13412 2848
rect 14832 2796 14884 2848
rect 17408 2796 17460 2848
rect 20076 2796 20128 2848
rect 21824 2796 21876 2848
rect 24952 2864 25004 2916
rect 26976 3068 27028 3120
rect 27344 3111 27396 3120
rect 27344 3077 27346 3111
rect 27346 3077 27380 3111
rect 27380 3077 27396 3111
rect 27344 3068 27396 3077
rect 27620 3068 27672 3120
rect 28356 3043 28408 3052
rect 28356 3009 28365 3043
rect 28365 3009 28399 3043
rect 28399 3009 28408 3043
rect 28356 3000 28408 3009
rect 29092 3000 29144 3052
rect 26148 2932 26200 2984
rect 27252 2975 27304 2984
rect 27252 2941 27261 2975
rect 27261 2941 27295 2975
rect 27295 2941 27304 2975
rect 27252 2932 27304 2941
rect 27344 2932 27396 2984
rect 26424 2907 26476 2916
rect 26424 2873 26433 2907
rect 26433 2873 26467 2907
rect 26467 2873 26476 2907
rect 26424 2864 26476 2873
rect 26976 2864 27028 2916
rect 28908 2932 28960 2984
rect 30380 3068 30432 3120
rect 29552 3000 29604 3052
rect 29920 3000 29972 3052
rect 31576 3043 31628 3052
rect 31576 3009 31585 3043
rect 31585 3009 31619 3043
rect 31619 3009 31628 3043
rect 31576 3000 31628 3009
rect 31852 3000 31904 3052
rect 32404 3000 32456 3052
rect 30656 2932 30708 2984
rect 31944 2864 31996 2916
rect 35440 3000 35492 3052
rect 37832 3000 37884 3052
rect 37924 3000 37976 3052
rect 34612 2864 34664 2916
rect 28448 2839 28500 2848
rect 28448 2805 28457 2839
rect 28457 2805 28491 2839
rect 28491 2805 28500 2839
rect 28448 2796 28500 2805
rect 29736 2839 29788 2848
rect 29736 2805 29745 2839
rect 29745 2805 29779 2839
rect 29779 2805 29788 2839
rect 29736 2796 29788 2805
rect 30380 2839 30432 2848
rect 30380 2805 30389 2839
rect 30389 2805 30423 2839
rect 30423 2805 30432 2839
rect 30380 2796 30432 2805
rect 30472 2796 30524 2848
rect 31668 2839 31720 2848
rect 31668 2805 31677 2839
rect 31677 2805 31711 2839
rect 31711 2805 31720 2839
rect 31668 2796 31720 2805
rect 38660 2796 38712 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 4988 2592 5040 2644
rect 7472 2592 7524 2644
rect 20 2524 72 2576
rect 4620 2456 4672 2508
rect 7012 2456 7064 2508
rect 7748 2456 7800 2508
rect 16304 2567 16356 2576
rect 16304 2533 16313 2567
rect 16313 2533 16347 2567
rect 16347 2533 16356 2567
rect 16304 2524 16356 2533
rect 13268 2456 13320 2508
rect 13912 2456 13964 2508
rect 15476 2456 15528 2508
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 2504 2388 2556 2440
rect 3148 2431 3200 2440
rect 3148 2397 3157 2431
rect 3157 2397 3191 2431
rect 3191 2397 3200 2431
rect 3148 2388 3200 2397
rect 4528 2363 4580 2372
rect 4528 2329 4537 2363
rect 4537 2329 4571 2363
rect 4571 2329 4580 2363
rect 4528 2320 4580 2329
rect 5816 2320 5868 2372
rect 6368 2320 6420 2372
rect 7472 2320 7524 2372
rect 12256 2363 12308 2372
rect 1952 2252 2004 2304
rect 3240 2252 3292 2304
rect 5540 2252 5592 2304
rect 8484 2295 8536 2304
rect 8484 2261 8493 2295
rect 8493 2261 8527 2295
rect 8527 2261 8536 2295
rect 8484 2252 8536 2261
rect 9772 2252 9824 2304
rect 11152 2295 11204 2304
rect 11152 2261 11161 2295
rect 11161 2261 11195 2295
rect 11195 2261 11204 2295
rect 11152 2252 11204 2261
rect 12256 2329 12265 2363
rect 12265 2329 12299 2363
rect 12299 2329 12308 2363
rect 12256 2320 12308 2329
rect 15292 2320 15344 2372
rect 13636 2252 13688 2304
rect 16212 2252 16264 2304
rect 20444 2592 20496 2644
rect 18972 2524 19024 2576
rect 16948 2456 17000 2508
rect 19248 2456 19300 2508
rect 22928 2592 22980 2644
rect 22376 2524 22428 2576
rect 26608 2592 26660 2644
rect 26700 2592 26752 2644
rect 28356 2592 28408 2644
rect 23940 2456 23992 2508
rect 25136 2456 25188 2508
rect 21272 2388 21324 2440
rect 24860 2431 24912 2440
rect 19432 2320 19484 2372
rect 19708 2363 19760 2372
rect 19708 2329 19717 2363
rect 19717 2329 19751 2363
rect 19751 2329 19760 2363
rect 19708 2320 19760 2329
rect 23112 2363 23164 2372
rect 23112 2329 23121 2363
rect 23121 2329 23155 2363
rect 23155 2329 23164 2363
rect 23112 2320 23164 2329
rect 23204 2320 23256 2372
rect 24860 2397 24869 2431
rect 24869 2397 24903 2431
rect 24903 2397 24912 2431
rect 24860 2388 24912 2397
rect 30564 2524 30616 2576
rect 37096 2524 37148 2576
rect 25964 2499 26016 2508
rect 25964 2465 25973 2499
rect 25973 2465 26007 2499
rect 26007 2465 26016 2499
rect 25964 2456 26016 2465
rect 26424 2499 26476 2508
rect 26424 2465 26433 2499
rect 26433 2465 26467 2499
rect 26467 2465 26476 2499
rect 26424 2456 26476 2465
rect 26608 2456 26660 2508
rect 28448 2456 28500 2508
rect 32588 2499 32640 2508
rect 32588 2465 32597 2499
rect 32597 2465 32631 2499
rect 32631 2465 32640 2499
rect 32588 2456 32640 2465
rect 35348 2456 35400 2508
rect 37740 2499 37792 2508
rect 27160 2431 27212 2440
rect 27160 2397 27169 2431
rect 27169 2397 27203 2431
rect 27203 2397 27212 2431
rect 27160 2388 27212 2397
rect 27712 2388 27764 2440
rect 29368 2388 29420 2440
rect 31024 2388 31076 2440
rect 31300 2388 31352 2440
rect 32220 2388 32272 2440
rect 33416 2388 33468 2440
rect 34796 2388 34848 2440
rect 35532 2388 35584 2440
rect 37740 2465 37749 2499
rect 37749 2465 37783 2499
rect 37783 2465 37792 2499
rect 37740 2456 37792 2465
rect 37372 2388 37424 2440
rect 18696 2252 18748 2304
rect 19156 2252 19208 2304
rect 21180 2295 21232 2304
rect 21180 2261 21189 2295
rect 21189 2261 21223 2295
rect 21223 2261 21232 2295
rect 21180 2252 21232 2261
rect 22560 2252 22612 2304
rect 27712 2252 27764 2304
rect 29000 2252 29052 2304
rect 30288 2252 30340 2304
rect 31300 2295 31352 2304
rect 31300 2261 31309 2295
rect 31309 2261 31343 2295
rect 31343 2261 31352 2295
rect 31300 2252 31352 2261
rect 33508 2252 33560 2304
rect 34152 2252 34204 2304
rect 36728 2252 36780 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 3424 2048 3476 2100
rect 7472 2048 7524 2100
rect 3792 1980 3844 2032
rect 18052 2048 18104 2100
rect 18512 2048 18564 2100
rect 22744 2048 22796 2100
rect 22928 2048 22980 2100
rect 31116 2048 31168 2100
rect 4712 1844 4764 1896
rect 15292 1980 15344 2032
rect 19064 1980 19116 2032
rect 23020 1980 23072 2032
rect 23112 1980 23164 2032
rect 30380 1980 30432 2032
rect 11152 1912 11204 1964
rect 15476 1912 15528 1964
rect 15752 1912 15804 1964
rect 27160 1912 27212 1964
rect 16304 1844 16356 1896
rect 22836 1844 22888 1896
rect 24952 1844 25004 1896
rect 31300 1844 31352 1896
rect 4528 1776 4580 1828
rect 11060 1776 11112 1828
rect 13452 1776 13504 1828
rect 21180 1776 21232 1828
rect 27896 1776 27948 1828
rect 2320 1708 2372 1760
rect 8484 1708 8536 1760
rect 11704 1708 11756 1760
rect 8668 1640 8720 1692
rect 24860 1708 24912 1760
rect 25780 1708 25832 1760
rect 27620 1708 27672 1760
rect 18788 1640 18840 1692
rect 19984 1640 20036 1692
rect 23020 1640 23072 1692
rect 30472 1640 30524 1692
rect 6276 1572 6328 1624
rect 12256 1572 12308 1624
rect 16212 1572 16264 1624
rect 29092 1572 29144 1624
rect 19432 1504 19484 1556
rect 31668 1504 31720 1556
<< metal2 >>
rect 662 39200 718 39800
rect 1950 39200 2006 39800
rect 2594 39200 2650 39800
rect 2962 39536 3018 39545
rect 2962 39471 3018 39480
rect 676 36922 704 39200
rect 1766 37496 1822 37505
rect 1766 37431 1822 37440
rect 664 36916 716 36922
rect 664 36858 716 36864
rect 1780 36378 1808 37431
rect 1964 37330 1992 39200
rect 1952 37324 2004 37330
rect 1952 37266 2004 37272
rect 2504 37256 2556 37262
rect 2504 37198 2556 37204
rect 1860 36644 1912 36650
rect 1860 36586 1912 36592
rect 1768 36372 1820 36378
rect 1768 36314 1820 36320
rect 1584 36168 1636 36174
rect 1584 36110 1636 36116
rect 1766 36136 1822 36145
rect 1492 29640 1544 29646
rect 1492 29582 1544 29588
rect 1504 19514 1532 29582
rect 1596 28506 1624 36110
rect 1766 36071 1822 36080
rect 1780 35698 1808 36071
rect 1872 35894 1900 36586
rect 1872 35866 2268 35894
rect 1768 35692 1820 35698
rect 1768 35634 1820 35640
rect 1768 34400 1820 34406
rect 1768 34342 1820 34348
rect 1780 34105 1808 34342
rect 1766 34096 1822 34105
rect 1766 34031 1822 34040
rect 1768 32768 1820 32774
rect 1766 32736 1768 32745
rect 1820 32736 1822 32745
rect 1766 32671 1822 32680
rect 1860 32428 1912 32434
rect 1860 32370 1912 32376
rect 1768 32224 1820 32230
rect 1768 32166 1820 32172
rect 1780 32065 1808 32166
rect 1766 32056 1822 32065
rect 1766 31991 1822 32000
rect 1766 30696 1822 30705
rect 1766 30631 1822 30640
rect 1780 30598 1808 30631
rect 1768 30592 1820 30598
rect 1768 30534 1820 30540
rect 1768 29504 1820 29510
rect 1768 29446 1820 29452
rect 1780 29345 1808 29446
rect 1766 29336 1822 29345
rect 1766 29271 1822 29280
rect 1768 29164 1820 29170
rect 1768 29106 1820 29112
rect 1780 28665 1808 29106
rect 1766 28656 1822 28665
rect 1766 28591 1822 28600
rect 1596 28478 1808 28506
rect 1584 27464 1636 27470
rect 1584 27406 1636 27412
rect 1596 27305 1624 27406
rect 1582 27296 1638 27305
rect 1582 27231 1638 27240
rect 1676 26308 1728 26314
rect 1676 26250 1728 26256
rect 1688 25945 1716 26250
rect 1780 25974 1808 28478
rect 1768 25968 1820 25974
rect 1674 25936 1730 25945
rect 1768 25910 1820 25916
rect 1674 25871 1730 25880
rect 1768 24608 1820 24614
rect 1766 24576 1768 24585
rect 1820 24576 1822 24585
rect 1872 24562 1900 32370
rect 1952 29028 2004 29034
rect 1952 28970 2004 28976
rect 1964 25294 1992 28970
rect 1952 25288 2004 25294
rect 1952 25230 2004 25236
rect 2136 25288 2188 25294
rect 2136 25230 2188 25236
rect 1872 24534 2084 24562
rect 1766 24511 1822 24520
rect 1584 24200 1636 24206
rect 1584 24142 1636 24148
rect 1860 24200 1912 24206
rect 1860 24142 1912 24148
rect 1596 23905 1624 24142
rect 1582 23896 1638 23905
rect 1872 23866 1900 24142
rect 1582 23831 1638 23840
rect 1860 23860 1912 23866
rect 1860 23802 1912 23808
rect 1952 23520 2004 23526
rect 1950 23488 1952 23497
rect 2004 23488 2006 23497
rect 1950 23423 2006 23432
rect 2056 22778 2084 24534
rect 2148 23730 2176 25230
rect 2136 23724 2188 23730
rect 2136 23666 2188 23672
rect 2044 22772 2096 22778
rect 2044 22714 2096 22720
rect 1768 22636 1820 22642
rect 1768 22578 1820 22584
rect 1780 22545 1808 22578
rect 1766 22536 1822 22545
rect 1766 22471 1822 22480
rect 1676 21548 1728 21554
rect 1676 21490 1728 21496
rect 1688 21185 1716 21490
rect 1674 21176 1730 21185
rect 2240 21146 2268 35866
rect 2516 32910 2544 37198
rect 2608 36802 2636 39200
rect 2870 38856 2926 38865
rect 2870 38791 2926 38800
rect 2608 36786 2820 36802
rect 2608 36780 2832 36786
rect 2608 36774 2780 36780
rect 2780 36722 2832 36728
rect 2884 36174 2912 38791
rect 2976 36854 3004 39471
rect 3882 39200 3938 39800
rect 5170 39200 5226 39800
rect 5814 39200 5870 39800
rect 7102 39200 7158 39800
rect 8390 39200 8446 39800
rect 9034 39200 9090 39800
rect 10322 39200 10378 39800
rect 11610 39200 11666 39800
rect 12254 39200 12310 39800
rect 13542 39200 13598 39800
rect 14830 39200 14886 39800
rect 14936 39222 15148 39250
rect 3896 37330 3924 39200
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 3884 37324 3936 37330
rect 3884 37266 3936 37272
rect 5184 37262 5212 39200
rect 5828 37262 5856 39200
rect 7116 37262 7144 39200
rect 8404 37330 8432 39200
rect 8392 37324 8444 37330
rect 8392 37266 8444 37272
rect 5172 37256 5224 37262
rect 5172 37198 5224 37204
rect 5816 37256 5868 37262
rect 5816 37198 5868 37204
rect 7104 37256 7156 37262
rect 7104 37198 7156 37204
rect 8300 37256 8352 37262
rect 8300 37198 8352 37204
rect 6184 37120 6236 37126
rect 6184 37062 6236 37068
rect 6552 37120 6604 37126
rect 6552 37062 6604 37068
rect 7932 37120 7984 37126
rect 7932 37062 7984 37068
rect 2964 36848 3016 36854
rect 2964 36790 3016 36796
rect 3240 36576 3292 36582
rect 3240 36518 3292 36524
rect 2872 36168 2924 36174
rect 2872 36110 2924 36116
rect 3252 34610 3280 36518
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 5540 35488 5592 35494
rect 5540 35430 5592 35436
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 3056 34604 3108 34610
rect 3056 34546 3108 34552
rect 3240 34604 3292 34610
rect 3240 34546 3292 34552
rect 2504 32904 2556 32910
rect 2504 32846 2556 32852
rect 2516 26382 2544 32846
rect 3068 30938 3096 34546
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 3056 30932 3108 30938
rect 3056 30874 3108 30880
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 5552 28082 5580 35430
rect 6196 31414 6224 37062
rect 6564 36922 6592 37062
rect 6552 36916 6604 36922
rect 6552 36858 6604 36864
rect 6552 36576 6604 36582
rect 6552 36518 6604 36524
rect 6460 36032 6512 36038
rect 6460 35974 6512 35980
rect 6184 31408 6236 31414
rect 6184 31350 6236 31356
rect 6276 30660 6328 30666
rect 6276 30602 6328 30608
rect 6288 28762 6316 30602
rect 6472 30258 6500 35974
rect 6564 31346 6592 36518
rect 6736 34536 6788 34542
rect 6736 34478 6788 34484
rect 6552 31340 6604 31346
rect 6552 31282 6604 31288
rect 6460 30252 6512 30258
rect 6460 30194 6512 30200
rect 6644 30048 6696 30054
rect 6644 29990 6696 29996
rect 6276 28756 6328 28762
rect 6276 28698 6328 28704
rect 5540 28076 5592 28082
rect 5540 28018 5592 28024
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 5540 27464 5592 27470
rect 5540 27406 5592 27412
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 2504 26376 2556 26382
rect 2504 26318 2556 26324
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4068 24812 4120 24818
rect 4068 24754 4120 24760
rect 4080 23594 4108 24754
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4068 23588 4120 23594
rect 4068 23530 4120 23536
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 1674 21111 1730 21120
rect 2228 21140 2280 21146
rect 2228 21082 2280 21088
rect 4804 21004 4856 21010
rect 4804 20946 4856 20952
rect 1584 20936 1636 20942
rect 1584 20878 1636 20884
rect 1860 20936 1912 20942
rect 1860 20878 1912 20884
rect 1596 20505 1624 20878
rect 1872 20534 1900 20878
rect 4528 20868 4580 20874
rect 4528 20810 4580 20816
rect 4540 20777 4568 20810
rect 4526 20768 4582 20777
rect 4526 20703 4582 20712
rect 1860 20528 1912 20534
rect 1582 20496 1638 20505
rect 1860 20470 1912 20476
rect 1582 20431 1638 20440
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 3976 19780 4028 19786
rect 3976 19722 4028 19728
rect 1492 19508 1544 19514
rect 1492 19450 1544 19456
rect 1860 19372 1912 19378
rect 1860 19314 1912 19320
rect 1766 19136 1822 19145
rect 1766 19071 1822 19080
rect 1780 18766 1808 19071
rect 1768 18760 1820 18766
rect 1768 18702 1820 18708
rect 1584 18216 1636 18222
rect 1584 18158 1636 18164
rect 1596 17785 1624 18158
rect 1582 17776 1638 17785
rect 1872 17746 1900 19314
rect 1582 17711 1638 17720
rect 1860 17740 1912 17746
rect 1860 17682 1912 17688
rect 1768 17196 1820 17202
rect 1768 17138 1820 17144
rect 1780 17105 1808 17138
rect 1766 17096 1822 17105
rect 1766 17031 1822 17040
rect 1584 16992 1636 16998
rect 1584 16934 1636 16940
rect 1596 16658 1624 16934
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 1492 16040 1544 16046
rect 1492 15982 1544 15988
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1412 6905 1440 8434
rect 1398 6896 1454 6905
rect 1398 6831 1454 6840
rect 1504 6662 1532 15982
rect 1768 15904 1820 15910
rect 1768 15846 1820 15852
rect 1780 15745 1808 15846
rect 1766 15736 1822 15745
rect 1766 15671 1822 15680
rect 1676 15496 1728 15502
rect 1676 15438 1728 15444
rect 1688 15026 1716 15438
rect 1676 15020 1728 15026
rect 1676 14962 1728 14968
rect 1584 13932 1636 13938
rect 1584 13874 1636 13880
rect 1596 8401 1624 13874
rect 1582 8392 1638 8401
rect 1582 8327 1638 8336
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1492 6656 1544 6662
rect 1492 6598 1544 6604
rect 1596 5545 1624 7822
rect 1688 6769 1716 14962
rect 1872 14618 1900 17682
rect 1952 17060 2004 17066
rect 1952 17002 2004 17008
rect 1860 14612 1912 14618
rect 1860 14554 1912 14560
rect 1768 14408 1820 14414
rect 1766 14376 1768 14385
rect 1820 14376 1822 14385
rect 1766 14311 1822 14320
rect 1768 13728 1820 13734
rect 1766 13696 1768 13705
rect 1820 13696 1822 13705
rect 1766 13631 1822 13640
rect 1860 12844 1912 12850
rect 1860 12786 1912 12792
rect 1768 12640 1820 12646
rect 1768 12582 1820 12588
rect 1780 12345 1808 12582
rect 1766 12336 1822 12345
rect 1766 12271 1822 12280
rect 1768 11144 1820 11150
rect 1768 11086 1820 11092
rect 1780 10985 1808 11086
rect 1766 10976 1822 10985
rect 1766 10911 1822 10920
rect 1768 10668 1820 10674
rect 1768 10610 1820 10616
rect 1780 10305 1808 10610
rect 1766 10296 1822 10305
rect 1766 10231 1822 10240
rect 1766 8936 1822 8945
rect 1766 8871 1822 8880
rect 1780 8838 1808 8871
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 1872 8634 1900 12786
rect 1964 10810 1992 17002
rect 3700 16788 3752 16794
rect 3700 16730 3752 16736
rect 2504 16108 2556 16114
rect 2504 16050 2556 16056
rect 2516 15706 2544 16050
rect 2596 15904 2648 15910
rect 2596 15846 2648 15852
rect 2504 15700 2556 15706
rect 2504 15642 2556 15648
rect 2412 15360 2464 15366
rect 2412 15302 2464 15308
rect 2424 15026 2452 15302
rect 2608 15026 2636 15846
rect 3608 15428 3660 15434
rect 3608 15370 3660 15376
rect 2412 15020 2464 15026
rect 2412 14962 2464 14968
rect 2596 15020 2648 15026
rect 2596 14962 2648 14968
rect 2688 14816 2740 14822
rect 2688 14758 2740 14764
rect 3056 14816 3108 14822
rect 3056 14758 3108 14764
rect 2700 14482 2728 14758
rect 3068 14618 3096 14758
rect 3056 14612 3108 14618
rect 3056 14554 3108 14560
rect 2688 14476 2740 14482
rect 2688 14418 2740 14424
rect 2504 14408 2556 14414
rect 2504 14350 2556 14356
rect 2320 11008 2372 11014
rect 2320 10950 2372 10956
rect 1952 10804 2004 10810
rect 1952 10746 2004 10752
rect 1952 10600 2004 10606
rect 1952 10542 2004 10548
rect 1860 8628 1912 8634
rect 1860 8570 1912 8576
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 1766 7576 1822 7585
rect 1766 7511 1822 7520
rect 1780 6798 1808 7511
rect 1768 6792 1820 6798
rect 1674 6760 1730 6769
rect 1768 6734 1820 6740
rect 1674 6695 1730 6704
rect 1582 5536 1638 5545
rect 1582 5471 1638 5480
rect 1582 5400 1638 5409
rect 1582 5335 1638 5344
rect 1596 4622 1624 5335
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 1768 4480 1820 4486
rect 1768 4422 1820 4428
rect 1780 4185 1808 4422
rect 1766 4176 1822 4185
rect 1766 4111 1822 4120
rect 1766 3496 1822 3505
rect 1766 3431 1822 3440
rect 1780 3398 1808 3431
rect 1768 3392 1820 3398
rect 1768 3334 1820 3340
rect 664 2848 716 2854
rect 664 2790 716 2796
rect 20 2576 72 2582
rect 20 2518 72 2524
rect 32 800 60 2518
rect 676 800 704 2790
rect 1674 2680 1730 2689
rect 1674 2615 1730 2624
rect 1688 2446 1716 2615
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 1872 2145 1900 8434
rect 1964 8090 1992 10542
rect 2228 9648 2280 9654
rect 2228 9590 2280 9596
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 2148 7426 2176 9522
rect 2240 8634 2268 9590
rect 2332 9178 2360 10950
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 2228 8628 2280 8634
rect 2228 8570 2280 8576
rect 2148 7398 2268 7426
rect 2240 7342 2268 7398
rect 1952 7336 2004 7342
rect 1952 7278 2004 7284
rect 2136 7336 2188 7342
rect 2136 7278 2188 7284
rect 2228 7336 2280 7342
rect 2228 7278 2280 7284
rect 1964 6934 1992 7278
rect 1952 6928 2004 6934
rect 1952 6870 2004 6876
rect 2148 5370 2176 7278
rect 2332 6914 2360 9114
rect 2516 7546 2544 14350
rect 3068 14006 3096 14554
rect 3516 14068 3568 14074
rect 3516 14010 3568 14016
rect 3056 14000 3108 14006
rect 3056 13942 3108 13948
rect 3240 12912 3292 12918
rect 3240 12854 3292 12860
rect 2964 12368 3016 12374
rect 2964 12310 3016 12316
rect 2596 12096 2648 12102
rect 2596 12038 2648 12044
rect 2608 9586 2636 12038
rect 2780 10668 2832 10674
rect 2780 10610 2832 10616
rect 2792 10062 2820 10610
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2596 9580 2648 9586
rect 2596 9522 2648 9528
rect 2596 9104 2648 9110
rect 2596 9046 2648 9052
rect 2504 7540 2556 7546
rect 2504 7482 2556 7488
rect 2608 7426 2636 9046
rect 2976 8974 3004 12310
rect 3252 9586 3280 12854
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 3252 9058 3280 9522
rect 3330 9480 3386 9489
rect 3330 9415 3332 9424
rect 3384 9415 3386 9424
rect 3332 9386 3384 9392
rect 3252 9030 3372 9058
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 2872 8832 2924 8838
rect 2872 8774 2924 8780
rect 2688 7540 2740 7546
rect 2688 7482 2740 7488
rect 2516 7398 2636 7426
rect 2332 6886 2452 6914
rect 2228 6792 2280 6798
rect 2228 6734 2280 6740
rect 2240 6254 2268 6734
rect 2228 6248 2280 6254
rect 2228 6190 2280 6196
rect 2240 5914 2268 6190
rect 2228 5908 2280 5914
rect 2228 5850 2280 5856
rect 2424 5710 2452 6886
rect 2228 5704 2280 5710
rect 2228 5646 2280 5652
rect 2412 5704 2464 5710
rect 2412 5646 2464 5652
rect 2136 5364 2188 5370
rect 2136 5306 2188 5312
rect 2240 5302 2268 5646
rect 2228 5296 2280 5302
rect 2228 5238 2280 5244
rect 2320 5228 2372 5234
rect 2320 5170 2372 5176
rect 2226 3632 2282 3641
rect 2226 3567 2228 3576
rect 2280 3567 2282 3576
rect 2228 3538 2280 3544
rect 1952 2304 2004 2310
rect 1952 2246 2004 2252
rect 1858 2136 1914 2145
rect 1858 2071 1914 2080
rect 1964 800 1992 2246
rect 2332 1766 2360 5170
rect 2412 3120 2464 3126
rect 2410 3088 2412 3097
rect 2464 3088 2466 3097
rect 2410 3023 2466 3032
rect 2516 2446 2544 7398
rect 2596 7336 2648 7342
rect 2596 7278 2648 7284
rect 2608 3534 2636 7278
rect 2700 7002 2728 7482
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2688 6996 2740 7002
rect 2688 6938 2740 6944
rect 2596 3528 2648 3534
rect 2596 3470 2648 3476
rect 2792 3194 2820 7142
rect 2884 6866 2912 8774
rect 2872 6860 2924 6866
rect 2872 6802 2924 6808
rect 2976 6730 3004 8910
rect 3056 8492 3108 8498
rect 3056 8434 3108 8440
rect 2964 6724 3016 6730
rect 2964 6666 3016 6672
rect 2964 6384 3016 6390
rect 2964 6326 3016 6332
rect 2976 5370 3004 6326
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 2872 5024 2924 5030
rect 2872 4966 2924 4972
rect 2780 3188 2832 3194
rect 2780 3130 2832 3136
rect 2884 3058 2912 4966
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 2976 3398 3004 3878
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 2504 2440 2556 2446
rect 2504 2382 2556 2388
rect 2320 1760 2372 1766
rect 2320 1702 2372 1708
rect 3068 921 3096 8434
rect 3148 7744 3200 7750
rect 3148 7686 3200 7692
rect 3160 3369 3188 7686
rect 3252 5846 3280 8910
rect 3344 6798 3372 9030
rect 3424 7744 3476 7750
rect 3424 7686 3476 7692
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 3240 5840 3292 5846
rect 3240 5782 3292 5788
rect 3344 5710 3372 6734
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 3330 5536 3386 5545
rect 3330 5471 3386 5480
rect 3344 5234 3372 5471
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 3238 4720 3294 4729
rect 3238 4655 3294 4664
rect 3252 4622 3280 4655
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 3252 4214 3280 4558
rect 3240 4208 3292 4214
rect 3240 4150 3292 4156
rect 3240 4072 3292 4078
rect 3240 4014 3292 4020
rect 3146 3360 3202 3369
rect 3146 3295 3202 3304
rect 3146 3224 3202 3233
rect 3146 3159 3148 3168
rect 3200 3159 3202 3168
rect 3148 3130 3200 3136
rect 3252 3058 3280 4014
rect 3240 3052 3292 3058
rect 3240 2994 3292 3000
rect 3146 2680 3202 2689
rect 3146 2615 3202 2624
rect 3160 2446 3188 2615
rect 3148 2440 3200 2446
rect 3148 2382 3200 2388
rect 3240 2304 3292 2310
rect 3240 2246 3292 2252
rect 3054 912 3110 921
rect 3054 847 3110 856
rect 3252 800 3280 2246
rect 3436 2106 3464 7686
rect 3528 4146 3556 14010
rect 3620 12646 3648 15370
rect 3712 13841 3740 16730
rect 3792 14816 3844 14822
rect 3792 14758 3844 14764
rect 3698 13832 3754 13841
rect 3698 13767 3754 13776
rect 3608 12640 3660 12646
rect 3608 12582 3660 12588
rect 3804 9761 3832 14758
rect 3988 12986 4016 19722
rect 4816 19242 4844 20946
rect 5080 19780 5132 19786
rect 5080 19722 5132 19728
rect 5092 19514 5120 19722
rect 5080 19508 5132 19514
rect 5080 19450 5132 19456
rect 5552 19394 5580 27406
rect 5632 21480 5684 21486
rect 5632 21422 5684 21428
rect 5644 21010 5672 21422
rect 5632 21004 5684 21010
rect 5632 20946 5684 20952
rect 5552 19378 5672 19394
rect 5552 19372 5684 19378
rect 5552 19366 5632 19372
rect 5632 19314 5684 19320
rect 4804 19236 4856 19242
rect 4804 19178 4856 19184
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4816 18358 4844 19178
rect 5448 18624 5500 18630
rect 5448 18566 5500 18572
rect 5460 18358 5488 18566
rect 5644 18442 5672 19314
rect 5816 19304 5868 19310
rect 5816 19246 5868 19252
rect 5724 19168 5776 19174
rect 5724 19110 5776 19116
rect 5552 18414 5672 18442
rect 4620 18352 4672 18358
rect 4620 18294 4672 18300
rect 4804 18352 4856 18358
rect 4804 18294 4856 18300
rect 5448 18352 5500 18358
rect 5448 18294 5500 18300
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4632 17882 4660 18294
rect 4620 17876 4672 17882
rect 4620 17818 4672 17824
rect 5172 17876 5224 17882
rect 5172 17818 5224 17824
rect 4252 17672 4304 17678
rect 4250 17640 4252 17649
rect 4304 17640 4306 17649
rect 4250 17575 4306 17584
rect 4252 17536 4304 17542
rect 4252 17478 4304 17484
rect 4264 17270 4292 17478
rect 5184 17270 5212 17818
rect 5448 17672 5500 17678
rect 5448 17614 5500 17620
rect 4252 17264 4304 17270
rect 4252 17206 4304 17212
rect 5172 17264 5224 17270
rect 5172 17206 5224 17212
rect 4804 17128 4856 17134
rect 4804 17070 4856 17076
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4068 16108 4120 16114
rect 4068 16050 4120 16056
rect 4080 14074 4108 16050
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4712 14408 4764 14414
rect 4710 14376 4712 14385
rect 4764 14376 4766 14385
rect 4710 14311 4766 14320
rect 4712 14272 4764 14278
rect 4712 14214 4764 14220
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 4620 13932 4672 13938
rect 4620 13874 4672 13880
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4632 13394 4660 13874
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 4724 13326 4752 14214
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4620 13184 4672 13190
rect 4620 13126 4672 13132
rect 4712 13184 4764 13190
rect 4712 13126 4764 13132
rect 3976 12980 4028 12986
rect 3976 12922 4028 12928
rect 3976 12640 4028 12646
rect 3976 12582 4028 12588
rect 3884 9988 3936 9994
rect 3884 9930 3936 9936
rect 3790 9752 3846 9761
rect 3790 9687 3846 9696
rect 3896 9586 3924 9930
rect 3884 9580 3936 9586
rect 3884 9522 3936 9528
rect 3792 9512 3844 9518
rect 3792 9454 3844 9460
rect 3988 9466 4016 12582
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4540 9625 4568 9658
rect 4526 9616 4582 9625
rect 4252 9580 4304 9586
rect 4526 9551 4582 9560
rect 4252 9522 4304 9528
rect 4160 9512 4212 9518
rect 3988 9460 4160 9466
rect 3988 9454 4212 9460
rect 3608 7948 3660 7954
rect 3608 7890 3660 7896
rect 3620 5234 3648 7890
rect 3698 7440 3754 7449
rect 3698 7375 3700 7384
rect 3752 7375 3754 7384
rect 3700 7346 3752 7352
rect 3700 6724 3752 6730
rect 3700 6666 3752 6672
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3712 4214 3740 6666
rect 3804 5273 3832 9454
rect 3988 9438 4200 9454
rect 4264 9364 4292 9522
rect 4080 9336 4292 9364
rect 4080 9081 4108 9336
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4528 9172 4580 9178
rect 4528 9114 4580 9120
rect 4066 9072 4122 9081
rect 4066 9007 4122 9016
rect 4540 8566 4568 9114
rect 4632 8906 4660 13126
rect 4724 12646 4752 13126
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 4620 8900 4672 8906
rect 4620 8842 4672 8848
rect 4528 8560 4580 8566
rect 4528 8502 4580 8508
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 3790 5264 3846 5273
rect 3790 5199 3846 5208
rect 3792 4752 3844 4758
rect 3792 4694 3844 4700
rect 3700 4208 3752 4214
rect 3804 4185 3832 4694
rect 3700 4150 3752 4156
rect 3790 4176 3846 4185
rect 3516 4140 3568 4146
rect 3516 4082 3568 4088
rect 3712 3534 3740 4150
rect 3790 4111 3846 4120
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 3804 3194 3832 3878
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 3424 2100 3476 2106
rect 3424 2042 3476 2048
rect 3804 2038 3832 2994
rect 3792 2032 3844 2038
rect 3792 1974 3844 1980
rect 3896 800 3924 8434
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 3988 7886 4016 8230
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4068 8016 4120 8022
rect 4066 7984 4068 7993
rect 4120 7984 4122 7993
rect 4066 7919 4122 7928
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 4620 7812 4672 7818
rect 4620 7754 4672 7760
rect 4526 7712 4582 7721
rect 4526 7647 4582 7656
rect 4540 7274 4568 7647
rect 4528 7268 4580 7274
rect 4528 7210 4580 7216
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4342 6896 4398 6905
rect 4342 6831 4398 6840
rect 4356 6798 4384 6831
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 4068 6384 4120 6390
rect 4066 6352 4068 6361
rect 4120 6352 4122 6361
rect 4066 6287 4122 6296
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4632 5794 4660 7754
rect 4724 7478 4752 12582
rect 4816 10810 4844 17070
rect 5264 15632 5316 15638
rect 5264 15574 5316 15580
rect 4896 15496 4948 15502
rect 4896 15438 4948 15444
rect 5080 15496 5132 15502
rect 5080 15438 5132 15444
rect 4908 14414 4936 15438
rect 5092 15094 5120 15438
rect 5172 15360 5224 15366
rect 5172 15302 5224 15308
rect 5080 15088 5132 15094
rect 5080 15030 5132 15036
rect 4988 15020 5040 15026
rect 4988 14962 5040 14968
rect 4896 14408 4948 14414
rect 4896 14350 4948 14356
rect 4908 13190 4936 14350
rect 4896 13184 4948 13190
rect 4896 13126 4948 13132
rect 4894 12880 4950 12889
rect 4894 12815 4950 12824
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 4816 10062 4844 10610
rect 4804 10056 4856 10062
rect 4804 9998 4856 10004
rect 4802 9752 4858 9761
rect 4802 9687 4804 9696
rect 4856 9687 4858 9696
rect 4804 9658 4856 9664
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4712 7472 4764 7478
rect 4712 7414 4764 7420
rect 4632 5766 4752 5794
rect 4528 5704 4580 5710
rect 4580 5664 4660 5692
rect 4528 5646 4580 5652
rect 4632 5302 4660 5664
rect 4620 5296 4672 5302
rect 4620 5238 4672 5244
rect 4528 5160 4580 5166
rect 4526 5128 4528 5137
rect 4580 5128 4582 5137
rect 4526 5063 4582 5072
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4632 4706 4660 5238
rect 4540 4678 4660 4706
rect 4540 4622 4568 4678
rect 4528 4616 4580 4622
rect 4528 4558 4580 4564
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 3974 4176 4030 4185
rect 3974 4111 4030 4120
rect 3988 3534 4016 4111
rect 4080 3738 4108 4218
rect 4540 4196 4568 4558
rect 4540 4168 4660 4196
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 4172 4049 4200 4082
rect 4158 4040 4214 4049
rect 4158 3975 4214 3984
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 4528 3732 4580 3738
rect 4632 3720 4660 4168
rect 4724 4146 4752 5766
rect 4816 4457 4844 8774
rect 4908 4690 4936 12815
rect 5000 10062 5028 14962
rect 5092 13977 5120 15030
rect 5078 13968 5134 13977
rect 5078 13903 5134 13912
rect 5092 12850 5120 13903
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 4988 10056 5040 10062
rect 4988 9998 5040 10004
rect 4988 9920 5040 9926
rect 4988 9862 5040 9868
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 5000 4570 5028 9862
rect 5092 7886 5120 12786
rect 5184 8974 5212 15302
rect 5276 13394 5304 15574
rect 5356 15360 5408 15366
rect 5356 15302 5408 15308
rect 5264 13388 5316 13394
rect 5264 13330 5316 13336
rect 5276 9058 5304 13330
rect 5368 9926 5396 15302
rect 5460 13954 5488 17614
rect 5552 14074 5580 18414
rect 5736 18222 5764 19110
rect 5828 18766 5856 19246
rect 5816 18760 5868 18766
rect 5816 18702 5868 18708
rect 5724 18216 5776 18222
rect 5724 18158 5776 18164
rect 5828 16810 5856 18702
rect 6656 18358 6684 29990
rect 6748 26450 6776 34478
rect 7944 31822 7972 37062
rect 7932 31816 7984 31822
rect 7932 31758 7984 31764
rect 8116 31816 8168 31822
rect 8116 31758 8168 31764
rect 6828 31136 6880 31142
rect 6828 31078 6880 31084
rect 7380 31136 7432 31142
rect 7380 31078 7432 31084
rect 6736 26444 6788 26450
rect 6736 26386 6788 26392
rect 6736 21616 6788 21622
rect 6736 21558 6788 21564
rect 6748 20602 6776 21558
rect 6736 20596 6788 20602
rect 6736 20538 6788 20544
rect 6736 19780 6788 19786
rect 6736 19722 6788 19728
rect 6748 19514 6776 19722
rect 6736 19508 6788 19514
rect 6736 19450 6788 19456
rect 6644 18352 6696 18358
rect 6644 18294 6696 18300
rect 6748 18170 6776 19450
rect 6656 18142 6776 18170
rect 6368 17264 6420 17270
rect 6368 17206 6420 17212
rect 5736 16782 5856 16810
rect 5632 16108 5684 16114
rect 5632 16050 5684 16056
rect 5644 14890 5672 16050
rect 5632 14884 5684 14890
rect 5632 14826 5684 14832
rect 5644 14414 5672 14826
rect 5632 14408 5684 14414
rect 5632 14350 5684 14356
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 5460 13926 5580 13954
rect 5448 13864 5500 13870
rect 5448 13806 5500 13812
rect 5460 12442 5488 13806
rect 5552 12617 5580 13926
rect 5538 12608 5594 12617
rect 5538 12543 5594 12552
rect 5448 12436 5500 12442
rect 5448 12378 5500 12384
rect 5644 11558 5672 14214
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5736 11354 5764 16782
rect 5816 15496 5868 15502
rect 5816 15438 5868 15444
rect 5828 15026 5856 15438
rect 5816 15020 5868 15026
rect 5816 14962 5868 14968
rect 6000 15020 6052 15026
rect 6000 14962 6052 14968
rect 5828 13326 5856 14962
rect 5908 14816 5960 14822
rect 5908 14758 5960 14764
rect 5920 13530 5948 14758
rect 5908 13524 5960 13530
rect 5908 13466 5960 13472
rect 5816 13320 5868 13326
rect 5816 13262 5868 13268
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 5356 9920 5408 9926
rect 5356 9862 5408 9868
rect 5276 9030 5396 9058
rect 5172 8968 5224 8974
rect 5172 8910 5224 8916
rect 5264 8900 5316 8906
rect 5264 8842 5316 8848
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 5080 7880 5132 7886
rect 5080 7822 5132 7828
rect 5092 7410 5120 7822
rect 5080 7404 5132 7410
rect 5080 7346 5132 7352
rect 5078 7304 5134 7313
rect 5078 7239 5080 7248
rect 5132 7239 5134 7248
rect 5080 7210 5132 7216
rect 5080 6792 5132 6798
rect 5080 6734 5132 6740
rect 5092 6633 5120 6734
rect 5078 6624 5134 6633
rect 5078 6559 5134 6568
rect 5184 6202 5212 8774
rect 5092 6174 5212 6202
rect 5092 4865 5120 6174
rect 5276 5642 5304 8842
rect 5368 7750 5396 9030
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 5354 7576 5410 7585
rect 5354 7511 5410 7520
rect 5368 7478 5396 7511
rect 5356 7472 5408 7478
rect 5356 7414 5408 7420
rect 5460 7290 5488 9998
rect 5552 9722 5580 10066
rect 5828 10062 5856 13262
rect 5908 12844 5960 12850
rect 5908 12786 5960 12792
rect 5920 12374 5948 12786
rect 5908 12368 5960 12374
rect 5908 12310 5960 12316
rect 6012 11082 6040 14962
rect 6090 14512 6146 14521
rect 6090 14447 6146 14456
rect 6104 13938 6132 14447
rect 6276 14408 6328 14414
rect 6196 14368 6276 14396
rect 6092 13932 6144 13938
rect 6092 13874 6144 13880
rect 6196 13818 6224 14368
rect 6276 14350 6328 14356
rect 6104 13790 6224 13818
rect 6000 11076 6052 11082
rect 6000 11018 6052 11024
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 6104 9994 6132 13790
rect 6184 13728 6236 13734
rect 6184 13670 6236 13676
rect 6196 12850 6224 13670
rect 6184 12844 6236 12850
rect 6184 12786 6236 12792
rect 6182 12608 6238 12617
rect 6182 12543 6238 12552
rect 5724 9988 5776 9994
rect 5724 9930 5776 9936
rect 6092 9988 6144 9994
rect 6092 9930 6144 9936
rect 5540 9716 5592 9722
rect 5540 9658 5592 9664
rect 5632 9444 5684 9450
rect 5632 9386 5684 9392
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 5552 8090 5580 8502
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5368 7262 5488 7290
rect 5264 5636 5316 5642
rect 5264 5578 5316 5584
rect 5368 5114 5396 7262
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 5460 6934 5488 7142
rect 5448 6928 5500 6934
rect 5448 6870 5500 6876
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5552 6322 5580 6734
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5368 5098 5580 5114
rect 5368 5092 5592 5098
rect 5368 5086 5540 5092
rect 5540 5034 5592 5040
rect 5078 4856 5134 4865
rect 5078 4791 5134 4800
rect 4908 4542 5028 4570
rect 4802 4448 4858 4457
rect 4802 4383 4858 4392
rect 4712 4140 4764 4146
rect 4712 4082 4764 4088
rect 4580 3692 4660 3720
rect 4528 3674 4580 3680
rect 4540 3602 4568 3674
rect 4528 3596 4580 3602
rect 4528 3538 4580 3544
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 4526 3496 4582 3505
rect 4526 3431 4582 3440
rect 4540 2990 4568 3431
rect 4632 3126 4660 3538
rect 4804 3460 4856 3466
rect 4724 3420 4804 3448
rect 4620 3120 4672 3126
rect 4620 3062 4672 3068
rect 4528 2984 4580 2990
rect 4528 2926 4580 2932
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2514 4660 3062
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 4528 2372 4580 2378
rect 4528 2314 4580 2320
rect 4540 1834 4568 2314
rect 4724 1902 4752 3420
rect 4804 3402 4856 3408
rect 4804 3120 4856 3126
rect 4908 3108 4936 4542
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 5172 3936 5224 3942
rect 5172 3878 5224 3884
rect 4988 3460 5040 3466
rect 4988 3402 5040 3408
rect 4856 3080 4936 3108
rect 4804 3062 4856 3068
rect 5000 2650 5028 3402
rect 5092 2990 5120 3878
rect 5080 2984 5132 2990
rect 5080 2926 5132 2932
rect 4988 2644 5040 2650
rect 4988 2586 5040 2592
rect 4712 1896 4764 1902
rect 4712 1838 4764 1844
rect 4528 1828 4580 1834
rect 4528 1770 4580 1776
rect 5184 800 5212 3878
rect 5644 3466 5672 9386
rect 5736 6798 5764 9930
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5736 4593 5764 6258
rect 5722 4584 5778 4593
rect 5828 4554 5856 9318
rect 6196 9058 6224 12543
rect 6012 9030 6224 9058
rect 5908 8016 5960 8022
rect 5908 7958 5960 7964
rect 5920 6458 5948 7958
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 6012 5914 6040 9030
rect 6276 8900 6328 8906
rect 6276 8842 6328 8848
rect 6288 7954 6316 8842
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 6092 7744 6144 7750
rect 6092 7686 6144 7692
rect 6000 5908 6052 5914
rect 6000 5850 6052 5856
rect 6104 5302 6132 7686
rect 6184 6928 6236 6934
rect 6184 6870 6236 6876
rect 6092 5296 6144 5302
rect 6092 5238 6144 5244
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 5908 5024 5960 5030
rect 5908 4966 5960 4972
rect 5920 4758 5948 4966
rect 5908 4752 5960 4758
rect 6012 4729 6040 5170
rect 5908 4694 5960 4700
rect 5998 4720 6054 4729
rect 5998 4655 6054 4664
rect 5722 4519 5778 4528
rect 5816 4548 5868 4554
rect 5816 4490 5868 4496
rect 6196 4321 6224 6870
rect 6274 5944 6330 5953
rect 6274 5879 6276 5888
rect 6328 5879 6330 5888
rect 6276 5850 6328 5856
rect 6182 4312 6238 4321
rect 6182 4247 6238 4256
rect 5816 4208 5868 4214
rect 5816 4150 5868 4156
rect 5632 3460 5684 3466
rect 5632 3402 5684 3408
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5552 2310 5580 3130
rect 5828 2378 5856 4150
rect 5816 2372 5868 2378
rect 5816 2314 5868 2320
rect 5540 2304 5592 2310
rect 5540 2246 5592 2252
rect 6288 1630 6316 5850
rect 6380 3194 6408 17206
rect 6552 15904 6604 15910
rect 6552 15846 6604 15852
rect 6460 15700 6512 15706
rect 6460 15642 6512 15648
rect 6472 15502 6500 15642
rect 6460 15496 6512 15502
rect 6460 15438 6512 15444
rect 6472 14414 6500 15438
rect 6460 14408 6512 14414
rect 6460 14350 6512 14356
rect 6460 11280 6512 11286
rect 6458 11248 6460 11257
rect 6512 11248 6514 11257
rect 6458 11183 6514 11192
rect 6564 11082 6592 15846
rect 6552 11076 6604 11082
rect 6552 11018 6604 11024
rect 6460 10192 6512 10198
rect 6460 10134 6512 10140
rect 6472 4214 6500 10134
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6564 9761 6592 9998
rect 6550 9752 6606 9761
rect 6550 9687 6606 9696
rect 6564 7886 6592 9687
rect 6656 8566 6684 18142
rect 6840 16726 6868 31078
rect 7012 23724 7064 23730
rect 7012 23666 7064 23672
rect 7024 22098 7052 23666
rect 7012 22092 7064 22098
rect 7012 22034 7064 22040
rect 7104 22024 7156 22030
rect 7104 21966 7156 21972
rect 7116 21554 7144 21966
rect 7392 21622 7420 31078
rect 7564 22568 7616 22574
rect 7564 22510 7616 22516
rect 7472 21888 7524 21894
rect 7472 21830 7524 21836
rect 7484 21622 7512 21830
rect 7380 21616 7432 21622
rect 7380 21558 7432 21564
rect 7472 21616 7524 21622
rect 7472 21558 7524 21564
rect 7104 21548 7156 21554
rect 7104 21490 7156 21496
rect 6920 21412 6972 21418
rect 6920 21354 6972 21360
rect 6932 19310 6960 21354
rect 7116 20330 7144 21490
rect 7472 20936 7524 20942
rect 7472 20878 7524 20884
rect 7104 20324 7156 20330
rect 7104 20266 7156 20272
rect 7116 19990 7144 20266
rect 7104 19984 7156 19990
rect 7104 19926 7156 19932
rect 7116 19310 7144 19926
rect 6920 19304 6972 19310
rect 6920 19246 6972 19252
rect 7104 19304 7156 19310
rect 7104 19246 7156 19252
rect 6932 18222 6960 19246
rect 7012 18624 7064 18630
rect 7012 18566 7064 18572
rect 7104 18624 7156 18630
rect 7104 18566 7156 18572
rect 6920 18216 6972 18222
rect 6920 18158 6972 18164
rect 6828 16720 6880 16726
rect 6828 16662 6880 16668
rect 7024 16658 7052 18566
rect 7012 16652 7064 16658
rect 7012 16594 7064 16600
rect 7116 16522 7144 18566
rect 7104 16516 7156 16522
rect 7104 16458 7156 16464
rect 7380 16176 7432 16182
rect 7380 16118 7432 16124
rect 6736 16108 6788 16114
rect 6736 16050 6788 16056
rect 7288 16108 7340 16114
rect 7288 16050 7340 16056
rect 6748 13734 6776 16050
rect 6828 15360 6880 15366
rect 6828 15302 6880 15308
rect 7196 15360 7248 15366
rect 7196 15302 7248 15308
rect 6736 13728 6788 13734
rect 6736 13670 6788 13676
rect 6840 13569 6868 15302
rect 7104 14340 7156 14346
rect 7104 14282 7156 14288
rect 6920 14272 6972 14278
rect 6920 14214 6972 14220
rect 6932 14074 6960 14214
rect 6920 14068 6972 14074
rect 6920 14010 6972 14016
rect 6918 13968 6974 13977
rect 6918 13903 6920 13912
rect 6972 13903 6974 13912
rect 6920 13874 6972 13880
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 6826 13560 6882 13569
rect 6826 13495 6882 13504
rect 6826 13424 6882 13433
rect 6736 13388 6788 13394
rect 6826 13359 6882 13368
rect 6736 13330 6788 13336
rect 6748 12306 6776 13330
rect 6840 12850 6868 13359
rect 6828 12844 6880 12850
rect 6828 12786 6880 12792
rect 6932 12714 6960 13670
rect 7012 13252 7064 13258
rect 7012 13194 7064 13200
rect 6920 12708 6972 12714
rect 6920 12650 6972 12656
rect 6736 12300 6788 12306
rect 6736 12242 6788 12248
rect 6748 11218 6776 12242
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6840 10062 6868 10542
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6840 9518 6868 9998
rect 7024 9994 7052 13194
rect 7116 12170 7144 14282
rect 7208 13734 7236 15302
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 7196 13252 7248 13258
rect 7196 13194 7248 13200
rect 7208 12850 7236 13194
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7104 12164 7156 12170
rect 7104 12106 7156 12112
rect 7012 9988 7064 9994
rect 7012 9930 7064 9936
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6840 8974 6868 9454
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6932 9178 6960 9318
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6840 8634 6868 8910
rect 7196 8832 7248 8838
rect 7196 8774 7248 8780
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6644 8560 6696 8566
rect 6644 8502 6696 8508
rect 7208 8498 7236 8774
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6736 7948 6788 7954
rect 6736 7890 6788 7896
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6564 6934 6592 7822
rect 6748 7410 6776 7890
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6552 6928 6604 6934
rect 6552 6870 6604 6876
rect 6748 6866 6776 7346
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 6642 6080 6698 6089
rect 6564 5778 6592 6054
rect 6642 6015 6698 6024
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6550 5672 6606 5681
rect 6656 5642 6684 6015
rect 6748 5778 6776 6802
rect 6840 6662 6868 8230
rect 7116 7818 7144 8366
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 7104 7812 7156 7818
rect 7104 7754 7156 7760
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6932 5817 6960 7754
rect 7104 7200 7156 7206
rect 7104 7142 7156 7148
rect 7012 6724 7064 6730
rect 7012 6666 7064 6672
rect 6918 5808 6974 5817
rect 6736 5772 6788 5778
rect 7024 5778 7052 6666
rect 7116 6390 7144 7142
rect 7104 6384 7156 6390
rect 7104 6326 7156 6332
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 6918 5743 6974 5752
rect 7012 5772 7064 5778
rect 6736 5714 6788 5720
rect 7012 5714 7064 5720
rect 6550 5607 6606 5616
rect 6644 5636 6696 5642
rect 6460 4208 6512 4214
rect 6460 4150 6512 4156
rect 6564 3670 6592 5607
rect 6644 5578 6696 5584
rect 6748 4690 6776 5714
rect 6826 5400 6882 5409
rect 6826 5335 6882 5344
rect 6840 5098 6868 5335
rect 6918 5264 6974 5273
rect 6918 5199 6974 5208
rect 6828 5092 6880 5098
rect 6828 5034 6880 5040
rect 6736 4684 6788 4690
rect 6736 4626 6788 4632
rect 6932 4554 6960 5199
rect 6920 4548 6972 4554
rect 6920 4490 6972 4496
rect 7010 4176 7066 4185
rect 7116 4146 7144 6190
rect 7196 5568 7248 5574
rect 7196 5510 7248 5516
rect 7208 5409 7236 5510
rect 7194 5400 7250 5409
rect 7194 5335 7250 5344
rect 7196 5296 7248 5302
rect 7194 5264 7196 5273
rect 7248 5264 7250 5273
rect 7194 5199 7250 5208
rect 7196 5160 7248 5166
rect 7196 5102 7248 5108
rect 7208 4706 7236 5102
rect 7300 4842 7328 16050
rect 7392 15502 7420 16118
rect 7380 15496 7432 15502
rect 7380 15438 7432 15444
rect 7484 15026 7512 20878
rect 7576 16250 7604 22510
rect 7748 20868 7800 20874
rect 7748 20810 7800 20816
rect 7656 20460 7708 20466
rect 7656 20402 7708 20408
rect 7668 19990 7696 20402
rect 7656 19984 7708 19990
rect 7656 19926 7708 19932
rect 7656 16992 7708 16998
rect 7656 16934 7708 16940
rect 7564 16244 7616 16250
rect 7564 16186 7616 16192
rect 7562 15464 7618 15473
rect 7562 15399 7564 15408
rect 7616 15399 7618 15408
rect 7564 15370 7616 15376
rect 7472 15020 7524 15026
rect 7472 14962 7524 14968
rect 7564 14952 7616 14958
rect 7564 14894 7616 14900
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7392 14090 7420 14350
rect 7576 14346 7604 14894
rect 7668 14346 7696 16934
rect 7564 14340 7616 14346
rect 7564 14282 7616 14288
rect 7656 14340 7708 14346
rect 7656 14282 7708 14288
rect 7392 14074 7512 14090
rect 7392 14068 7524 14074
rect 7392 14062 7472 14068
rect 7472 14010 7524 14016
rect 7760 14006 7788 20810
rect 7932 20596 7984 20602
rect 7932 20538 7984 20544
rect 7840 19440 7892 19446
rect 7840 19382 7892 19388
rect 7852 18970 7880 19382
rect 7840 18964 7892 18970
rect 7840 18906 7892 18912
rect 7944 18442 7972 20538
rect 8128 20534 8156 31758
rect 8312 31754 8340 37198
rect 9048 36786 9076 39200
rect 10336 37126 10364 39200
rect 11624 37262 11652 39200
rect 10416 37256 10468 37262
rect 10416 37198 10468 37204
rect 11612 37256 11664 37262
rect 12268 37244 12296 39200
rect 13556 37262 13584 39200
rect 14844 39114 14872 39200
rect 14936 39114 14964 39222
rect 14844 39086 14964 39114
rect 12440 37256 12492 37262
rect 12268 37216 12440 37244
rect 11612 37198 11664 37204
rect 12440 37198 12492 37204
rect 13544 37256 13596 37262
rect 15120 37244 15148 39222
rect 16118 39200 16174 39800
rect 16762 39200 16818 39800
rect 18050 39200 18106 39800
rect 19338 39200 19394 39800
rect 19982 39200 20038 39800
rect 21270 39200 21326 39800
rect 22558 39200 22614 39800
rect 23202 39200 23258 39800
rect 24490 39200 24546 39800
rect 25778 39200 25834 39800
rect 26422 39200 26478 39800
rect 27710 39200 27766 39800
rect 28998 39200 29054 39800
rect 29642 39200 29698 39800
rect 30930 39200 30986 39800
rect 32218 39200 32274 39800
rect 32862 39200 32918 39800
rect 34150 39200 34206 39800
rect 34256 39222 34468 39250
rect 15200 37256 15252 37262
rect 15120 37216 15200 37244
rect 13544 37198 13596 37204
rect 15200 37198 15252 37204
rect 16028 37256 16080 37262
rect 16028 37198 16080 37204
rect 10324 37120 10376 37126
rect 10324 37062 10376 37068
rect 10428 36922 10456 37198
rect 10508 37188 10560 37194
rect 10508 37130 10560 37136
rect 9956 36916 10008 36922
rect 9956 36858 10008 36864
rect 10416 36916 10468 36922
rect 10416 36858 10468 36864
rect 9036 36780 9088 36786
rect 9036 36722 9088 36728
rect 9772 36576 9824 36582
rect 9772 36518 9824 36524
rect 8312 31726 8432 31754
rect 8208 28552 8260 28558
rect 8208 28494 8260 28500
rect 8220 26314 8248 28494
rect 8208 26308 8260 26314
rect 8208 26250 8260 26256
rect 8300 22432 8352 22438
rect 8300 22374 8352 22380
rect 8208 22160 8260 22166
rect 8208 22102 8260 22108
rect 8220 21418 8248 22102
rect 8312 22030 8340 22374
rect 8300 22024 8352 22030
rect 8300 21966 8352 21972
rect 8404 21434 8432 31726
rect 8484 30728 8536 30734
rect 8484 30670 8536 30676
rect 8496 25974 8524 30670
rect 9784 29646 9812 36518
rect 9968 30734 9996 36858
rect 10520 36786 10548 37130
rect 11704 37120 11756 37126
rect 11704 37062 11756 37068
rect 15016 37120 15068 37126
rect 15016 37062 15068 37068
rect 10508 36780 10560 36786
rect 10508 36722 10560 36728
rect 9956 30728 10008 30734
rect 9956 30670 10008 30676
rect 10232 30592 10284 30598
rect 10232 30534 10284 30540
rect 9772 29640 9824 29646
rect 9772 29582 9824 29588
rect 9220 27872 9272 27878
rect 9220 27814 9272 27820
rect 9232 27674 9260 27814
rect 9220 27668 9272 27674
rect 9220 27610 9272 27616
rect 10048 26988 10100 26994
rect 10048 26930 10100 26936
rect 9404 26920 9456 26926
rect 9404 26862 9456 26868
rect 9416 26586 9444 26862
rect 10060 26586 10088 26930
rect 9404 26580 9456 26586
rect 9404 26522 9456 26528
rect 10048 26580 10100 26586
rect 10048 26522 10100 26528
rect 8484 25968 8536 25974
rect 8484 25910 8536 25916
rect 9956 25900 10008 25906
rect 9956 25842 10008 25848
rect 8668 24812 8720 24818
rect 8668 24754 8720 24760
rect 8576 22500 8628 22506
rect 8576 22442 8628 22448
rect 8588 21690 8616 22442
rect 8576 21684 8628 21690
rect 8576 21626 8628 21632
rect 8208 21412 8260 21418
rect 8208 21354 8260 21360
rect 8312 21406 8432 21434
rect 8116 20528 8168 20534
rect 8116 20470 8168 20476
rect 8208 19712 8260 19718
rect 8208 19654 8260 19660
rect 8116 19508 8168 19514
rect 8116 19450 8168 19456
rect 7944 18414 8064 18442
rect 7932 18352 7984 18358
rect 7932 18294 7984 18300
rect 7944 17338 7972 18294
rect 7932 17332 7984 17338
rect 7932 17274 7984 17280
rect 7840 17196 7892 17202
rect 7840 17138 7892 17144
rect 7852 16697 7880 17138
rect 7838 16688 7894 16697
rect 8036 16674 8064 18414
rect 7838 16623 7894 16632
rect 7944 16646 8064 16674
rect 7840 14476 7892 14482
rect 7840 14418 7892 14424
rect 7852 14385 7880 14418
rect 7838 14376 7894 14385
rect 7838 14311 7894 14320
rect 7380 14000 7432 14006
rect 7748 14000 7800 14006
rect 7432 13948 7604 13954
rect 7380 13942 7604 13948
rect 7748 13942 7800 13948
rect 7392 13926 7604 13942
rect 7380 13864 7432 13870
rect 7380 13806 7432 13812
rect 7392 12918 7420 13806
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 7380 12912 7432 12918
rect 7380 12854 7432 12860
rect 7484 12782 7512 13126
rect 7472 12776 7524 12782
rect 7378 12744 7434 12753
rect 7472 12718 7524 12724
rect 7378 12679 7380 12688
rect 7432 12679 7434 12688
rect 7380 12650 7432 12656
rect 7576 12594 7604 13926
rect 7760 13734 7788 13942
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 7748 13728 7800 13734
rect 7748 13670 7800 13676
rect 7852 13394 7880 13806
rect 7840 13388 7892 13394
rect 7840 13330 7892 13336
rect 7748 12844 7800 12850
rect 7852 12832 7880 13330
rect 7800 12804 7880 12832
rect 7748 12786 7800 12792
rect 7656 12776 7708 12782
rect 7944 12730 7972 16646
rect 8024 16516 8076 16522
rect 8024 16458 8076 16464
rect 8036 16425 8064 16458
rect 8022 16416 8078 16425
rect 8022 16351 8078 16360
rect 8022 15600 8078 15609
rect 8022 15535 8024 15544
rect 8076 15535 8078 15544
rect 8024 15506 8076 15512
rect 8024 15020 8076 15026
rect 8024 14962 8076 14968
rect 7708 12724 7972 12730
rect 7656 12718 7972 12724
rect 7668 12702 7972 12718
rect 7484 12566 7604 12594
rect 7380 11008 7432 11014
rect 7380 10950 7432 10956
rect 7392 10810 7420 10950
rect 7380 10804 7432 10810
rect 7380 10746 7432 10752
rect 7484 10742 7512 12566
rect 7562 12472 7618 12481
rect 7562 12407 7618 12416
rect 7472 10736 7524 10742
rect 7472 10678 7524 10684
rect 7576 8430 7604 12407
rect 7944 10810 7972 12702
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 7930 9208 7986 9217
rect 7840 9172 7892 9178
rect 7892 9152 7930 9160
rect 7892 9143 7986 9152
rect 7892 9132 7972 9143
rect 7840 9114 7892 9120
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7392 7342 7420 8026
rect 7472 7812 7524 7818
rect 7472 7754 7524 7760
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 7484 7002 7512 7754
rect 7576 7002 7604 8366
rect 7656 7744 7708 7750
rect 7656 7686 7708 7692
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7562 6896 7618 6905
rect 7562 6831 7618 6840
rect 7576 6730 7604 6831
rect 7564 6724 7616 6730
rect 7564 6666 7616 6672
rect 7470 5400 7526 5409
rect 7470 5335 7526 5344
rect 7484 5302 7512 5335
rect 7472 5296 7524 5302
rect 7472 5238 7524 5244
rect 7564 5296 7616 5302
rect 7564 5238 7616 5244
rect 7300 4814 7512 4842
rect 7576 4826 7604 5238
rect 7208 4690 7420 4706
rect 7208 4684 7432 4690
rect 7208 4678 7380 4684
rect 7010 4111 7066 4120
rect 7104 4140 7156 4146
rect 7024 4078 7052 4111
rect 7104 4082 7156 4088
rect 7012 4072 7064 4078
rect 7012 4014 7064 4020
rect 6920 3732 6972 3738
rect 7116 3720 7144 4082
rect 6972 3692 7144 3720
rect 6920 3674 6972 3680
rect 6552 3664 6604 3670
rect 6552 3606 6604 3612
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6748 3380 6776 3538
rect 6920 3392 6972 3398
rect 6748 3352 6920 3380
rect 6920 3334 6972 3340
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 6380 2378 6408 3130
rect 7116 2938 7144 3692
rect 7208 3602 7236 4678
rect 7380 4626 7432 4632
rect 7196 3596 7248 3602
rect 7196 3538 7248 3544
rect 7208 3058 7236 3538
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 7024 2910 7144 2938
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 6368 2372 6420 2378
rect 6368 2314 6420 2320
rect 6276 1624 6328 1630
rect 6276 1566 6328 1572
rect 6472 800 6500 2790
rect 7024 2514 7052 2910
rect 7104 2848 7156 2854
rect 7104 2790 7156 2796
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 7116 800 7144 2790
rect 7484 2650 7512 4814
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7668 2854 7696 7686
rect 7760 5914 7788 8774
rect 7840 7472 7892 7478
rect 7838 7440 7840 7449
rect 7892 7440 7894 7449
rect 7838 7375 7894 7384
rect 7944 7342 7972 9132
rect 8036 8294 8064 14962
rect 8128 12481 8156 19450
rect 8220 18970 8248 19654
rect 8208 18964 8260 18970
rect 8208 18906 8260 18912
rect 8312 17202 8340 21406
rect 8392 21344 8444 21350
rect 8392 21286 8444 21292
rect 8404 19446 8432 21286
rect 8680 20874 8708 24754
rect 9864 23520 9916 23526
rect 9864 23462 9916 23468
rect 9772 22976 9824 22982
rect 9772 22918 9824 22924
rect 9784 22710 9812 22918
rect 9876 22710 9904 23462
rect 9772 22704 9824 22710
rect 9772 22646 9824 22652
rect 9864 22704 9916 22710
rect 9864 22646 9916 22652
rect 8852 22228 8904 22234
rect 8852 22170 8904 22176
rect 8760 21684 8812 21690
rect 8760 21626 8812 21632
rect 8668 20868 8720 20874
rect 8668 20810 8720 20816
rect 8484 20800 8536 20806
rect 8484 20742 8536 20748
rect 8496 19786 8524 20742
rect 8484 19780 8536 19786
rect 8484 19722 8536 19728
rect 8576 19780 8628 19786
rect 8576 19722 8628 19728
rect 8588 19530 8616 19722
rect 8496 19502 8616 19530
rect 8392 19440 8444 19446
rect 8392 19382 8444 19388
rect 8496 17513 8524 19502
rect 8576 19440 8628 19446
rect 8576 19382 8628 19388
rect 8588 18222 8616 19382
rect 8668 18828 8720 18834
rect 8668 18770 8720 18776
rect 8680 18290 8708 18770
rect 8772 18426 8800 21626
rect 8864 20602 8892 22170
rect 9036 21956 9088 21962
rect 9036 21898 9088 21904
rect 9048 21078 9076 21898
rect 9968 21486 9996 25842
rect 10048 23724 10100 23730
rect 10048 23666 10100 23672
rect 10060 22234 10088 23666
rect 10244 23186 10272 30534
rect 10520 29170 10548 36722
rect 11716 33522 11744 37062
rect 14464 35692 14516 35698
rect 14464 35634 14516 35640
rect 13912 35080 13964 35086
rect 13912 35022 13964 35028
rect 11704 33516 11756 33522
rect 11704 33458 11756 33464
rect 13924 30326 13952 35022
rect 13912 30320 13964 30326
rect 13912 30262 13964 30268
rect 13452 30252 13504 30258
rect 13452 30194 13504 30200
rect 13084 30048 13136 30054
rect 13084 29990 13136 29996
rect 11428 29504 11480 29510
rect 11428 29446 11480 29452
rect 10508 29164 10560 29170
rect 10508 29106 10560 29112
rect 11336 29028 11388 29034
rect 11336 28970 11388 28976
rect 10324 28552 10376 28558
rect 10324 28494 10376 28500
rect 10336 28218 10364 28494
rect 10324 28212 10376 28218
rect 10324 28154 10376 28160
rect 11152 28076 11204 28082
rect 11152 28018 11204 28024
rect 11164 27606 11192 28018
rect 11152 27600 11204 27606
rect 11152 27542 11204 27548
rect 10968 27396 11020 27402
rect 10968 27338 11020 27344
rect 10980 27062 11008 27338
rect 11152 27328 11204 27334
rect 11152 27270 11204 27276
rect 10968 27056 11020 27062
rect 10968 26998 11020 27004
rect 11060 26784 11112 26790
rect 11060 26726 11112 26732
rect 10692 26580 10744 26586
rect 10692 26522 10744 26528
rect 10704 26382 10732 26522
rect 10508 26376 10560 26382
rect 10508 26318 10560 26324
rect 10692 26376 10744 26382
rect 10692 26318 10744 26324
rect 10520 25906 10548 26318
rect 10784 25968 10836 25974
rect 10784 25910 10836 25916
rect 10508 25900 10560 25906
rect 10508 25842 10560 25848
rect 10520 25809 10548 25842
rect 10506 25800 10562 25809
rect 10506 25735 10562 25744
rect 10796 25498 10824 25910
rect 10784 25492 10836 25498
rect 10784 25434 10836 25440
rect 10692 25288 10744 25294
rect 10692 25230 10744 25236
rect 10704 24818 10732 25230
rect 10692 24812 10744 24818
rect 10692 24754 10744 24760
rect 10324 24608 10376 24614
rect 10324 24550 10376 24556
rect 10232 23180 10284 23186
rect 10232 23122 10284 23128
rect 10140 22432 10192 22438
rect 10140 22374 10192 22380
rect 10048 22228 10100 22234
rect 10048 22170 10100 22176
rect 10152 21962 10180 22374
rect 10140 21956 10192 21962
rect 10140 21898 10192 21904
rect 9956 21480 10008 21486
rect 9956 21422 10008 21428
rect 9404 21412 9456 21418
rect 9404 21354 9456 21360
rect 9036 21072 9088 21078
rect 9036 21014 9088 21020
rect 9312 20936 9364 20942
rect 9312 20878 9364 20884
rect 9220 20800 9272 20806
rect 9220 20742 9272 20748
rect 8852 20596 8904 20602
rect 8852 20538 8904 20544
rect 9232 20534 9260 20742
rect 9220 20528 9272 20534
rect 9220 20470 9272 20476
rect 9220 20392 9272 20398
rect 9220 20334 9272 20340
rect 8944 19848 8996 19854
rect 8944 19790 8996 19796
rect 8760 18420 8812 18426
rect 8760 18362 8812 18368
rect 8668 18284 8720 18290
rect 8668 18226 8720 18232
rect 8576 18216 8628 18222
rect 8576 18158 8628 18164
rect 8680 17678 8708 18226
rect 8668 17672 8720 17678
rect 8668 17614 8720 17620
rect 8482 17504 8538 17513
rect 8482 17439 8538 17448
rect 8300 17196 8352 17202
rect 8300 17138 8352 17144
rect 8312 16538 8340 17138
rect 8496 16538 8524 17439
rect 8576 16992 8628 16998
rect 8576 16934 8628 16940
rect 8588 16726 8616 16934
rect 8576 16720 8628 16726
rect 8576 16662 8628 16668
rect 8220 16510 8340 16538
rect 8404 16510 8524 16538
rect 8220 16182 8248 16510
rect 8208 16176 8260 16182
rect 8208 16118 8260 16124
rect 8298 15600 8354 15609
rect 8298 15535 8354 15544
rect 8312 14006 8340 15535
rect 8404 14958 8432 16510
rect 8484 16448 8536 16454
rect 8484 16390 8536 16396
rect 8496 16182 8524 16390
rect 8484 16176 8536 16182
rect 8484 16118 8536 16124
rect 8576 15904 8628 15910
rect 8576 15846 8628 15852
rect 8484 15632 8536 15638
rect 8482 15600 8484 15609
rect 8536 15600 8538 15609
rect 8482 15535 8538 15544
rect 8496 15502 8524 15535
rect 8484 15496 8536 15502
rect 8484 15438 8536 15444
rect 8392 14952 8444 14958
rect 8392 14894 8444 14900
rect 8392 14544 8444 14550
rect 8484 14544 8536 14550
rect 8392 14486 8444 14492
rect 8482 14512 8484 14521
rect 8536 14512 8538 14521
rect 8300 14000 8352 14006
rect 8300 13942 8352 13948
rect 8208 13728 8260 13734
rect 8208 13670 8260 13676
rect 8220 12730 8248 13670
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8312 13394 8340 13466
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 8220 12702 8340 12730
rect 8208 12640 8260 12646
rect 8208 12582 8260 12588
rect 8114 12472 8170 12481
rect 8114 12407 8170 12416
rect 8220 11830 8248 12582
rect 8208 11824 8260 11830
rect 8208 11766 8260 11772
rect 8312 11642 8340 12702
rect 8220 11614 8340 11642
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 8024 8288 8076 8294
rect 8024 8230 8076 8236
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 8036 6322 8064 7482
rect 8128 6474 8156 10950
rect 8220 9092 8248 11614
rect 8404 9217 8432 14486
rect 8482 14447 8538 14456
rect 8484 13728 8536 13734
rect 8484 13670 8536 13676
rect 8496 13190 8524 13670
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 8588 12646 8616 15846
rect 8576 12640 8628 12646
rect 8576 12582 8628 12588
rect 8680 12434 8708 17614
rect 8852 15564 8904 15570
rect 8852 15506 8904 15512
rect 8760 14272 8812 14278
rect 8760 14214 8812 14220
rect 8772 12986 8800 14214
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 8680 12406 8800 12434
rect 8484 12096 8536 12102
rect 8484 12038 8536 12044
rect 8496 11354 8524 12038
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8668 11280 8720 11286
rect 8574 11248 8630 11257
rect 8668 11222 8720 11228
rect 8574 11183 8630 11192
rect 8588 10538 8616 11183
rect 8576 10532 8628 10538
rect 8576 10474 8628 10480
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8390 9208 8446 9217
rect 8390 9143 8446 9152
rect 8392 9104 8444 9110
rect 8220 9064 8392 9092
rect 8392 9046 8444 9052
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 8496 8362 8524 8910
rect 8588 8430 8616 9998
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8484 8356 8536 8362
rect 8484 8298 8536 8304
rect 8588 7954 8616 8366
rect 8680 8022 8708 11222
rect 8668 8016 8720 8022
rect 8668 7958 8720 7964
rect 8772 7970 8800 12406
rect 8864 9874 8892 15506
rect 8956 11082 8984 19790
rect 9232 19334 9260 20334
rect 9140 19306 9260 19334
rect 9036 18624 9088 18630
rect 9036 18566 9088 18572
rect 9048 12986 9076 18566
rect 9140 15552 9168 19306
rect 9220 18624 9272 18630
rect 9220 18566 9272 18572
rect 9232 16522 9260 18566
rect 9220 16516 9272 16522
rect 9220 16458 9272 16464
rect 9220 16108 9272 16114
rect 9220 16050 9272 16056
rect 9232 15910 9260 16050
rect 9220 15904 9272 15910
rect 9220 15846 9272 15852
rect 9220 15564 9272 15570
rect 9140 15524 9220 15552
rect 9220 15506 9272 15512
rect 9128 14952 9180 14958
rect 9128 14894 9180 14900
rect 9140 14385 9168 14894
rect 9126 14376 9182 14385
rect 9126 14311 9182 14320
rect 9220 14340 9272 14346
rect 9220 14282 9272 14288
rect 9232 13802 9260 14282
rect 9220 13796 9272 13802
rect 9220 13738 9272 13744
rect 9126 13560 9182 13569
rect 9126 13495 9128 13504
rect 9180 13495 9182 13504
rect 9128 13466 9180 13472
rect 9128 13388 9180 13394
rect 9232 13376 9260 13738
rect 9180 13348 9260 13376
rect 9128 13330 9180 13336
rect 9324 13258 9352 20878
rect 9416 19446 9444 21354
rect 9968 21010 9996 21422
rect 9956 21004 10008 21010
rect 9956 20946 10008 20952
rect 10140 20868 10192 20874
rect 10140 20810 10192 20816
rect 9956 20800 10008 20806
rect 9586 20768 9642 20777
rect 9956 20742 10008 20748
rect 9586 20703 9642 20712
rect 9600 20398 9628 20703
rect 9588 20392 9640 20398
rect 9588 20334 9640 20340
rect 9968 20058 9996 20742
rect 9956 20052 10008 20058
rect 9956 19994 10008 20000
rect 9772 19848 9824 19854
rect 9772 19790 9824 19796
rect 9404 19440 9456 19446
rect 9404 19382 9456 19388
rect 9784 18766 9812 19790
rect 10152 19786 10180 20810
rect 10244 20602 10272 23122
rect 10336 23050 10364 24550
rect 11072 24313 11100 26726
rect 11058 24304 11114 24313
rect 11058 24239 11114 24248
rect 10416 23724 10468 23730
rect 10416 23666 10468 23672
rect 10324 23044 10376 23050
rect 10324 22986 10376 22992
rect 10232 20596 10284 20602
rect 10232 20538 10284 20544
rect 10140 19780 10192 19786
rect 10140 19722 10192 19728
rect 10048 19712 10100 19718
rect 10048 19654 10100 19660
rect 10232 19712 10284 19718
rect 10232 19654 10284 19660
rect 9772 18760 9824 18766
rect 9772 18702 9824 18708
rect 9404 18692 9456 18698
rect 9404 18634 9456 18640
rect 9416 15586 9444 18634
rect 9956 18284 10008 18290
rect 9956 18226 10008 18232
rect 9680 18148 9732 18154
rect 9680 18090 9732 18096
rect 9588 18080 9640 18086
rect 9588 18022 9640 18028
rect 9600 17270 9628 18022
rect 9588 17264 9640 17270
rect 9588 17206 9640 17212
rect 9692 17082 9720 18090
rect 9864 17536 9916 17542
rect 9864 17478 9916 17484
rect 9770 17232 9826 17241
rect 9876 17202 9904 17478
rect 9770 17167 9772 17176
rect 9824 17167 9826 17176
rect 9864 17196 9916 17202
rect 9772 17138 9824 17144
rect 9864 17138 9916 17144
rect 9692 17054 9812 17082
rect 9678 16960 9734 16969
rect 9678 16895 9734 16904
rect 9692 16794 9720 16895
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9496 16176 9548 16182
rect 9692 16130 9720 16526
rect 9784 16182 9812 17054
rect 9864 16992 9916 16998
rect 9864 16934 9916 16940
rect 9876 16794 9904 16934
rect 9864 16788 9916 16794
rect 9864 16730 9916 16736
rect 9548 16124 9720 16130
rect 9496 16118 9720 16124
rect 9772 16176 9824 16182
rect 9772 16118 9824 16124
rect 9508 16102 9720 16118
rect 9770 15736 9826 15745
rect 9770 15671 9826 15680
rect 9588 15632 9640 15638
rect 9586 15600 9588 15609
rect 9640 15600 9642 15609
rect 9416 15558 9536 15586
rect 9312 13252 9364 13258
rect 9232 13212 9312 13240
rect 9126 13152 9182 13161
rect 9126 13087 9182 13096
rect 9036 12980 9088 12986
rect 9036 12922 9088 12928
rect 9036 12708 9088 12714
rect 9036 12650 9088 12656
rect 8944 11076 8996 11082
rect 8944 11018 8996 11024
rect 9048 10266 9076 12650
rect 9140 12238 9168 13087
rect 9232 12714 9260 13212
rect 9312 13194 9364 13200
rect 9312 12980 9364 12986
rect 9312 12922 9364 12928
rect 9220 12708 9272 12714
rect 9220 12650 9272 12656
rect 9220 12436 9272 12442
rect 9220 12378 9272 12384
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9232 11626 9260 12378
rect 9220 11620 9272 11626
rect 9220 11562 9272 11568
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 8864 9846 9168 9874
rect 9036 9716 9088 9722
rect 9036 9658 9088 9664
rect 8852 9104 8904 9110
rect 8852 9046 8904 9052
rect 8864 8974 8892 9046
rect 8852 8968 8904 8974
rect 8852 8910 8904 8916
rect 8850 8664 8906 8673
rect 8850 8599 8906 8608
rect 8864 8430 8892 8599
rect 8852 8424 8904 8430
rect 8852 8366 8904 8372
rect 8944 8424 8996 8430
rect 8944 8366 8996 8372
rect 8956 8294 8984 8366
rect 8944 8288 8996 8294
rect 8944 8230 8996 8236
rect 8576 7948 8628 7954
rect 8772 7942 8892 7970
rect 8576 7890 8628 7896
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 8300 7812 8352 7818
rect 8300 7754 8352 7760
rect 8312 7721 8340 7754
rect 8298 7712 8354 7721
rect 8298 7647 8354 7656
rect 8772 7546 8800 7822
rect 8760 7540 8812 7546
rect 8760 7482 8812 7488
rect 8668 6792 8720 6798
rect 8390 6760 8446 6769
rect 8668 6734 8720 6740
rect 8390 6695 8446 6704
rect 8404 6497 8432 6695
rect 8484 6656 8536 6662
rect 8680 6633 8708 6734
rect 8484 6598 8536 6604
rect 8666 6624 8722 6633
rect 8390 6488 8446 6497
rect 8128 6446 8248 6474
rect 8116 6384 8168 6390
rect 8116 6326 8168 6332
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 8128 5914 8156 6326
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 7930 5808 7986 5817
rect 8220 5794 8248 6446
rect 8390 6423 8446 6432
rect 7930 5743 7986 5752
rect 8128 5766 8248 5794
rect 8300 5772 8352 5778
rect 7944 4214 7972 5743
rect 8128 4434 8156 5766
rect 8300 5714 8352 5720
rect 8312 5658 8340 5714
rect 8220 5630 8340 5658
rect 8220 4758 8248 5630
rect 8300 4820 8352 4826
rect 8300 4762 8352 4768
rect 8208 4752 8260 4758
rect 8208 4694 8260 4700
rect 8128 4406 8248 4434
rect 8024 4276 8076 4282
rect 8024 4218 8076 4224
rect 8116 4276 8168 4282
rect 8116 4218 8168 4224
rect 7932 4208 7984 4214
rect 7932 4150 7984 4156
rect 8036 4078 8064 4218
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 8024 4072 8076 4078
rect 8024 4014 8076 4020
rect 7944 3913 7972 4014
rect 7930 3904 7986 3913
rect 7930 3839 7986 3848
rect 8128 3126 8156 4218
rect 8220 3670 8248 4406
rect 8312 4185 8340 4762
rect 8404 4486 8432 6423
rect 8496 6186 8524 6598
rect 8666 6559 8722 6568
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8484 6180 8536 6186
rect 8484 6122 8536 6128
rect 8588 6066 8616 6258
rect 8666 6216 8722 6225
rect 8666 6151 8668 6160
rect 8720 6151 8722 6160
rect 8668 6122 8720 6128
rect 8588 6038 8708 6066
rect 8484 5840 8536 5846
rect 8482 5808 8484 5817
rect 8536 5808 8538 5817
rect 8482 5743 8538 5752
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 8298 4176 8354 4185
rect 8298 4111 8354 4120
rect 8392 4004 8444 4010
rect 8392 3946 8444 3952
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 8404 3505 8432 3946
rect 8390 3496 8446 3505
rect 8390 3431 8446 3440
rect 8574 3360 8630 3369
rect 8574 3295 8630 3304
rect 8588 3126 8616 3295
rect 8116 3120 8168 3126
rect 8116 3062 8168 3068
rect 8576 3120 8628 3126
rect 8576 3062 8628 3068
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 7656 2848 7708 2854
rect 7656 2790 7708 2796
rect 7472 2644 7524 2650
rect 7472 2586 7524 2592
rect 7760 2514 7788 2994
rect 7748 2508 7800 2514
rect 7748 2450 7800 2456
rect 7472 2372 7524 2378
rect 7472 2314 7524 2320
rect 7484 2106 7512 2314
rect 8484 2304 8536 2310
rect 8484 2246 8536 2252
rect 7472 2100 7524 2106
rect 7472 2042 7524 2048
rect 8496 1766 8524 2246
rect 8484 1760 8536 1766
rect 8484 1702 8536 1708
rect 8680 1698 8708 6038
rect 8864 3913 8892 7942
rect 9048 5574 9076 9658
rect 9036 5568 9088 5574
rect 9036 5510 9088 5516
rect 9140 5137 9168 9846
rect 9324 9382 9352 12922
rect 9508 12434 9536 15558
rect 9784 15570 9812 15671
rect 9772 15564 9824 15570
rect 9586 15535 9642 15544
rect 9692 15524 9772 15552
rect 9692 14958 9720 15524
rect 9772 15506 9824 15512
rect 9864 15564 9916 15570
rect 9864 15506 9916 15512
rect 9770 15464 9826 15473
rect 9770 15399 9772 15408
rect 9824 15399 9826 15408
rect 9772 15370 9824 15376
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 9588 14544 9640 14550
rect 9588 14486 9640 14492
rect 9770 14512 9826 14521
rect 9600 13161 9628 14486
rect 9770 14447 9826 14456
rect 9784 14006 9812 14447
rect 9772 14000 9824 14006
rect 9772 13942 9824 13948
rect 9772 13796 9824 13802
rect 9772 13738 9824 13744
rect 9784 13394 9812 13738
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9586 13152 9642 13161
rect 9586 13087 9642 13096
rect 9678 12880 9734 12889
rect 9678 12815 9734 12824
rect 9692 12646 9720 12815
rect 9772 12776 9824 12782
rect 9772 12718 9824 12724
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9784 12481 9812 12718
rect 9416 12406 9536 12434
rect 9770 12472 9826 12481
rect 9876 12442 9904 15506
rect 9770 12407 9826 12416
rect 9864 12436 9916 12442
rect 9312 9376 9364 9382
rect 9312 9318 9364 9324
rect 9416 9042 9444 12406
rect 9864 12378 9916 12384
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 9692 12209 9720 12242
rect 9678 12200 9734 12209
rect 9678 12135 9734 12144
rect 9494 11792 9550 11801
rect 9494 11727 9550 11736
rect 9508 11286 9536 11727
rect 9862 11656 9918 11665
rect 9862 11591 9864 11600
rect 9916 11591 9918 11600
rect 9864 11562 9916 11568
rect 9496 11280 9548 11286
rect 9496 11222 9548 11228
rect 9496 11144 9548 11150
rect 9496 11086 9548 11092
rect 9508 10062 9536 11086
rect 9680 11076 9732 11082
rect 9968 11064 9996 18226
rect 10060 16590 10088 19654
rect 10140 18760 10192 18766
rect 10140 18702 10192 18708
rect 10048 16584 10100 16590
rect 10048 16526 10100 16532
rect 10152 16402 10180 18702
rect 10244 17814 10272 19654
rect 10324 18284 10376 18290
rect 10324 18226 10376 18232
rect 10336 17814 10364 18226
rect 10232 17808 10284 17814
rect 10232 17750 10284 17756
rect 10324 17808 10376 17814
rect 10324 17750 10376 17756
rect 10324 17672 10376 17678
rect 10324 17614 10376 17620
rect 10232 17196 10284 17202
rect 10232 17138 10284 17144
rect 10244 17105 10272 17138
rect 10230 17096 10286 17105
rect 10230 17031 10286 17040
rect 10060 16374 10180 16402
rect 10060 12442 10088 16374
rect 10244 14958 10272 17031
rect 10336 16998 10364 17614
rect 10324 16992 10376 16998
rect 10324 16934 10376 16940
rect 10232 14952 10284 14958
rect 10232 14894 10284 14900
rect 10232 14408 10284 14414
rect 10232 14350 10284 14356
rect 10244 13938 10272 14350
rect 10232 13932 10284 13938
rect 10152 13892 10232 13920
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 9732 11036 9996 11064
rect 9680 11018 9732 11024
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 9508 9654 9536 9998
rect 9586 9752 9642 9761
rect 9586 9687 9588 9696
rect 9640 9687 9642 9696
rect 9588 9658 9640 9664
rect 9496 9648 9548 9654
rect 9496 9590 9548 9596
rect 9494 9072 9550 9081
rect 9404 9036 9456 9042
rect 9494 9007 9496 9016
rect 9404 8978 9456 8984
rect 9548 9007 9550 9016
rect 9496 8978 9548 8984
rect 9586 8936 9642 8945
rect 9312 8900 9364 8906
rect 9312 8842 9364 8848
rect 9404 8900 9456 8906
rect 9586 8871 9642 8880
rect 9404 8842 9456 8848
rect 9324 8566 9352 8842
rect 9312 8560 9364 8566
rect 9312 8502 9364 8508
rect 9312 7336 9364 7342
rect 9416 7313 9444 8842
rect 9600 8838 9628 8871
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9692 7342 9720 11018
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9772 9920 9824 9926
rect 9770 9888 9772 9897
rect 9824 9888 9826 9897
rect 9770 9823 9826 9832
rect 9770 9616 9826 9625
rect 9770 9551 9826 9560
rect 9784 8838 9812 9551
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9680 7336 9732 7342
rect 9312 7278 9364 7284
rect 9402 7304 9458 7313
rect 9220 6384 9272 6390
rect 9324 6372 9352 7278
rect 9680 7278 9732 7284
rect 9402 7239 9458 7248
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9416 6390 9444 6598
rect 9272 6344 9352 6372
rect 9220 6326 9272 6332
rect 9324 5778 9352 6344
rect 9404 6384 9456 6390
rect 9404 6326 9456 6332
rect 9586 6216 9642 6225
rect 9586 6151 9642 6160
rect 9600 6118 9628 6151
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9312 5772 9364 5778
rect 9312 5714 9364 5720
rect 9218 5536 9274 5545
rect 9218 5471 9274 5480
rect 9126 5128 9182 5137
rect 9126 5063 9182 5072
rect 9140 5030 9168 5063
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 9126 4720 9182 4729
rect 9126 4655 9182 4664
rect 9140 4146 9168 4655
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 8850 3904 8906 3913
rect 8850 3839 8906 3848
rect 8760 3460 8812 3466
rect 8760 3402 8812 3408
rect 8668 1692 8720 1698
rect 8668 1634 8720 1640
rect 8404 870 8524 898
rect 8404 800 8432 870
rect 18 200 74 800
rect 662 200 718 800
rect 1950 200 2006 800
rect 3238 200 3294 800
rect 3882 200 3938 800
rect 5170 200 5226 800
rect 6458 200 6514 800
rect 7102 200 7158 800
rect 8390 200 8446 800
rect 8496 762 8524 870
rect 8772 762 8800 3402
rect 8864 2938 8892 3839
rect 9140 3670 9168 4082
rect 9232 4010 9260 5471
rect 9324 5234 9352 5714
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 9496 4752 9548 4758
rect 9496 4694 9548 4700
rect 9508 4321 9536 4694
rect 9588 4684 9640 4690
rect 9588 4626 9640 4632
rect 9494 4312 9550 4321
rect 9494 4247 9550 4256
rect 9220 4004 9272 4010
rect 9220 3946 9272 3952
rect 9494 3768 9550 3777
rect 9494 3703 9496 3712
rect 9548 3703 9550 3712
rect 9496 3674 9548 3680
rect 9128 3664 9180 3670
rect 9128 3606 9180 3612
rect 9600 3534 9628 4626
rect 9680 4004 9732 4010
rect 9680 3946 9732 3952
rect 9588 3528 9640 3534
rect 9402 3496 9458 3505
rect 9588 3470 9640 3476
rect 9402 3431 9404 3440
rect 9456 3431 9458 3440
rect 9404 3402 9456 3408
rect 8864 2922 9168 2938
rect 8864 2916 9180 2922
rect 8864 2910 9128 2916
rect 9128 2858 9180 2864
rect 9692 800 9720 3946
rect 9784 2310 9812 6598
rect 9876 3466 9904 10406
rect 9954 10024 10010 10033
rect 9954 9959 9956 9968
rect 10008 9959 10010 9968
rect 9956 9930 10008 9936
rect 10060 8294 10088 12378
rect 10152 9586 10180 13892
rect 10232 13874 10284 13880
rect 10324 12776 10376 12782
rect 10244 12753 10324 12764
rect 10230 12744 10324 12753
rect 10286 12736 10324 12744
rect 10324 12718 10376 12724
rect 10230 12679 10286 12688
rect 10244 10674 10272 12679
rect 10428 12434 10456 23666
rect 10876 22636 10928 22642
rect 10876 22578 10928 22584
rect 10888 22234 10916 22578
rect 10876 22228 10928 22234
rect 10876 22170 10928 22176
rect 10876 21956 10928 21962
rect 10876 21898 10928 21904
rect 10692 21616 10744 21622
rect 10692 21558 10744 21564
rect 10704 20806 10732 21558
rect 10692 20800 10744 20806
rect 10692 20742 10744 20748
rect 10704 19854 10732 20742
rect 10784 20528 10836 20534
rect 10784 20470 10836 20476
rect 10796 20058 10824 20470
rect 10784 20052 10836 20058
rect 10784 19994 10836 20000
rect 10888 19938 10916 21898
rect 10968 20528 11020 20534
rect 10968 20470 11020 20476
rect 10796 19910 10916 19938
rect 10692 19848 10744 19854
rect 10692 19790 10744 19796
rect 10508 18624 10560 18630
rect 10508 18566 10560 18572
rect 10600 18624 10652 18630
rect 10600 18566 10652 18572
rect 10520 18358 10548 18566
rect 10508 18352 10560 18358
rect 10508 18294 10560 18300
rect 10612 18222 10640 18566
rect 10600 18216 10652 18222
rect 10600 18158 10652 18164
rect 10796 17898 10824 19910
rect 10980 19718 11008 20470
rect 11060 19780 11112 19786
rect 11060 19722 11112 19728
rect 10968 19712 11020 19718
rect 10968 19654 11020 19660
rect 10874 19408 10930 19417
rect 10874 19343 10876 19352
rect 10928 19343 10930 19352
rect 10876 19314 10928 19320
rect 11072 19242 11100 19722
rect 11060 19236 11112 19242
rect 11060 19178 11112 19184
rect 10796 17870 11008 17898
rect 10784 17740 10836 17746
rect 10784 17682 10836 17688
rect 10600 17672 10652 17678
rect 10600 17614 10652 17620
rect 10508 17536 10560 17542
rect 10508 17478 10560 17484
rect 10520 13954 10548 17478
rect 10612 16833 10640 17614
rect 10692 17536 10744 17542
rect 10692 17478 10744 17484
rect 10704 17134 10732 17478
rect 10692 17128 10744 17134
rect 10692 17070 10744 17076
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 10598 16824 10654 16833
rect 10598 16759 10654 16768
rect 10600 16516 10652 16522
rect 10600 16458 10652 16464
rect 10612 15978 10640 16458
rect 10600 15972 10652 15978
rect 10600 15914 10652 15920
rect 10600 15088 10652 15094
rect 10600 15030 10652 15036
rect 10612 14618 10640 15030
rect 10600 14612 10652 14618
rect 10600 14554 10652 14560
rect 10520 13926 10640 13954
rect 10508 13864 10560 13870
rect 10508 13806 10560 13812
rect 10336 12406 10456 12434
rect 10336 11762 10364 12406
rect 10416 12368 10468 12374
rect 10414 12336 10416 12345
rect 10468 12336 10470 12345
rect 10414 12271 10470 12280
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10428 11898 10456 12174
rect 10416 11892 10468 11898
rect 10416 11834 10468 11840
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 10336 10742 10364 11698
rect 10428 11694 10456 11834
rect 10416 11688 10468 11694
rect 10416 11630 10468 11636
rect 10520 10996 10548 13806
rect 10428 10968 10548 10996
rect 10324 10736 10376 10742
rect 10324 10678 10376 10684
rect 10232 10668 10284 10674
rect 10232 10610 10284 10616
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 10232 9988 10284 9994
rect 10232 9930 10284 9936
rect 10244 9897 10272 9930
rect 10230 9888 10286 9897
rect 10230 9823 10286 9832
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 10152 8634 10180 9522
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10152 8362 10180 8570
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 10140 8356 10192 8362
rect 10140 8298 10192 8304
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 10152 6798 10180 8298
rect 10244 7585 10272 8434
rect 10336 8378 10364 10406
rect 10428 9625 10456 10968
rect 10508 10736 10560 10742
rect 10508 10678 10560 10684
rect 10414 9616 10470 9625
rect 10414 9551 10470 9560
rect 10520 8498 10548 10678
rect 10612 10033 10640 13926
rect 10704 12617 10732 16934
rect 10796 16182 10824 17682
rect 10876 17264 10928 17270
rect 10876 17206 10928 17212
rect 10888 17105 10916 17206
rect 10874 17096 10930 17105
rect 10874 17031 10930 17040
rect 10874 16688 10930 16697
rect 10874 16623 10876 16632
rect 10928 16623 10930 16632
rect 10876 16594 10928 16600
rect 10980 16538 11008 17870
rect 11072 17066 11100 19178
rect 11060 17060 11112 17066
rect 11060 17002 11112 17008
rect 10888 16510 11008 16538
rect 10784 16176 10836 16182
rect 10784 16118 10836 16124
rect 10888 15434 10916 16510
rect 10968 16108 11020 16114
rect 10968 16050 11020 16056
rect 10980 15434 11008 16050
rect 10876 15428 10928 15434
rect 10876 15370 10928 15376
rect 10968 15428 11020 15434
rect 10968 15370 11020 15376
rect 10966 15056 11022 15065
rect 10966 14991 11022 15000
rect 10980 14890 11008 14991
rect 10784 14884 10836 14890
rect 10784 14826 10836 14832
rect 10968 14884 11020 14890
rect 10968 14826 11020 14832
rect 10690 12608 10746 12617
rect 10690 12543 10746 12552
rect 10796 12458 10824 14826
rect 10966 14512 11022 14521
rect 10966 14447 11022 14456
rect 10704 12430 10824 12458
rect 10704 11762 10732 12430
rect 10980 12288 11008 14447
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 11072 13870 11100 14350
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 10888 12260 11008 12288
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 10796 11898 10824 12038
rect 10784 11892 10836 11898
rect 10784 11834 10836 11840
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 10704 10742 10732 11698
rect 10888 11370 10916 12260
rect 10968 12164 11020 12170
rect 10968 12106 11020 12112
rect 10980 11558 11008 12106
rect 11072 11762 11100 13806
rect 11060 11756 11112 11762
rect 11060 11698 11112 11704
rect 11164 11694 11192 27270
rect 11348 21010 11376 28970
rect 11336 21004 11388 21010
rect 11336 20946 11388 20952
rect 11336 19984 11388 19990
rect 11336 19926 11388 19932
rect 11244 19304 11296 19310
rect 11244 19246 11296 19252
rect 11256 19009 11284 19246
rect 11242 19000 11298 19009
rect 11242 18935 11298 18944
rect 11244 18760 11296 18766
rect 11244 18702 11296 18708
rect 11256 13802 11284 18702
rect 11348 18465 11376 19926
rect 11440 19174 11468 29446
rect 11520 28416 11572 28422
rect 11520 28358 11572 28364
rect 11532 26994 11560 28358
rect 11980 28076 12032 28082
rect 11980 28018 12032 28024
rect 12992 28076 13044 28082
rect 12992 28018 13044 28024
rect 11612 28008 11664 28014
rect 11612 27950 11664 27956
rect 11520 26988 11572 26994
rect 11520 26930 11572 26936
rect 11624 26382 11652 27950
rect 11888 27872 11940 27878
rect 11888 27814 11940 27820
rect 11900 27538 11928 27814
rect 11888 27532 11940 27538
rect 11888 27474 11940 27480
rect 11992 27334 12020 28018
rect 12072 27940 12124 27946
rect 12072 27882 12124 27888
rect 11980 27328 12032 27334
rect 11980 27270 12032 27276
rect 12084 26994 12112 27882
rect 12716 27872 12768 27878
rect 12716 27814 12768 27820
rect 12728 27538 12756 27814
rect 12532 27532 12584 27538
rect 12532 27474 12584 27480
rect 12716 27532 12768 27538
rect 12716 27474 12768 27480
rect 12440 27464 12492 27470
rect 12440 27406 12492 27412
rect 12452 27130 12480 27406
rect 12440 27124 12492 27130
rect 12440 27066 12492 27072
rect 12256 27056 12308 27062
rect 12256 26998 12308 27004
rect 12072 26988 12124 26994
rect 12072 26930 12124 26936
rect 11796 26920 11848 26926
rect 11796 26862 11848 26868
rect 11612 26376 11664 26382
rect 11612 26318 11664 26324
rect 11624 24818 11652 26318
rect 11808 25838 11836 26862
rect 12072 26376 12124 26382
rect 12072 26318 12124 26324
rect 11796 25832 11848 25838
rect 11796 25774 11848 25780
rect 11808 25430 11836 25774
rect 11796 25424 11848 25430
rect 11796 25366 11848 25372
rect 12084 24818 12112 26318
rect 12164 25696 12216 25702
rect 12164 25638 12216 25644
rect 12176 25294 12204 25638
rect 12164 25288 12216 25294
rect 12164 25230 12216 25236
rect 11612 24812 11664 24818
rect 11612 24754 11664 24760
rect 12072 24812 12124 24818
rect 12072 24754 12124 24760
rect 11888 24336 11940 24342
rect 11888 24278 11940 24284
rect 11520 23520 11572 23526
rect 11520 23462 11572 23468
rect 11532 21962 11560 23462
rect 11900 23118 11928 24278
rect 11888 23112 11940 23118
rect 11888 23054 11940 23060
rect 11612 22568 11664 22574
rect 11612 22510 11664 22516
rect 11624 22098 11652 22510
rect 11704 22500 11756 22506
rect 11704 22442 11756 22448
rect 11612 22092 11664 22098
rect 11612 22034 11664 22040
rect 11520 21956 11572 21962
rect 11520 21898 11572 21904
rect 11624 21842 11652 22034
rect 11532 21814 11652 21842
rect 11532 20398 11560 21814
rect 11612 21548 11664 21554
rect 11612 21490 11664 21496
rect 11520 20392 11572 20398
rect 11520 20334 11572 20340
rect 11428 19168 11480 19174
rect 11428 19110 11480 19116
rect 11334 18456 11390 18465
rect 11334 18391 11390 18400
rect 11336 18284 11388 18290
rect 11336 18226 11388 18232
rect 11348 17649 11376 18226
rect 11440 17746 11468 19110
rect 11532 18222 11560 20334
rect 11624 19854 11652 21490
rect 11612 19848 11664 19854
rect 11612 19790 11664 19796
rect 11624 18272 11652 19790
rect 11716 18766 11744 22442
rect 11796 20392 11848 20398
rect 11796 20334 11848 20340
rect 11808 20058 11836 20334
rect 11796 20052 11848 20058
rect 11796 19994 11848 20000
rect 11796 19168 11848 19174
rect 11796 19110 11848 19116
rect 11808 18766 11836 19110
rect 11900 18986 11928 23054
rect 12268 22094 12296 26998
rect 12544 24274 12572 27474
rect 12900 26920 12952 26926
rect 12900 26862 12952 26868
rect 12808 26852 12860 26858
rect 12808 26794 12860 26800
rect 12624 26580 12676 26586
rect 12624 26522 12676 26528
rect 12636 25498 12664 26522
rect 12820 26450 12848 26794
rect 12808 26444 12860 26450
rect 12808 26386 12860 26392
rect 12912 26246 12940 26862
rect 13004 26314 13032 28018
rect 12992 26308 13044 26314
rect 12992 26250 13044 26256
rect 12900 26240 12952 26246
rect 12900 26182 12952 26188
rect 12624 25492 12676 25498
rect 12624 25434 12676 25440
rect 12900 24812 12952 24818
rect 12900 24754 12952 24760
rect 12716 24744 12768 24750
rect 12716 24686 12768 24692
rect 12624 24608 12676 24614
rect 12624 24550 12676 24556
rect 12532 24268 12584 24274
rect 12532 24210 12584 24216
rect 12636 24138 12664 24550
rect 12624 24132 12676 24138
rect 12624 24074 12676 24080
rect 12348 22976 12400 22982
rect 12348 22918 12400 22924
rect 12176 22066 12296 22094
rect 12070 19272 12126 19281
rect 12176 19258 12204 22066
rect 12256 21004 12308 21010
rect 12256 20946 12308 20952
rect 12268 20602 12296 20946
rect 12360 20874 12388 22918
rect 12440 22704 12492 22710
rect 12440 22646 12492 22652
rect 12348 20868 12400 20874
rect 12348 20810 12400 20816
rect 12256 20596 12308 20602
rect 12256 20538 12308 20544
rect 12452 19938 12480 22646
rect 12532 21956 12584 21962
rect 12532 21898 12584 21904
rect 12544 21418 12572 21898
rect 12532 21412 12584 21418
rect 12532 21354 12584 21360
rect 12624 20868 12676 20874
rect 12624 20810 12676 20816
rect 12360 19910 12480 19938
rect 12256 19780 12308 19786
rect 12360 19768 12388 19910
rect 12532 19780 12584 19786
rect 12308 19740 12388 19768
rect 12452 19740 12532 19768
rect 12256 19722 12308 19728
rect 12176 19230 12388 19258
rect 12070 19207 12072 19216
rect 12124 19207 12126 19216
rect 12072 19178 12124 19184
rect 12256 19168 12308 19174
rect 12256 19110 12308 19116
rect 11900 18958 12204 18986
rect 12072 18828 12124 18834
rect 12072 18770 12124 18776
rect 11704 18760 11756 18766
rect 11702 18728 11704 18737
rect 11796 18760 11848 18766
rect 11756 18728 11758 18737
rect 11796 18702 11848 18708
rect 11702 18663 11758 18672
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 11794 18456 11850 18465
rect 11992 18426 12020 18566
rect 11794 18391 11796 18400
rect 11848 18391 11850 18400
rect 11980 18420 12032 18426
rect 11796 18362 11848 18368
rect 11980 18362 12032 18368
rect 11624 18244 11928 18272
rect 11520 18216 11572 18222
rect 11520 18158 11572 18164
rect 11702 18184 11758 18193
rect 11702 18119 11758 18128
rect 11428 17740 11480 17746
rect 11428 17682 11480 17688
rect 11334 17640 11390 17649
rect 11520 17604 11572 17610
rect 11334 17575 11390 17584
rect 11440 17564 11520 17592
rect 11440 17202 11468 17564
rect 11520 17546 11572 17552
rect 11520 17332 11572 17338
rect 11520 17274 11572 17280
rect 11612 17332 11664 17338
rect 11612 17274 11664 17280
rect 11428 17196 11480 17202
rect 11428 17138 11480 17144
rect 11440 16590 11468 17138
rect 11532 16658 11560 17274
rect 11624 16969 11652 17274
rect 11610 16960 11666 16969
rect 11610 16895 11666 16904
rect 11520 16652 11572 16658
rect 11520 16594 11572 16600
rect 11428 16584 11480 16590
rect 11428 16526 11480 16532
rect 11612 16584 11664 16590
rect 11612 16526 11664 16532
rect 11624 15026 11652 16526
rect 11612 15020 11664 15026
rect 11612 14962 11664 14968
rect 11336 14952 11388 14958
rect 11336 14894 11388 14900
rect 11348 14346 11376 14894
rect 11336 14340 11388 14346
rect 11336 14282 11388 14288
rect 11244 13796 11296 13802
rect 11244 13738 11296 13744
rect 11244 12300 11296 12306
rect 11244 12242 11296 12248
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 10968 11552 11020 11558
rect 10968 11494 11020 11500
rect 10888 11342 11008 11370
rect 11164 11354 11192 11630
rect 11256 11558 11284 12242
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 10784 11212 10836 11218
rect 10784 11154 10836 11160
rect 10796 10849 10824 11154
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 10782 10840 10838 10849
rect 10888 10810 10916 11086
rect 10782 10775 10838 10784
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10692 10736 10744 10742
rect 10692 10678 10744 10684
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 10598 10024 10654 10033
rect 10598 9959 10654 9968
rect 10612 9178 10640 9959
rect 10600 9172 10652 9178
rect 10600 9114 10652 9120
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10336 8350 10456 8378
rect 10230 7576 10286 7585
rect 10230 7511 10286 7520
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 9956 6452 10008 6458
rect 10152 6440 10180 6734
rect 10008 6412 10180 6440
rect 10322 6488 10378 6497
rect 10322 6423 10378 6432
rect 9956 6394 10008 6400
rect 9956 6180 10008 6186
rect 9956 6122 10008 6128
rect 9968 6089 9996 6122
rect 9954 6080 10010 6089
rect 9954 6015 10010 6024
rect 9956 5296 10008 5302
rect 9956 5238 10008 5244
rect 9968 4826 9996 5238
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 10060 4486 10088 5102
rect 10048 4480 10100 4486
rect 9954 4448 10010 4457
rect 10048 4422 10100 4428
rect 9954 4383 10010 4392
rect 9968 3670 9996 4383
rect 10152 4214 10180 6412
rect 10336 6390 10364 6423
rect 10324 6384 10376 6390
rect 10324 6326 10376 6332
rect 10230 6216 10286 6225
rect 10230 6151 10286 6160
rect 10140 4208 10192 4214
rect 10140 4150 10192 4156
rect 10048 4072 10100 4078
rect 10048 4014 10100 4020
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 10060 3534 10088 4014
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 9864 3460 9916 3466
rect 9864 3402 9916 3408
rect 10244 3058 10272 6151
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 10428 2774 10456 8350
rect 10600 8288 10652 8294
rect 10600 8230 10652 8236
rect 10612 8022 10640 8230
rect 10600 8016 10652 8022
rect 10600 7958 10652 7964
rect 10796 6322 10824 10610
rect 10980 9602 11008 11342
rect 11152 11348 11204 11354
rect 11152 11290 11204 11296
rect 11348 10266 11376 14282
rect 11518 13968 11574 13977
rect 11518 13903 11574 13912
rect 11428 12708 11480 12714
rect 11428 12650 11480 12656
rect 11440 12617 11468 12650
rect 11426 12608 11482 12617
rect 11426 12543 11482 12552
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11440 12345 11468 12378
rect 11426 12336 11482 12345
rect 11426 12271 11482 12280
rect 11532 12220 11560 13903
rect 11624 12986 11652 14962
rect 11716 14958 11744 18119
rect 11796 17128 11848 17134
rect 11796 17070 11848 17076
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11808 13977 11836 17070
rect 11900 15450 11928 18244
rect 12084 18222 12112 18770
rect 12072 18216 12124 18222
rect 12072 18158 12124 18164
rect 11980 17808 12032 17814
rect 11980 17750 12032 17756
rect 11992 15609 12020 17750
rect 12072 16652 12124 16658
rect 12072 16594 12124 16600
rect 11978 15600 12034 15609
rect 11978 15535 12034 15544
rect 11900 15422 12020 15450
rect 11888 15360 11940 15366
rect 11888 15302 11940 15308
rect 11900 14929 11928 15302
rect 11886 14920 11942 14929
rect 11886 14855 11942 14864
rect 11794 13968 11850 13977
rect 11794 13903 11850 13912
rect 11888 13932 11940 13938
rect 11888 13874 11940 13880
rect 11900 13841 11928 13874
rect 11886 13832 11942 13841
rect 11886 13767 11942 13776
rect 11992 13546 12020 15422
rect 11716 13518 12020 13546
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11716 12866 11744 13518
rect 11888 13320 11940 13326
rect 11940 13280 12020 13308
rect 11888 13262 11940 13268
rect 11992 12986 12020 13280
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 11440 12192 11560 12220
rect 11624 12838 11744 12866
rect 11992 12850 12020 12922
rect 11980 12844 12032 12850
rect 11440 10606 11468 12192
rect 11518 11928 11574 11937
rect 11518 11863 11574 11872
rect 11532 11830 11560 11863
rect 11520 11824 11572 11830
rect 11520 11766 11572 11772
rect 11520 11008 11572 11014
rect 11520 10950 11572 10956
rect 11428 10600 11480 10606
rect 11428 10542 11480 10548
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 11532 10198 11560 10950
rect 11520 10192 11572 10198
rect 11520 10134 11572 10140
rect 10980 9574 11100 9602
rect 10876 8832 10928 8838
rect 10876 8774 10928 8780
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 10598 5536 10654 5545
rect 10598 5471 10654 5480
rect 10506 5264 10562 5273
rect 10506 5199 10562 5208
rect 10520 4826 10548 5199
rect 10508 4820 10560 4826
rect 10508 4762 10560 4768
rect 10520 3058 10548 4762
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 10612 2990 10640 5471
rect 10690 3768 10746 3777
rect 10690 3703 10692 3712
rect 10744 3703 10746 3712
rect 10692 3674 10744 3680
rect 10888 3058 10916 8774
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10980 7886 11008 8434
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 10980 7002 11008 7142
rect 10968 6996 11020 7002
rect 10968 6938 11020 6944
rect 11072 4078 11100 9574
rect 11244 9036 11296 9042
rect 11244 8978 11296 8984
rect 11150 6896 11206 6905
rect 11150 6831 11206 6840
rect 11164 5681 11192 6831
rect 11150 5672 11206 5681
rect 11150 5607 11206 5616
rect 11152 5568 11204 5574
rect 11152 5510 11204 5516
rect 11164 5166 11192 5510
rect 11152 5160 11204 5166
rect 11152 5102 11204 5108
rect 11164 4690 11192 5102
rect 11152 4684 11204 4690
rect 11152 4626 11204 4632
rect 11060 4072 11112 4078
rect 11060 4014 11112 4020
rect 11152 3120 11204 3126
rect 11152 3062 11204 3068
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 11164 2990 11192 3062
rect 10600 2984 10652 2990
rect 10600 2926 10652 2932
rect 11152 2984 11204 2990
rect 11152 2926 11204 2932
rect 10336 2746 10456 2774
rect 11256 2774 11284 8978
rect 11624 7426 11652 12838
rect 11980 12786 12032 12792
rect 11704 12776 11756 12782
rect 11704 12718 11756 12724
rect 11716 11218 11744 12718
rect 12084 12356 12112 16594
rect 12176 13394 12204 18958
rect 12268 17270 12296 19110
rect 12360 17377 12388 19230
rect 12452 18426 12480 19740
rect 12532 19722 12584 19728
rect 12532 19440 12584 19446
rect 12636 19417 12664 20810
rect 12532 19382 12584 19388
rect 12622 19408 12678 19417
rect 12544 18698 12572 19382
rect 12622 19343 12678 19352
rect 12622 19272 12678 19281
rect 12622 19207 12678 19216
rect 12636 18902 12664 19207
rect 12624 18896 12676 18902
rect 12624 18838 12676 18844
rect 12532 18692 12584 18698
rect 12532 18634 12584 18640
rect 12440 18420 12492 18426
rect 12440 18362 12492 18368
rect 12346 17368 12402 17377
rect 12346 17303 12402 17312
rect 12256 17264 12308 17270
rect 12256 17206 12308 17212
rect 12254 17096 12310 17105
rect 12254 17031 12310 17040
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 11979 12328 12112 12356
rect 11979 12288 12007 12328
rect 12268 12306 12296 17031
rect 12360 16046 12388 17303
rect 12728 17252 12756 24686
rect 12912 24274 12940 24754
rect 13096 24750 13124 29990
rect 13268 27872 13320 27878
rect 13268 27814 13320 27820
rect 13176 25900 13228 25906
rect 13176 25842 13228 25848
rect 13084 24744 13136 24750
rect 13084 24686 13136 24692
rect 12900 24268 12952 24274
rect 12900 24210 12952 24216
rect 12992 23792 13044 23798
rect 12992 23734 13044 23740
rect 13004 22778 13032 23734
rect 13096 23662 13124 24686
rect 13084 23656 13136 23662
rect 13084 23598 13136 23604
rect 12992 22772 13044 22778
rect 12992 22714 13044 22720
rect 13188 22094 13216 25842
rect 13280 25362 13308 27814
rect 13464 27606 13492 30194
rect 13452 27600 13504 27606
rect 13452 27542 13504 27548
rect 13464 27130 13492 27542
rect 13452 27124 13504 27130
rect 13452 27066 13504 27072
rect 14004 26988 14056 26994
rect 14004 26930 14056 26936
rect 13452 26240 13504 26246
rect 13452 26182 13504 26188
rect 13464 25498 13492 26182
rect 14016 26042 14044 26930
rect 14188 26376 14240 26382
rect 14188 26318 14240 26324
rect 14004 26036 14056 26042
rect 14004 25978 14056 25984
rect 14200 25906 14228 26318
rect 14188 25900 14240 25906
rect 14188 25842 14240 25848
rect 13452 25492 13504 25498
rect 13452 25434 13504 25440
rect 13268 25356 13320 25362
rect 13268 25298 13320 25304
rect 14372 25152 14424 25158
rect 14372 25094 14424 25100
rect 14384 24886 14412 25094
rect 14372 24880 14424 24886
rect 14372 24822 14424 24828
rect 13360 24744 13412 24750
rect 13360 24686 13412 24692
rect 13268 24268 13320 24274
rect 13268 24210 13320 24216
rect 13096 22066 13216 22094
rect 13280 22094 13308 24210
rect 13372 23186 13400 24686
rect 13728 24132 13780 24138
rect 13728 24074 13780 24080
rect 13452 23588 13504 23594
rect 13452 23530 13504 23536
rect 13464 23186 13492 23530
rect 13360 23180 13412 23186
rect 13360 23122 13412 23128
rect 13452 23180 13504 23186
rect 13452 23122 13504 23128
rect 13360 22704 13412 22710
rect 13464 22658 13492 23122
rect 13412 22652 13492 22658
rect 13360 22646 13492 22652
rect 13372 22630 13492 22646
rect 13740 22574 13768 24074
rect 14188 23588 14240 23594
rect 14188 23530 14240 23536
rect 13912 23112 13964 23118
rect 13912 23054 13964 23060
rect 13728 22568 13780 22574
rect 13728 22510 13780 22516
rect 13740 22166 13768 22510
rect 13728 22160 13780 22166
rect 13728 22102 13780 22108
rect 13280 22066 13400 22094
rect 12992 21888 13044 21894
rect 12992 21830 13044 21836
rect 12808 21616 12860 21622
rect 12808 21558 12860 21564
rect 12820 18086 12848 21558
rect 13004 21049 13032 21830
rect 12990 21040 13046 21049
rect 12990 20975 13046 20984
rect 12900 19712 12952 19718
rect 12900 19654 12952 19660
rect 12808 18080 12860 18086
rect 12808 18022 12860 18028
rect 12452 17224 12756 17252
rect 12348 16040 12400 16046
rect 12348 15982 12400 15988
rect 12348 15632 12400 15638
rect 12348 15574 12400 15580
rect 12360 15473 12388 15574
rect 12346 15464 12402 15473
rect 12346 15399 12402 15408
rect 12348 14476 12400 14482
rect 12348 14418 12400 14424
rect 12360 13977 12388 14418
rect 12346 13968 12402 13977
rect 12346 13903 12402 13912
rect 12348 13728 12400 13734
rect 12348 13670 12400 13676
rect 12256 12300 12308 12306
rect 11979 12260 12112 12288
rect 11888 11824 11940 11830
rect 11808 11801 11888 11812
rect 11794 11792 11888 11801
rect 11850 11784 11888 11792
rect 11888 11766 11940 11772
rect 11794 11727 11850 11736
rect 11704 11212 11756 11218
rect 11704 11154 11756 11160
rect 11980 11076 12032 11082
rect 11980 11018 12032 11024
rect 11992 10674 12020 11018
rect 11980 10668 12032 10674
rect 11980 10610 12032 10616
rect 11704 10600 11756 10606
rect 12084 10554 12112 12260
rect 12256 12242 12308 12248
rect 11704 10542 11756 10548
rect 11716 10266 11744 10542
rect 11992 10526 12112 10554
rect 11704 10260 11756 10266
rect 11704 10202 11756 10208
rect 11888 10056 11940 10062
rect 11888 9998 11940 10004
rect 11900 9518 11928 9998
rect 11888 9512 11940 9518
rect 11888 9454 11940 9460
rect 11532 7398 11652 7426
rect 11532 6254 11560 7398
rect 11612 7336 11664 7342
rect 11612 7278 11664 7284
rect 11520 6248 11572 6254
rect 11520 6190 11572 6196
rect 11334 6080 11390 6089
rect 11334 6015 11390 6024
rect 11348 5846 11376 6015
rect 11336 5840 11388 5846
rect 11336 5782 11388 5788
rect 11348 4010 11376 5782
rect 11624 5624 11652 7278
rect 11886 7032 11942 7041
rect 11886 6967 11942 6976
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11716 6254 11744 6734
rect 11704 6248 11756 6254
rect 11704 6190 11756 6196
rect 11716 5692 11744 6190
rect 11796 5704 11848 5710
rect 11716 5664 11796 5692
rect 11796 5646 11848 5652
rect 11624 5596 11744 5624
rect 11716 5166 11744 5596
rect 11704 5160 11756 5166
rect 11704 5102 11756 5108
rect 11716 4146 11744 5102
rect 11808 4690 11836 5646
rect 11796 4684 11848 4690
rect 11796 4626 11848 4632
rect 11796 4548 11848 4554
rect 11796 4490 11848 4496
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 11336 4004 11388 4010
rect 11336 3946 11388 3952
rect 11808 2774 11836 4490
rect 11900 3738 11928 6967
rect 11992 6730 12020 10526
rect 12268 9674 12296 12242
rect 12360 10810 12388 13670
rect 12452 12434 12480 17224
rect 12912 16522 12940 19654
rect 13004 19310 13032 20975
rect 13096 19530 13124 22066
rect 13176 21888 13228 21894
rect 13176 21830 13228 21836
rect 13188 21486 13216 21830
rect 13176 21480 13228 21486
rect 13176 21422 13228 21428
rect 13174 21312 13230 21321
rect 13174 21247 13230 21256
rect 13188 20398 13216 21247
rect 13268 21004 13320 21010
rect 13268 20946 13320 20952
rect 13280 20777 13308 20946
rect 13266 20768 13322 20777
rect 13266 20703 13322 20712
rect 13268 20528 13320 20534
rect 13268 20470 13320 20476
rect 13176 20392 13228 20398
rect 13176 20334 13228 20340
rect 13096 19502 13216 19530
rect 13280 19514 13308 20470
rect 13084 19440 13136 19446
rect 13084 19382 13136 19388
rect 12992 19304 13044 19310
rect 12992 19246 13044 19252
rect 12990 19136 13046 19145
rect 12990 19071 13046 19080
rect 13004 18850 13032 19071
rect 13096 18970 13124 19382
rect 13188 19334 13216 19502
rect 13268 19508 13320 19514
rect 13268 19450 13320 19456
rect 13188 19306 13308 19334
rect 13084 18964 13136 18970
rect 13084 18906 13136 18912
rect 13004 18822 13124 18850
rect 12992 17604 13044 17610
rect 12992 17546 13044 17552
rect 12624 16516 12676 16522
rect 12624 16458 12676 16464
rect 12900 16516 12952 16522
rect 12900 16458 12952 16464
rect 12636 15706 12664 16458
rect 12808 16040 12860 16046
rect 12808 15982 12860 15988
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 12624 15700 12676 15706
rect 12624 15642 12676 15648
rect 12544 15586 12572 15642
rect 12544 15558 12756 15586
rect 12532 15088 12584 15094
rect 12530 15056 12532 15065
rect 12584 15056 12586 15065
rect 12530 14991 12586 15000
rect 12624 14952 12676 14958
rect 12624 14894 12676 14900
rect 12636 14414 12664 14894
rect 12624 14408 12676 14414
rect 12624 14350 12676 14356
rect 12532 13524 12584 13530
rect 12532 13466 12584 13472
rect 12544 13433 12572 13466
rect 12530 13424 12586 13433
rect 12728 13394 12756 15558
rect 12820 15337 12848 15982
rect 13004 15473 13032 17546
rect 12990 15464 13046 15473
rect 12912 15422 12990 15450
rect 12806 15328 12862 15337
rect 12806 15263 12862 15272
rect 12530 13359 12586 13368
rect 12716 13388 12768 13394
rect 12716 13330 12768 13336
rect 12806 12744 12862 12753
rect 12806 12679 12862 12688
rect 12452 12406 12572 12434
rect 12544 12209 12572 12406
rect 12716 12300 12768 12306
rect 12716 12242 12768 12248
rect 12530 12200 12586 12209
rect 12530 12135 12586 12144
rect 12440 11824 12492 11830
rect 12440 11766 12492 11772
rect 12452 11665 12480 11766
rect 12438 11656 12494 11665
rect 12438 11591 12494 11600
rect 12544 11218 12572 12135
rect 12728 12102 12756 12242
rect 12820 12238 12848 12679
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12912 11529 12940 15422
rect 12990 15399 13046 15408
rect 13096 15366 13124 18822
rect 13176 18216 13228 18222
rect 13176 18158 13228 18164
rect 13084 15360 13136 15366
rect 13084 15302 13136 15308
rect 13082 15192 13138 15201
rect 13082 15127 13138 15136
rect 13096 15094 13124 15127
rect 13084 15088 13136 15094
rect 13084 15030 13136 15036
rect 13084 14272 13136 14278
rect 13084 14214 13136 14220
rect 13096 14006 13124 14214
rect 13084 14000 13136 14006
rect 13084 13942 13136 13948
rect 13188 13818 13216 18158
rect 13096 13790 13216 13818
rect 12990 13696 13046 13705
rect 12990 13631 13046 13640
rect 12898 11520 12954 11529
rect 12898 11455 12954 11464
rect 13004 11370 13032 13631
rect 12820 11342 13032 11370
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 12438 10976 12494 10985
rect 12438 10911 12494 10920
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 12084 9646 12296 9674
rect 12084 7002 12112 9646
rect 12452 9602 12480 10911
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 12532 10668 12584 10674
rect 12532 10610 12584 10616
rect 12544 9722 12572 10610
rect 12636 9994 12664 10746
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12624 9988 12676 9994
rect 12624 9930 12676 9936
rect 12532 9716 12584 9722
rect 12532 9658 12584 9664
rect 12268 9586 12480 9602
rect 12256 9580 12480 9586
rect 12308 9574 12480 9580
rect 12256 9522 12308 9528
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12254 9072 12310 9081
rect 12360 9042 12388 9454
rect 12254 9007 12310 9016
rect 12348 9036 12400 9042
rect 12268 8498 12296 9007
rect 12348 8978 12400 8984
rect 12452 8809 12480 9574
rect 12728 8974 12756 10406
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 12438 8800 12494 8809
rect 12438 8735 12494 8744
rect 12348 8560 12400 8566
rect 12346 8528 12348 8537
rect 12400 8528 12402 8537
rect 12256 8492 12308 8498
rect 12346 8463 12402 8472
rect 12256 8434 12308 8440
rect 12440 8424 12492 8430
rect 12440 8366 12492 8372
rect 12164 7336 12216 7342
rect 12164 7278 12216 7284
rect 12176 7177 12204 7278
rect 12162 7168 12218 7177
rect 12162 7103 12218 7112
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 12164 6996 12216 7002
rect 12164 6938 12216 6944
rect 12176 6905 12204 6938
rect 12162 6896 12218 6905
rect 12072 6860 12124 6866
rect 12162 6831 12218 6840
rect 12348 6860 12400 6866
rect 12072 6802 12124 6808
rect 12348 6802 12400 6808
rect 12084 6769 12112 6802
rect 12070 6760 12126 6769
rect 11980 6724 12032 6730
rect 12070 6695 12126 6704
rect 11980 6666 12032 6672
rect 11992 5846 12020 6666
rect 12072 6656 12124 6662
rect 12360 6610 12388 6802
rect 12452 6730 12480 8366
rect 12440 6724 12492 6730
rect 12440 6666 12492 6672
rect 12124 6604 12388 6610
rect 12072 6598 12388 6604
rect 12084 6582 12388 6598
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 12440 6384 12492 6390
rect 12440 6326 12492 6332
rect 12254 5944 12310 5953
rect 12254 5879 12310 5888
rect 11980 5840 12032 5846
rect 11980 5782 12032 5788
rect 12268 5658 12296 5879
rect 12346 5672 12402 5681
rect 12268 5630 12346 5658
rect 12346 5607 12402 5616
rect 12070 4992 12126 5001
rect 12070 4927 12126 4936
rect 12084 4554 12112 4927
rect 12072 4548 12124 4554
rect 12072 4490 12124 4496
rect 12256 4480 12308 4486
rect 12256 4422 12308 4428
rect 12268 4282 12296 4422
rect 12256 4276 12308 4282
rect 12256 4218 12308 4224
rect 12452 4026 12480 6326
rect 12728 5642 12756 6394
rect 12716 5636 12768 5642
rect 12716 5578 12768 5584
rect 12820 5409 12848 11342
rect 12992 11280 13044 11286
rect 12992 11222 13044 11228
rect 12900 9036 12952 9042
rect 12900 8978 12952 8984
rect 12912 8498 12940 8978
rect 13004 8838 13032 11222
rect 13096 9874 13124 13790
rect 13280 13716 13308 19306
rect 13188 13688 13308 13716
rect 13188 12481 13216 13688
rect 13174 12472 13230 12481
rect 13174 12407 13230 12416
rect 13268 12436 13320 12442
rect 13268 12378 13320 12384
rect 13096 9846 13216 9874
rect 13084 9648 13136 9654
rect 13082 9616 13084 9625
rect 13136 9616 13138 9625
rect 13082 9551 13138 9560
rect 13188 8838 13216 9846
rect 12992 8832 13044 8838
rect 12992 8774 13044 8780
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 13188 8566 13216 8774
rect 13176 8560 13228 8566
rect 13176 8502 13228 8508
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 12900 8356 12952 8362
rect 12900 8298 12952 8304
rect 12912 7886 12940 8298
rect 12900 7880 12952 7886
rect 12900 7822 12952 7828
rect 13176 7540 13228 7546
rect 13176 7482 13228 7488
rect 13188 6118 13216 7482
rect 13280 6934 13308 12378
rect 13372 11558 13400 22066
rect 13452 21480 13504 21486
rect 13452 21422 13504 21428
rect 13464 20398 13492 21422
rect 13728 21412 13780 21418
rect 13728 21354 13780 21360
rect 13544 21072 13596 21078
rect 13544 21014 13596 21020
rect 13452 20392 13504 20398
rect 13452 20334 13504 20340
rect 13452 19780 13504 19786
rect 13452 19722 13504 19728
rect 13464 19446 13492 19722
rect 13556 19718 13584 21014
rect 13740 20942 13768 21354
rect 13728 20936 13780 20942
rect 13728 20878 13780 20884
rect 13820 20392 13872 20398
rect 13820 20334 13872 20340
rect 13544 19712 13596 19718
rect 13544 19654 13596 19660
rect 13452 19440 13504 19446
rect 13452 19382 13504 19388
rect 13464 18426 13492 19382
rect 13452 18420 13504 18426
rect 13452 18362 13504 18368
rect 13556 17218 13584 19654
rect 13728 18828 13780 18834
rect 13728 18770 13780 18776
rect 13740 18222 13768 18770
rect 13728 18216 13780 18222
rect 13728 18158 13780 18164
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 13740 17377 13768 17818
rect 13832 17678 13860 20334
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 13726 17368 13782 17377
rect 13726 17303 13782 17312
rect 13556 17190 13676 17218
rect 13544 17128 13596 17134
rect 13544 17070 13596 17076
rect 13452 16992 13504 16998
rect 13452 16934 13504 16940
rect 13464 16182 13492 16934
rect 13452 16176 13504 16182
rect 13452 16118 13504 16124
rect 13452 16040 13504 16046
rect 13450 16008 13452 16017
rect 13504 16008 13506 16017
rect 13450 15943 13506 15952
rect 13556 15910 13584 17070
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13452 15360 13504 15366
rect 13452 15302 13504 15308
rect 13464 11801 13492 15302
rect 13556 15201 13584 15846
rect 13542 15192 13598 15201
rect 13542 15127 13598 15136
rect 13648 15042 13676 17190
rect 13728 16040 13780 16046
rect 13728 15982 13780 15988
rect 13556 15014 13676 15042
rect 13556 13308 13584 15014
rect 13634 13696 13690 13705
rect 13634 13631 13690 13640
rect 13648 13462 13676 13631
rect 13636 13456 13688 13462
rect 13636 13398 13688 13404
rect 13740 13394 13768 15982
rect 13924 15570 13952 23054
rect 14004 22024 14056 22030
rect 14004 21966 14056 21972
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 13912 15564 13964 15570
rect 13912 15506 13964 15512
rect 13832 15473 13860 15506
rect 13818 15464 13874 15473
rect 14016 15450 14044 21966
rect 14096 20596 14148 20602
rect 14096 20538 14148 20544
rect 14108 19922 14136 20538
rect 14200 20210 14228 23530
rect 14372 22704 14424 22710
rect 14372 22646 14424 22652
rect 14384 22098 14412 22646
rect 14372 22092 14424 22098
rect 14372 22034 14424 22040
rect 14372 21344 14424 21350
rect 14372 21286 14424 21292
rect 14384 21185 14412 21286
rect 14370 21176 14426 21185
rect 14370 21111 14426 21120
rect 14280 20460 14332 20466
rect 14280 20402 14332 20408
rect 14292 20369 14320 20402
rect 14278 20360 14334 20369
rect 14278 20295 14334 20304
rect 14200 20182 14320 20210
rect 14096 19916 14148 19922
rect 14096 19858 14148 19864
rect 14188 18284 14240 18290
rect 14188 18226 14240 18232
rect 14096 17740 14148 17746
rect 14096 17682 14148 17688
rect 14108 16998 14136 17682
rect 14096 16992 14148 16998
rect 14096 16934 14148 16940
rect 14096 16516 14148 16522
rect 14096 16458 14148 16464
rect 14108 16153 14136 16458
rect 14094 16144 14150 16153
rect 14094 16079 14150 16088
rect 14094 15600 14150 15609
rect 14094 15535 14150 15544
rect 13818 15399 13874 15408
rect 13924 15422 14044 15450
rect 13818 14920 13874 14929
rect 13818 14855 13874 14864
rect 13832 14006 13860 14855
rect 13820 14000 13872 14006
rect 13820 13942 13872 13948
rect 13728 13388 13780 13394
rect 13728 13330 13780 13336
rect 13556 13280 13676 13308
rect 13450 11792 13506 11801
rect 13450 11727 13506 11736
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13372 11286 13400 11494
rect 13360 11280 13412 11286
rect 13360 11222 13412 11228
rect 13360 11076 13412 11082
rect 13360 11018 13412 11024
rect 13372 10674 13400 11018
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13372 7886 13400 8570
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13268 6928 13320 6934
rect 13268 6870 13320 6876
rect 13176 6112 13228 6118
rect 13176 6054 13228 6060
rect 12806 5400 12862 5409
rect 12806 5335 12862 5344
rect 13266 4992 13322 5001
rect 13266 4927 13322 4936
rect 12990 4856 13046 4865
rect 12990 4791 13046 4800
rect 12530 4312 12586 4321
rect 12530 4247 12586 4256
rect 12624 4276 12676 4282
rect 12544 4214 12572 4247
rect 12624 4218 12676 4224
rect 12532 4208 12584 4214
rect 12532 4150 12584 4156
rect 12636 4078 12664 4218
rect 12360 3998 12480 4026
rect 12624 4072 12676 4078
rect 12624 4014 12676 4020
rect 11888 3732 11940 3738
rect 11888 3674 11940 3680
rect 12360 3398 12388 3998
rect 12900 3732 12952 3738
rect 12900 3674 12952 3680
rect 12532 3596 12584 3602
rect 12532 3538 12584 3544
rect 12544 3482 12572 3538
rect 12544 3466 12664 3482
rect 12544 3460 12676 3466
rect 12544 3454 12624 3460
rect 12624 3402 12676 3408
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 12622 3360 12678 3369
rect 12622 3295 12678 3304
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 11900 3097 11928 3130
rect 11886 3088 11942 3097
rect 11886 3023 11942 3032
rect 11978 2952 12034 2961
rect 11978 2887 11980 2896
rect 12032 2887 12034 2896
rect 11980 2858 12032 2864
rect 12636 2825 12664 3295
rect 12912 3058 12940 3674
rect 12900 3052 12952 3058
rect 12900 2994 12952 3000
rect 11256 2746 11652 2774
rect 9772 2304 9824 2310
rect 9772 2246 9824 2252
rect 10336 800 10364 2746
rect 11152 2304 11204 2310
rect 11058 2272 11114 2281
rect 11152 2246 11204 2252
rect 11058 2207 11114 2216
rect 11072 1834 11100 2207
rect 11164 1970 11192 2246
rect 11152 1964 11204 1970
rect 11152 1906 11204 1912
rect 11060 1828 11112 1834
rect 11060 1770 11112 1776
rect 11624 800 11652 2746
rect 11716 2746 11836 2774
rect 12622 2816 12678 2825
rect 12622 2751 12678 2760
rect 11716 1766 11744 2746
rect 13004 2564 13032 4791
rect 13280 4690 13308 4927
rect 13268 4684 13320 4690
rect 13268 4626 13320 4632
rect 13372 4570 13400 7822
rect 13464 5302 13492 11727
rect 13648 10198 13676 13280
rect 13740 12238 13768 13330
rect 13820 12912 13872 12918
rect 13820 12854 13872 12860
rect 13832 12442 13860 12854
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13740 10198 13768 10406
rect 13636 10192 13688 10198
rect 13636 10134 13688 10140
rect 13728 10192 13780 10198
rect 13728 10134 13780 10140
rect 13648 9722 13676 10134
rect 13924 9926 13952 15422
rect 14004 13864 14056 13870
rect 14004 13806 14056 13812
rect 14016 13326 14044 13806
rect 14108 13734 14136 15535
rect 14096 13728 14148 13734
rect 14096 13670 14148 13676
rect 14004 13320 14056 13326
rect 14004 13262 14056 13268
rect 14016 12986 14044 13262
rect 14096 13184 14148 13190
rect 14096 13126 14148 13132
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 14016 12850 14044 12922
rect 14004 12844 14056 12850
rect 14004 12786 14056 12792
rect 14016 11694 14044 12786
rect 14108 12782 14136 13126
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 14200 12730 14228 18226
rect 14292 17513 14320 20182
rect 14476 19904 14504 35634
rect 15028 30258 15056 37062
rect 16040 35290 16068 37198
rect 16132 37126 16160 39200
rect 16776 37126 16804 39200
rect 18064 37262 18092 39200
rect 16948 37256 17000 37262
rect 16948 37198 17000 37204
rect 18052 37256 18104 37262
rect 18052 37198 18104 37204
rect 16120 37120 16172 37126
rect 16120 37062 16172 37068
rect 16764 37120 16816 37126
rect 16764 37062 16816 37068
rect 16028 35284 16080 35290
rect 16028 35226 16080 35232
rect 15476 31136 15528 31142
rect 15476 31078 15528 31084
rect 15016 30252 15068 30258
rect 15016 30194 15068 30200
rect 15016 29640 15068 29646
rect 15016 29582 15068 29588
rect 14740 27328 14792 27334
rect 14740 27270 14792 27276
rect 14556 26784 14608 26790
rect 14556 26726 14608 26732
rect 14568 24274 14596 26726
rect 14752 25906 14780 27270
rect 14740 25900 14792 25906
rect 14740 25842 14792 25848
rect 14648 25424 14700 25430
rect 14648 25366 14700 25372
rect 14660 24410 14688 25366
rect 14740 25220 14792 25226
rect 14740 25162 14792 25168
rect 14648 24404 14700 24410
rect 14648 24346 14700 24352
rect 14556 24268 14608 24274
rect 14556 24210 14608 24216
rect 14660 22778 14688 24346
rect 14648 22772 14700 22778
rect 14648 22714 14700 22720
rect 14752 22642 14780 25162
rect 14924 23724 14976 23730
rect 14924 23666 14976 23672
rect 14832 23520 14884 23526
rect 14832 23462 14884 23468
rect 14844 23050 14872 23462
rect 14832 23044 14884 23050
rect 14832 22986 14884 22992
rect 14936 22642 14964 23666
rect 15028 23474 15056 29582
rect 15384 26988 15436 26994
rect 15384 26930 15436 26936
rect 15200 26784 15252 26790
rect 15200 26726 15252 26732
rect 15108 26444 15160 26450
rect 15108 26386 15160 26392
rect 15120 25430 15148 26386
rect 15212 25906 15240 26726
rect 15396 26586 15424 26930
rect 15384 26580 15436 26586
rect 15384 26522 15436 26528
rect 15292 26240 15344 26246
rect 15292 26182 15344 26188
rect 15304 26042 15332 26182
rect 15292 26036 15344 26042
rect 15292 25978 15344 25984
rect 15200 25900 15252 25906
rect 15200 25842 15252 25848
rect 15200 25764 15252 25770
rect 15200 25706 15252 25712
rect 15108 25424 15160 25430
rect 15108 25366 15160 25372
rect 15212 25294 15240 25706
rect 15200 25288 15252 25294
rect 15252 25248 15332 25276
rect 15200 25230 15252 25236
rect 15200 25152 15252 25158
rect 15200 25094 15252 25100
rect 15212 24750 15240 25094
rect 15200 24744 15252 24750
rect 15200 24686 15252 24692
rect 15108 24676 15160 24682
rect 15108 24618 15160 24624
rect 15120 23594 15148 24618
rect 15212 24206 15240 24686
rect 15304 24206 15332 25248
rect 15200 24200 15252 24206
rect 15200 24142 15252 24148
rect 15292 24200 15344 24206
rect 15292 24142 15344 24148
rect 15292 23656 15344 23662
rect 15292 23598 15344 23604
rect 15108 23588 15160 23594
rect 15108 23530 15160 23536
rect 15304 23526 15332 23598
rect 15292 23520 15344 23526
rect 15028 23446 15148 23474
rect 15292 23462 15344 23468
rect 14740 22636 14792 22642
rect 14740 22578 14792 22584
rect 14924 22636 14976 22642
rect 14924 22578 14976 22584
rect 14556 22568 14608 22574
rect 14556 22510 14608 22516
rect 14568 21622 14596 22510
rect 14556 21616 14608 21622
rect 14556 21558 14608 21564
rect 14568 20856 14596 21558
rect 14648 20868 14700 20874
rect 14568 20828 14648 20856
rect 14648 20810 14700 20816
rect 14740 20868 14792 20874
rect 14740 20810 14792 20816
rect 14752 20602 14780 20810
rect 14740 20596 14792 20602
rect 14740 20538 14792 20544
rect 14384 19876 14504 19904
rect 14384 19446 14412 19876
rect 14464 19780 14516 19786
rect 14464 19722 14516 19728
rect 14372 19440 14424 19446
rect 14372 19382 14424 19388
rect 14372 19168 14424 19174
rect 14372 19110 14424 19116
rect 14384 18970 14412 19110
rect 14372 18964 14424 18970
rect 14372 18906 14424 18912
rect 14278 17504 14334 17513
rect 14278 17439 14334 17448
rect 14292 17202 14320 17439
rect 14280 17196 14332 17202
rect 14280 17138 14332 17144
rect 14384 16266 14412 18906
rect 14476 18426 14504 19722
rect 15120 19666 15148 23446
rect 15384 22024 15436 22030
rect 15382 21992 15384 22001
rect 15436 21992 15438 22001
rect 15200 21956 15252 21962
rect 15382 21927 15438 21936
rect 15200 21898 15252 21904
rect 15212 21690 15240 21898
rect 15200 21684 15252 21690
rect 15200 21626 15252 21632
rect 15384 21072 15436 21078
rect 15384 21014 15436 21020
rect 15292 20528 15344 20534
rect 15292 20470 15344 20476
rect 15028 19638 15148 19666
rect 14556 19168 14608 19174
rect 14556 19110 14608 19116
rect 14568 18698 14596 19110
rect 14556 18692 14608 18698
rect 14556 18634 14608 18640
rect 14740 18692 14792 18698
rect 14740 18634 14792 18640
rect 14464 18420 14516 18426
rect 14464 18362 14516 18368
rect 14648 18352 14700 18358
rect 14648 18294 14700 18300
rect 14660 18086 14688 18294
rect 14752 18086 14780 18634
rect 14924 18624 14976 18630
rect 14844 18584 14924 18612
rect 14648 18080 14700 18086
rect 14648 18022 14700 18028
rect 14740 18080 14792 18086
rect 14740 18022 14792 18028
rect 14648 17060 14700 17066
rect 14648 17002 14700 17008
rect 14464 16788 14516 16794
rect 14464 16730 14516 16736
rect 14476 16522 14504 16730
rect 14464 16516 14516 16522
rect 14464 16458 14516 16464
rect 14556 16448 14608 16454
rect 14556 16390 14608 16396
rect 14384 16238 14504 16266
rect 14372 16176 14424 16182
rect 14372 16118 14424 16124
rect 14384 15434 14412 16118
rect 14372 15428 14424 15434
rect 14372 15370 14424 15376
rect 14384 14958 14412 15370
rect 14372 14952 14424 14958
rect 14476 14940 14504 16238
rect 14568 15094 14596 16390
rect 14660 15434 14688 17002
rect 14752 16726 14780 18022
rect 14844 17678 14872 18584
rect 14924 18566 14976 18572
rect 14832 17672 14884 17678
rect 14832 17614 14884 17620
rect 14740 16720 14792 16726
rect 14740 16662 14792 16668
rect 14844 16574 14872 17614
rect 14924 17128 14976 17134
rect 14924 17070 14976 17076
rect 14936 16726 14964 17070
rect 14924 16720 14976 16726
rect 14924 16662 14976 16668
rect 14752 16546 14872 16574
rect 14648 15428 14700 15434
rect 14648 15370 14700 15376
rect 14556 15088 14608 15094
rect 14556 15030 14608 15036
rect 14476 14912 14596 14940
rect 14372 14894 14424 14900
rect 14280 14544 14332 14550
rect 14464 14544 14516 14550
rect 14332 14504 14464 14532
rect 14280 14486 14332 14492
rect 14464 14486 14516 14492
rect 14372 14340 14424 14346
rect 14372 14282 14424 14288
rect 14200 12702 14320 12730
rect 14188 12640 14240 12646
rect 14188 12582 14240 12588
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 14016 11082 14044 11630
rect 14096 11280 14148 11286
rect 14094 11248 14096 11257
rect 14148 11248 14150 11257
rect 14094 11183 14150 11192
rect 14004 11076 14056 11082
rect 14004 11018 14056 11024
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13636 9716 13688 9722
rect 13636 9658 13688 9664
rect 13542 9480 13598 9489
rect 13542 9415 13598 9424
rect 13452 5296 13504 5302
rect 13452 5238 13504 5244
rect 13556 5234 13584 9415
rect 13924 9110 13952 9862
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 14108 9178 14136 9318
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 13912 9104 13964 9110
rect 13912 9046 13964 9052
rect 14200 8906 14228 12582
rect 14292 9330 14320 12702
rect 14384 9654 14412 14282
rect 14464 13728 14516 13734
rect 14464 13670 14516 13676
rect 14476 12646 14504 13670
rect 14568 13394 14596 14912
rect 14556 13388 14608 13394
rect 14556 13330 14608 13336
rect 14752 12986 14780 16546
rect 15028 16182 15056 19638
rect 15304 19514 15332 20470
rect 15108 19508 15160 19514
rect 15108 19450 15160 19456
rect 15292 19508 15344 19514
rect 15292 19450 15344 19456
rect 15120 17626 15148 19450
rect 15396 18222 15424 21014
rect 15488 20398 15516 31078
rect 15568 30116 15620 30122
rect 15568 30058 15620 30064
rect 15580 23526 15608 30058
rect 15752 25900 15804 25906
rect 15752 25842 15804 25848
rect 15660 24064 15712 24070
rect 15660 24006 15712 24012
rect 15568 23520 15620 23526
rect 15672 23497 15700 24006
rect 15568 23462 15620 23468
rect 15658 23488 15714 23497
rect 15580 21486 15608 23462
rect 15658 23423 15714 23432
rect 15764 23050 15792 25842
rect 16396 25492 16448 25498
rect 16396 25434 16448 25440
rect 16408 25294 16436 25434
rect 16396 25288 16448 25294
rect 16396 25230 16448 25236
rect 16304 24812 16356 24818
rect 16304 24754 16356 24760
rect 15844 24132 15896 24138
rect 15844 24074 15896 24080
rect 15856 23866 15884 24074
rect 15844 23860 15896 23866
rect 15844 23802 15896 23808
rect 15856 23118 15884 23802
rect 15844 23112 15896 23118
rect 15844 23054 15896 23060
rect 15752 23044 15804 23050
rect 15752 22986 15804 22992
rect 16028 23044 16080 23050
rect 16028 22986 16080 22992
rect 15660 22976 15712 22982
rect 15660 22918 15712 22924
rect 15568 21480 15620 21486
rect 15568 21422 15620 21428
rect 15476 20392 15528 20398
rect 15476 20334 15528 20340
rect 15476 18692 15528 18698
rect 15476 18634 15528 18640
rect 15200 18216 15252 18222
rect 15200 18158 15252 18164
rect 15384 18216 15436 18222
rect 15384 18158 15436 18164
rect 15212 17746 15240 18158
rect 15488 18068 15516 18634
rect 15672 18204 15700 22918
rect 16040 22166 16068 22986
rect 16212 22568 16264 22574
rect 16212 22510 16264 22516
rect 16120 22500 16172 22506
rect 16120 22442 16172 22448
rect 16028 22160 16080 22166
rect 16028 22102 16080 22108
rect 16132 22030 16160 22442
rect 15844 22024 15896 22030
rect 15750 21992 15806 22001
rect 16120 22024 16172 22030
rect 15896 21984 15976 22012
rect 15844 21966 15896 21972
rect 15750 21927 15806 21936
rect 15764 21418 15792 21927
rect 15842 21856 15898 21865
rect 15842 21791 15898 21800
rect 15752 21412 15804 21418
rect 15752 21354 15804 21360
rect 15752 19372 15804 19378
rect 15752 19314 15804 19320
rect 15396 18040 15516 18068
rect 15580 18176 15700 18204
rect 15200 17740 15252 17746
rect 15200 17682 15252 17688
rect 15120 17610 15332 17626
rect 15120 17604 15344 17610
rect 15120 17598 15292 17604
rect 15292 17546 15344 17552
rect 15108 17060 15160 17066
rect 15108 17002 15160 17008
rect 15016 16176 15068 16182
rect 15016 16118 15068 16124
rect 14832 16108 14884 16114
rect 14832 16050 14884 16056
rect 14844 15337 14872 16050
rect 15120 15450 15148 17002
rect 15292 16516 15344 16522
rect 15292 16458 15344 16464
rect 15304 16046 15332 16458
rect 15292 16040 15344 16046
rect 15292 15982 15344 15988
rect 15200 15972 15252 15978
rect 15200 15914 15252 15920
rect 14936 15422 15148 15450
rect 14830 15328 14886 15337
rect 14830 15263 14886 15272
rect 14936 15178 14964 15422
rect 15016 15360 15068 15366
rect 15016 15302 15068 15308
rect 14844 15150 14964 15178
rect 14740 12980 14792 12986
rect 14740 12922 14792 12928
rect 14844 12866 14872 15150
rect 14924 15020 14976 15026
rect 14924 14962 14976 14968
rect 14936 14414 14964 14962
rect 15028 14822 15056 15302
rect 15212 15042 15240 15914
rect 15292 15700 15344 15706
rect 15292 15642 15344 15648
rect 15120 15014 15240 15042
rect 15120 14822 15148 15014
rect 15200 14952 15252 14958
rect 15200 14894 15252 14900
rect 15016 14816 15068 14822
rect 15016 14758 15068 14764
rect 15108 14816 15160 14822
rect 15108 14758 15160 14764
rect 14924 14408 14976 14414
rect 14924 14350 14976 14356
rect 15014 13968 15070 13977
rect 15014 13903 15070 13912
rect 14924 13388 14976 13394
rect 14924 13330 14976 13336
rect 14660 12838 14872 12866
rect 14464 12640 14516 12646
rect 14464 12582 14516 12588
rect 14660 12186 14688 12838
rect 14476 12158 14688 12186
rect 14832 12164 14884 12170
rect 14372 9648 14424 9654
rect 14372 9590 14424 9596
rect 14292 9302 14412 9330
rect 14280 9172 14332 9178
rect 14280 9114 14332 9120
rect 14188 8900 14240 8906
rect 14188 8842 14240 8848
rect 13636 8560 13688 8566
rect 13634 8528 13636 8537
rect 13688 8528 13690 8537
rect 13634 8463 13690 8472
rect 14096 7948 14148 7954
rect 14096 7890 14148 7896
rect 14188 7948 14240 7954
rect 14188 7890 14240 7896
rect 14108 7206 14136 7890
rect 14200 7410 14228 7890
rect 14292 7546 14320 9114
rect 14280 7540 14332 7546
rect 14280 7482 14332 7488
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 14200 7274 14228 7346
rect 14188 7268 14240 7274
rect 14188 7210 14240 7216
rect 14096 7200 14148 7206
rect 14096 7142 14148 7148
rect 13728 6928 13780 6934
rect 13728 6870 13780 6876
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13544 5228 13596 5234
rect 13544 5170 13596 5176
rect 13280 4542 13400 4570
rect 13280 4282 13308 4542
rect 13544 4480 13596 4486
rect 13544 4422 13596 4428
rect 13268 4276 13320 4282
rect 13268 4218 13320 4224
rect 13280 3602 13308 4218
rect 13360 3936 13412 3942
rect 13360 3878 13412 3884
rect 13452 3936 13504 3942
rect 13452 3878 13504 3884
rect 13268 3596 13320 3602
rect 13268 3538 13320 3544
rect 13176 3460 13228 3466
rect 13176 3402 13228 3408
rect 12912 2536 13032 2564
rect 12256 2372 12308 2378
rect 12256 2314 12308 2320
rect 11704 1760 11756 1766
rect 11704 1702 11756 1708
rect 12268 1630 12296 2314
rect 12256 1624 12308 1630
rect 12256 1566 12308 1572
rect 12912 800 12940 2536
rect 8496 734 8800 762
rect 9678 200 9734 800
rect 10322 200 10378 800
rect 11610 200 11666 800
rect 12898 200 12954 800
rect 13188 762 13216 3402
rect 13372 3398 13400 3878
rect 13360 3392 13412 3398
rect 13360 3334 13412 3340
rect 13268 3052 13320 3058
rect 13268 2994 13320 3000
rect 13280 2514 13308 2994
rect 13360 2848 13412 2854
rect 13358 2816 13360 2825
rect 13412 2816 13414 2825
rect 13358 2751 13414 2760
rect 13268 2508 13320 2514
rect 13268 2450 13320 2456
rect 13464 1834 13492 3878
rect 13556 3126 13584 4422
rect 13544 3120 13596 3126
rect 13648 3097 13676 6054
rect 13740 5778 13768 6870
rect 14200 6866 14228 7210
rect 14188 6860 14240 6866
rect 14188 6802 14240 6808
rect 14200 6390 14228 6802
rect 14384 6769 14412 9302
rect 14370 6760 14426 6769
rect 14370 6695 14426 6704
rect 14384 6390 14412 6695
rect 14188 6384 14240 6390
rect 14188 6326 14240 6332
rect 14372 6384 14424 6390
rect 14372 6326 14424 6332
rect 14200 5778 14228 6326
rect 14372 5908 14424 5914
rect 14372 5850 14424 5856
rect 13728 5772 13780 5778
rect 13728 5714 13780 5720
rect 14188 5772 14240 5778
rect 14188 5714 14240 5720
rect 14384 5574 14412 5850
rect 14372 5568 14424 5574
rect 14372 5510 14424 5516
rect 13820 5296 13872 5302
rect 13820 5238 13872 5244
rect 13832 5030 13860 5238
rect 14476 5166 14504 12158
rect 14832 12106 14884 12112
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 14568 11082 14596 11834
rect 14844 11082 14872 12106
rect 14556 11076 14608 11082
rect 14556 11018 14608 11024
rect 14832 11076 14884 11082
rect 14832 11018 14884 11024
rect 14740 9648 14792 9654
rect 14740 9590 14792 9596
rect 14648 9580 14700 9586
rect 14648 9522 14700 9528
rect 14660 8634 14688 9522
rect 14648 8628 14700 8634
rect 14648 8570 14700 8576
rect 14556 8288 14608 8294
rect 14556 8230 14608 8236
rect 14568 8022 14596 8230
rect 14556 8016 14608 8022
rect 14556 7958 14608 7964
rect 14646 5808 14702 5817
rect 14646 5743 14702 5752
rect 14660 5370 14688 5743
rect 14556 5364 14608 5370
rect 14556 5306 14608 5312
rect 14648 5364 14700 5370
rect 14648 5306 14700 5312
rect 14568 5166 14596 5306
rect 14188 5160 14240 5166
rect 14464 5160 14516 5166
rect 14240 5120 14320 5148
rect 14188 5102 14240 5108
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 14292 4622 14320 5120
rect 14464 5102 14516 5108
rect 14556 5160 14608 5166
rect 14556 5102 14608 5108
rect 14646 5128 14702 5137
rect 14476 4758 14504 5102
rect 14752 5114 14780 9590
rect 14702 5086 14780 5114
rect 14646 5063 14702 5072
rect 14464 4752 14516 4758
rect 14464 4694 14516 4700
rect 14280 4616 14332 4622
rect 14660 4593 14688 5063
rect 14280 4558 14332 4564
rect 14646 4584 14702 4593
rect 14292 4078 14320 4558
rect 14646 4519 14702 4528
rect 14830 4584 14886 4593
rect 14830 4519 14832 4528
rect 14884 4519 14886 4528
rect 14832 4490 14884 4496
rect 14280 4072 14332 4078
rect 14280 4014 14332 4020
rect 14554 4040 14610 4049
rect 14188 3664 14240 3670
rect 14188 3606 14240 3612
rect 13912 3460 13964 3466
rect 13912 3402 13964 3408
rect 13544 3062 13596 3068
rect 13634 3088 13690 3097
rect 13556 2774 13584 3062
rect 13634 3023 13690 3032
rect 13556 2746 13676 2774
rect 13648 2310 13676 2746
rect 13924 2514 13952 3402
rect 14200 3346 14228 3606
rect 14292 3534 14320 4014
rect 14554 3975 14610 3984
rect 14568 3942 14596 3975
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 14464 3460 14516 3466
rect 14464 3402 14516 3408
rect 14476 3346 14504 3402
rect 14200 3318 14504 3346
rect 14476 2689 14504 3318
rect 14830 3088 14886 3097
rect 14830 3023 14886 3032
rect 14844 2990 14872 3023
rect 14936 2990 14964 13330
rect 15028 13258 15056 13903
rect 15212 13530 15240 14894
rect 15304 14414 15332 15642
rect 15396 15473 15424 18040
rect 15580 16658 15608 18176
rect 15660 17536 15712 17542
rect 15660 17478 15712 17484
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 15476 16584 15528 16590
rect 15476 16526 15528 16532
rect 15382 15464 15438 15473
rect 15382 15399 15438 15408
rect 15488 15416 15516 16526
rect 15580 16046 15608 16594
rect 15672 16182 15700 17478
rect 15660 16176 15712 16182
rect 15660 16118 15712 16124
rect 15568 16040 15620 16046
rect 15568 15982 15620 15988
rect 15568 15428 15620 15434
rect 15488 15388 15568 15416
rect 15568 15370 15620 15376
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 15200 13524 15252 13530
rect 15200 13466 15252 13472
rect 15016 13252 15068 13258
rect 15016 13194 15068 13200
rect 15016 12980 15068 12986
rect 15016 12922 15068 12928
rect 15028 9586 15056 12922
rect 15212 10962 15240 13466
rect 15304 12434 15332 14350
rect 15396 14006 15424 14962
rect 15384 14000 15436 14006
rect 15436 13960 15516 13988
rect 15384 13942 15436 13948
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 15396 12782 15424 12922
rect 15384 12776 15436 12782
rect 15384 12718 15436 12724
rect 15304 12406 15424 12434
rect 15290 11248 15346 11257
rect 15290 11183 15346 11192
rect 15120 10934 15240 10962
rect 15120 10130 15148 10934
rect 15200 10804 15252 10810
rect 15200 10746 15252 10752
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 15212 9994 15240 10746
rect 15304 10742 15332 11183
rect 15292 10736 15344 10742
rect 15292 10678 15344 10684
rect 15200 9988 15252 9994
rect 15200 9930 15252 9936
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 15016 9580 15068 9586
rect 15016 9522 15068 9528
rect 15108 9444 15160 9450
rect 15108 9386 15160 9392
rect 15016 9376 15068 9382
rect 15016 9318 15068 9324
rect 15028 3126 15056 9318
rect 15120 8906 15148 9386
rect 15108 8900 15160 8906
rect 15108 8842 15160 8848
rect 15106 8664 15162 8673
rect 15106 8599 15162 8608
rect 15120 8566 15148 8599
rect 15108 8560 15160 8566
rect 15108 8502 15160 8508
rect 15200 7472 15252 7478
rect 15200 7414 15252 7420
rect 15212 6458 15240 7414
rect 15200 6452 15252 6458
rect 15200 6394 15252 6400
rect 15304 6390 15332 9862
rect 15396 9722 15424 12406
rect 15488 12238 15516 13960
rect 15580 12306 15608 15370
rect 15764 14618 15792 19314
rect 15856 18329 15884 21791
rect 15948 21622 15976 21984
rect 16120 21966 16172 21972
rect 16120 21888 16172 21894
rect 16120 21830 16172 21836
rect 16132 21706 16160 21830
rect 16040 21690 16160 21706
rect 16028 21684 16160 21690
rect 16080 21678 16160 21684
rect 16028 21626 16080 21632
rect 15936 21616 15988 21622
rect 15936 21558 15988 21564
rect 15948 21146 15976 21558
rect 15936 21140 15988 21146
rect 15936 21082 15988 21088
rect 15936 20868 15988 20874
rect 15936 20810 15988 20816
rect 15948 20534 15976 20810
rect 15936 20528 15988 20534
rect 15936 20470 15988 20476
rect 16120 19780 16172 19786
rect 16120 19722 16172 19728
rect 16132 19446 16160 19722
rect 16224 19514 16252 22510
rect 16212 19508 16264 19514
rect 16212 19450 16264 19456
rect 16120 19440 16172 19446
rect 15934 19408 15990 19417
rect 16120 19382 16172 19388
rect 15934 19343 15936 19352
rect 15988 19343 15990 19352
rect 15936 19314 15988 19320
rect 15842 18320 15898 18329
rect 15842 18255 15898 18264
rect 15856 18222 15884 18255
rect 15844 18216 15896 18222
rect 15844 18158 15896 18164
rect 15844 17604 15896 17610
rect 15844 17546 15896 17552
rect 15856 15978 15884 17546
rect 15948 17202 15976 19314
rect 16224 18834 16252 19450
rect 16212 18828 16264 18834
rect 16212 18770 16264 18776
rect 16120 18692 16172 18698
rect 16120 18634 16172 18640
rect 16132 18154 16160 18634
rect 16212 18216 16264 18222
rect 16212 18158 16264 18164
rect 16120 18148 16172 18154
rect 16120 18090 16172 18096
rect 16118 17640 16174 17649
rect 16118 17575 16174 17584
rect 16132 17202 16160 17575
rect 15936 17196 15988 17202
rect 15936 17138 15988 17144
rect 16120 17196 16172 17202
rect 16120 17138 16172 17144
rect 16028 16788 16080 16794
rect 16028 16730 16080 16736
rect 15936 16516 15988 16522
rect 15936 16458 15988 16464
rect 15844 15972 15896 15978
rect 15844 15914 15896 15920
rect 15844 15700 15896 15706
rect 15844 15642 15896 15648
rect 15752 14612 15804 14618
rect 15752 14554 15804 14560
rect 15658 13560 15714 13569
rect 15658 13495 15714 13504
rect 15672 12730 15700 13495
rect 15752 12776 15804 12782
rect 15672 12724 15752 12730
rect 15672 12718 15804 12724
rect 15672 12702 15792 12718
rect 15568 12300 15620 12306
rect 15568 12242 15620 12248
rect 15476 12232 15528 12238
rect 15476 12174 15528 12180
rect 15580 12073 15608 12242
rect 15566 12064 15622 12073
rect 15566 11999 15622 12008
rect 15476 10056 15528 10062
rect 15476 9998 15528 10004
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 15488 9654 15516 9998
rect 15476 9648 15528 9654
rect 15476 9590 15528 9596
rect 15384 9036 15436 9042
rect 15488 9024 15516 9590
rect 15436 8996 15516 9024
rect 15384 8978 15436 8984
rect 15672 7449 15700 12702
rect 15856 12594 15884 15642
rect 15764 12566 15884 12594
rect 15764 12442 15792 12566
rect 15752 12436 15804 12442
rect 15752 12378 15804 12384
rect 15764 11898 15792 12378
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 15844 10668 15896 10674
rect 15844 10610 15896 10616
rect 15750 8800 15806 8809
rect 15750 8735 15806 8744
rect 15658 7440 15714 7449
rect 15658 7375 15714 7384
rect 15292 6384 15344 6390
rect 15292 6326 15344 6332
rect 15108 5636 15160 5642
rect 15108 5578 15160 5584
rect 15120 5545 15148 5578
rect 15106 5536 15162 5545
rect 15106 5471 15162 5480
rect 15660 5160 15712 5166
rect 15660 5102 15712 5108
rect 15108 4548 15160 4554
rect 15108 4490 15160 4496
rect 15120 3233 15148 4490
rect 15106 3224 15162 3233
rect 15106 3159 15162 3168
rect 15016 3120 15068 3126
rect 15016 3062 15068 3068
rect 14832 2984 14884 2990
rect 14832 2926 14884 2932
rect 14924 2984 14976 2990
rect 14924 2926 14976 2932
rect 14832 2848 14884 2854
rect 14832 2790 14884 2796
rect 14462 2680 14518 2689
rect 14462 2615 14518 2624
rect 13912 2508 13964 2514
rect 13912 2450 13964 2456
rect 13636 2304 13688 2310
rect 13636 2246 13688 2252
rect 13452 1828 13504 1834
rect 13452 1770 13504 1776
rect 13464 870 13584 898
rect 13464 762 13492 870
rect 13556 800 13584 870
rect 14844 800 14872 2790
rect 15672 2774 15700 5102
rect 15488 2746 15700 2774
rect 15488 2514 15516 2746
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 15292 2372 15344 2378
rect 15292 2314 15344 2320
rect 15304 2038 15332 2314
rect 15292 2032 15344 2038
rect 15292 1974 15344 1980
rect 15488 1970 15516 2450
rect 15764 1970 15792 8735
rect 15856 8294 15884 10610
rect 15844 8288 15896 8294
rect 15844 8230 15896 8236
rect 15856 7546 15884 8230
rect 15844 7540 15896 7546
rect 15844 7482 15896 7488
rect 15948 5574 15976 16458
rect 16040 10810 16068 16730
rect 16120 16244 16172 16250
rect 16120 16186 16172 16192
rect 16132 15978 16160 16186
rect 16120 15972 16172 15978
rect 16120 15914 16172 15920
rect 16224 15858 16252 18158
rect 16316 16794 16344 24754
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 16132 15830 16252 15858
rect 16132 15706 16160 15830
rect 16408 15722 16436 25230
rect 16856 24336 16908 24342
rect 16856 24278 16908 24284
rect 16868 23730 16896 24278
rect 16856 23724 16908 23730
rect 16856 23666 16908 23672
rect 16488 23112 16540 23118
rect 16488 23054 16540 23060
rect 16500 22506 16528 23054
rect 16488 22500 16540 22506
rect 16488 22442 16540 22448
rect 16580 22432 16632 22438
rect 16580 22374 16632 22380
rect 16488 22024 16540 22030
rect 16488 21966 16540 21972
rect 16500 21486 16528 21966
rect 16488 21480 16540 21486
rect 16488 21422 16540 21428
rect 16592 20806 16620 22374
rect 16960 22094 16988 37198
rect 17132 37120 17184 37126
rect 17132 37062 17184 37068
rect 17144 31346 17172 37062
rect 19352 36922 19380 39200
rect 19996 37126 20024 39200
rect 20168 37392 20220 37398
rect 20168 37334 20220 37340
rect 20076 37256 20128 37262
rect 20076 37198 20128 37204
rect 19984 37120 20036 37126
rect 19984 37062 20036 37068
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19340 36916 19392 36922
rect 19340 36858 19392 36864
rect 19432 36780 19484 36786
rect 19432 36722 19484 36728
rect 19444 33658 19472 36722
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19432 33652 19484 33658
rect 19432 33594 19484 33600
rect 18604 33312 18656 33318
rect 18604 33254 18656 33260
rect 17132 31340 17184 31346
rect 17132 31282 17184 31288
rect 18420 30660 18472 30666
rect 18420 30602 18472 30608
rect 17960 30388 18012 30394
rect 17960 30330 18012 30336
rect 17592 29028 17644 29034
rect 17592 28970 17644 28976
rect 17224 25152 17276 25158
rect 17224 25094 17276 25100
rect 17040 23520 17092 23526
rect 17040 23462 17092 23468
rect 17052 23186 17080 23462
rect 17040 23180 17092 23186
rect 17040 23122 17092 23128
rect 17236 22710 17264 25094
rect 17224 22704 17276 22710
rect 17224 22646 17276 22652
rect 17224 22160 17276 22166
rect 17224 22102 17276 22108
rect 16960 22066 17172 22094
rect 16856 22024 16908 22030
rect 16856 21966 16908 21972
rect 16580 20800 16632 20806
rect 16580 20742 16632 20748
rect 16868 20602 16896 21966
rect 16946 21040 17002 21049
rect 16946 20975 16948 20984
rect 17000 20975 17002 20984
rect 16948 20946 17000 20952
rect 16856 20596 16908 20602
rect 16856 20538 16908 20544
rect 16580 20528 16632 20534
rect 16580 20470 16632 20476
rect 16488 19304 16540 19310
rect 16488 19246 16540 19252
rect 16500 18630 16528 19246
rect 16488 18624 16540 18630
rect 16488 18566 16540 18572
rect 16488 17604 16540 17610
rect 16488 17546 16540 17552
rect 16500 17338 16528 17546
rect 16488 17332 16540 17338
rect 16488 17274 16540 17280
rect 16488 16652 16540 16658
rect 16488 16594 16540 16600
rect 16120 15700 16172 15706
rect 16120 15642 16172 15648
rect 16224 15694 16436 15722
rect 16120 14476 16172 14482
rect 16120 14418 16172 14424
rect 16132 14385 16160 14418
rect 16118 14376 16174 14385
rect 16118 14311 16174 14320
rect 16120 13864 16172 13870
rect 16120 13806 16172 13812
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 16132 10674 16160 13806
rect 16224 12986 16252 15694
rect 16500 15552 16528 16594
rect 16592 16153 16620 20470
rect 17144 20262 17172 22066
rect 17132 20256 17184 20262
rect 17132 20198 17184 20204
rect 17236 20058 17264 22102
rect 17500 21616 17552 21622
rect 17500 21558 17552 21564
rect 17408 21344 17460 21350
rect 17408 21286 17460 21292
rect 17420 21049 17448 21286
rect 17406 21040 17462 21049
rect 17406 20975 17462 20984
rect 17316 20528 17368 20534
rect 17316 20470 17368 20476
rect 17224 20052 17276 20058
rect 17224 19994 17276 20000
rect 17040 19712 17092 19718
rect 17040 19654 17092 19660
rect 16670 19000 16726 19009
rect 16670 18935 16726 18944
rect 16684 18834 16712 18935
rect 16672 18828 16724 18834
rect 16672 18770 16724 18776
rect 16684 17134 16712 18770
rect 17052 18358 17080 19654
rect 17132 18964 17184 18970
rect 17132 18906 17184 18912
rect 17144 18766 17172 18906
rect 17132 18760 17184 18766
rect 17132 18702 17184 18708
rect 17040 18352 17092 18358
rect 17040 18294 17092 18300
rect 16764 17740 16816 17746
rect 16764 17682 16816 17688
rect 16776 17202 16804 17682
rect 17132 17264 17184 17270
rect 17132 17206 17184 17212
rect 16764 17196 16816 17202
rect 16764 17138 16816 17144
rect 16672 17128 16724 17134
rect 16672 17070 16724 17076
rect 17144 16794 17172 17206
rect 17132 16788 17184 16794
rect 17132 16730 17184 16736
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 16764 16584 16816 16590
rect 16764 16526 16816 16532
rect 16684 16182 16712 16526
rect 16672 16176 16724 16182
rect 16578 16144 16634 16153
rect 16672 16118 16724 16124
rect 16578 16079 16634 16088
rect 16408 15524 16528 15552
rect 16304 14952 16356 14958
rect 16304 14894 16356 14900
rect 16316 14385 16344 14894
rect 16302 14376 16358 14385
rect 16302 14311 16358 14320
rect 16304 13184 16356 13190
rect 16304 13126 16356 13132
rect 16212 12980 16264 12986
rect 16212 12922 16264 12928
rect 16120 10668 16172 10674
rect 16120 10610 16172 10616
rect 16120 10464 16172 10470
rect 16120 10406 16172 10412
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 16040 9586 16068 10202
rect 16028 9580 16080 9586
rect 16028 9522 16080 9528
rect 16132 8514 16160 10406
rect 16224 9518 16252 12922
rect 16316 12782 16344 13126
rect 16304 12776 16356 12782
rect 16304 12718 16356 12724
rect 16304 11076 16356 11082
rect 16304 11018 16356 11024
rect 16316 10849 16344 11018
rect 16302 10840 16358 10849
rect 16302 10775 16358 10784
rect 16304 10124 16356 10130
rect 16304 10066 16356 10072
rect 16212 9512 16264 9518
rect 16212 9454 16264 9460
rect 16316 9081 16344 10066
rect 16302 9072 16358 9081
rect 16302 9007 16358 9016
rect 16040 8486 16160 8514
rect 16040 6866 16068 8486
rect 16120 8424 16172 8430
rect 16120 8366 16172 8372
rect 16132 7954 16160 8366
rect 16120 7948 16172 7954
rect 16120 7890 16172 7896
rect 16408 7834 16436 15524
rect 16672 14816 16724 14822
rect 16672 14758 16724 14764
rect 16580 13796 16632 13802
rect 16580 13738 16632 13744
rect 16592 13326 16620 13738
rect 16580 13320 16632 13326
rect 16580 13262 16632 13268
rect 16592 12782 16620 13262
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 16592 12306 16620 12718
rect 16580 12300 16632 12306
rect 16580 12242 16632 12248
rect 16488 12164 16540 12170
rect 16488 12106 16540 12112
rect 16500 11898 16528 12106
rect 16488 11892 16540 11898
rect 16488 11834 16540 11840
rect 16592 11762 16620 12242
rect 16684 12170 16712 14758
rect 16672 12164 16724 12170
rect 16672 12106 16724 12112
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 16592 11218 16620 11698
rect 16672 11688 16724 11694
rect 16672 11630 16724 11636
rect 16684 11218 16712 11630
rect 16580 11212 16632 11218
rect 16580 11154 16632 11160
rect 16672 11212 16724 11218
rect 16672 11154 16724 11160
rect 16488 9172 16540 9178
rect 16488 9114 16540 9120
rect 16224 7806 16436 7834
rect 16224 7342 16252 7806
rect 16304 7744 16356 7750
rect 16500 7698 16528 9114
rect 16578 9072 16634 9081
rect 16578 9007 16634 9016
rect 16592 8974 16620 9007
rect 16580 8968 16632 8974
rect 16580 8910 16632 8916
rect 16672 8832 16724 8838
rect 16672 8774 16724 8780
rect 16684 7818 16712 8774
rect 16776 8090 16804 16526
rect 17132 16040 17184 16046
rect 17132 15982 17184 15988
rect 17144 15609 17172 15982
rect 17328 15978 17356 20470
rect 17408 19848 17460 19854
rect 17408 19790 17460 19796
rect 17420 19514 17448 19790
rect 17408 19508 17460 19514
rect 17408 19450 17460 19456
rect 17316 15972 17368 15978
rect 17316 15914 17368 15920
rect 17130 15600 17186 15609
rect 17130 15535 17186 15544
rect 17132 15428 17184 15434
rect 17132 15370 17184 15376
rect 16856 14612 16908 14618
rect 16856 14554 16908 14560
rect 17040 14612 17092 14618
rect 17040 14554 17092 14560
rect 16868 13258 16896 14554
rect 16948 14408 17000 14414
rect 16948 14350 17000 14356
rect 16856 13252 16908 13258
rect 16856 13194 16908 13200
rect 16868 10130 16896 13194
rect 16960 12753 16988 14350
rect 17052 14346 17080 14554
rect 17040 14340 17092 14346
rect 17040 14282 17092 14288
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 16946 12744 17002 12753
rect 16946 12679 17002 12688
rect 17052 11082 17080 13466
rect 17144 11642 17172 15370
rect 17316 14272 17368 14278
rect 17316 14214 17368 14220
rect 17224 13728 17276 13734
rect 17224 13670 17276 13676
rect 17236 12918 17264 13670
rect 17328 13258 17356 14214
rect 17512 13530 17540 21558
rect 17604 20398 17632 28970
rect 17684 27600 17736 27606
rect 17684 27542 17736 27548
rect 17696 24342 17724 27542
rect 17972 26314 18000 30330
rect 17960 26308 18012 26314
rect 17960 26250 18012 26256
rect 18236 26308 18288 26314
rect 18236 26250 18288 26256
rect 17960 25832 18012 25838
rect 17960 25774 18012 25780
rect 17972 25430 18000 25774
rect 17960 25424 18012 25430
rect 17960 25366 18012 25372
rect 17684 24336 17736 24342
rect 17684 24278 17736 24284
rect 17972 22574 18000 25366
rect 18052 24744 18104 24750
rect 18052 24686 18104 24692
rect 17960 22568 18012 22574
rect 17960 22510 18012 22516
rect 17960 22432 18012 22438
rect 17960 22374 18012 22380
rect 17972 22250 18000 22374
rect 17788 22222 18000 22250
rect 17788 21962 17816 22222
rect 17868 22160 17920 22166
rect 17868 22102 17920 22108
rect 17776 21956 17828 21962
rect 17776 21898 17828 21904
rect 17880 21622 17908 22102
rect 17960 22092 18012 22098
rect 17960 22034 18012 22040
rect 17868 21616 17920 21622
rect 17868 21558 17920 21564
rect 17972 21350 18000 22034
rect 17684 21344 17736 21350
rect 17960 21344 18012 21350
rect 17684 21286 17736 21292
rect 17958 21312 17960 21321
rect 18012 21312 18014 21321
rect 17696 20806 17724 21286
rect 17958 21247 18014 21256
rect 17972 21221 18000 21247
rect 18064 21146 18092 24686
rect 18248 22094 18276 26250
rect 18432 25974 18460 30602
rect 18420 25968 18472 25974
rect 18420 25910 18472 25916
rect 18328 24200 18380 24206
rect 18328 24142 18380 24148
rect 18340 24041 18368 24142
rect 18326 24032 18382 24041
rect 18326 23967 18382 23976
rect 18340 23526 18368 23967
rect 18616 23730 18644 33254
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 20088 26976 20116 37198
rect 20180 31754 20208 37334
rect 21180 37256 21232 37262
rect 21180 37198 21232 37204
rect 20180 31726 20484 31754
rect 20088 26948 20300 26976
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19524 25968 19576 25974
rect 19524 25910 19576 25916
rect 19340 25900 19392 25906
rect 19340 25842 19392 25848
rect 19248 25832 19300 25838
rect 19248 25774 19300 25780
rect 19260 24954 19288 25774
rect 19352 25294 19380 25842
rect 19536 25498 19564 25910
rect 19524 25492 19576 25498
rect 19524 25434 19576 25440
rect 19340 25288 19392 25294
rect 19340 25230 19392 25236
rect 19248 24948 19300 24954
rect 19248 24890 19300 24896
rect 18788 24064 18840 24070
rect 18788 24006 18840 24012
rect 18800 23730 18828 24006
rect 18604 23724 18656 23730
rect 18604 23666 18656 23672
rect 18788 23724 18840 23730
rect 18788 23666 18840 23672
rect 18328 23520 18380 23526
rect 18328 23462 18380 23468
rect 18972 23180 19024 23186
rect 18972 23122 19024 23128
rect 18604 22636 18656 22642
rect 18604 22578 18656 22584
rect 18248 22066 18368 22094
rect 18340 21486 18368 22066
rect 18616 21865 18644 22578
rect 18602 21856 18658 21865
rect 18602 21791 18658 21800
rect 18984 21622 19012 23122
rect 19260 22574 19288 24890
rect 19248 22568 19300 22574
rect 19248 22510 19300 22516
rect 18420 21616 18472 21622
rect 18420 21558 18472 21564
rect 18972 21616 19024 21622
rect 18972 21558 19024 21564
rect 18328 21480 18380 21486
rect 18328 21422 18380 21428
rect 18052 21140 18104 21146
rect 18052 21082 18104 21088
rect 18144 21072 18196 21078
rect 18144 21014 18196 21020
rect 17776 20868 17828 20874
rect 17776 20810 17828 20816
rect 17684 20800 17736 20806
rect 17684 20742 17736 20748
rect 17592 20392 17644 20398
rect 17592 20334 17644 20340
rect 17788 20330 17816 20810
rect 18156 20534 18184 21014
rect 18328 20868 18380 20874
rect 18328 20810 18380 20816
rect 18144 20528 18196 20534
rect 18144 20470 18196 20476
rect 18156 20330 18184 20470
rect 17776 20324 17828 20330
rect 17776 20266 17828 20272
rect 18144 20324 18196 20330
rect 18144 20266 18196 20272
rect 17684 19780 17736 19786
rect 17684 19722 17736 19728
rect 17696 18970 17724 19722
rect 17684 18964 17736 18970
rect 17684 18906 17736 18912
rect 17684 16584 17736 16590
rect 17684 16526 17736 16532
rect 17592 15904 17644 15910
rect 17592 15846 17644 15852
rect 17604 15094 17632 15846
rect 17592 15088 17644 15094
rect 17592 15030 17644 15036
rect 17592 14272 17644 14278
rect 17592 14214 17644 14220
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17316 13252 17368 13258
rect 17316 13194 17368 13200
rect 17224 12912 17276 12918
rect 17224 12854 17276 12860
rect 17500 12640 17552 12646
rect 17500 12582 17552 12588
rect 17512 12434 17540 12582
rect 17420 12406 17540 12434
rect 17420 11830 17448 12406
rect 17408 11824 17460 11830
rect 17408 11766 17460 11772
rect 17144 11614 17356 11642
rect 17132 11552 17184 11558
rect 17132 11494 17184 11500
rect 17040 11076 17092 11082
rect 17040 11018 17092 11024
rect 16948 10600 17000 10606
rect 16948 10542 17000 10548
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 16960 9586 16988 10542
rect 16948 9580 17000 9586
rect 16868 9540 16948 9568
rect 16868 9042 16896 9540
rect 16948 9522 17000 9528
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 16868 8498 16896 8978
rect 17144 8566 17172 11494
rect 17328 10198 17356 11614
rect 17316 10192 17368 10198
rect 17316 10134 17368 10140
rect 17132 8560 17184 8566
rect 17132 8502 17184 8508
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 16672 7812 16724 7818
rect 16672 7754 16724 7760
rect 16356 7692 16528 7698
rect 16304 7686 16528 7692
rect 16316 7670 16528 7686
rect 16500 7410 16528 7670
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 16212 7336 16264 7342
rect 16212 7278 16264 7284
rect 16028 6860 16080 6866
rect 16028 6802 16080 6808
rect 16224 5778 16252 7278
rect 16394 7168 16450 7177
rect 16394 7103 16450 7112
rect 16212 5772 16264 5778
rect 16212 5714 16264 5720
rect 15936 5568 15988 5574
rect 15936 5510 15988 5516
rect 15948 5370 15976 5510
rect 15936 5364 15988 5370
rect 15936 5306 15988 5312
rect 16120 5364 16172 5370
rect 16120 5306 16172 5312
rect 16026 5264 16082 5273
rect 16026 5199 16082 5208
rect 16040 4593 16068 5199
rect 16132 5166 16160 5306
rect 16120 5160 16172 5166
rect 16120 5102 16172 5108
rect 16304 5024 16356 5030
rect 16304 4966 16356 4972
rect 16316 4758 16344 4966
rect 16304 4752 16356 4758
rect 16304 4694 16356 4700
rect 16026 4584 16082 4593
rect 16026 4519 16082 4528
rect 16040 3738 16068 4519
rect 16210 4176 16266 4185
rect 16210 4111 16266 4120
rect 16028 3732 16080 3738
rect 16028 3674 16080 3680
rect 16120 3052 16172 3058
rect 16120 2994 16172 3000
rect 15476 1964 15528 1970
rect 15476 1906 15528 1912
rect 15752 1964 15804 1970
rect 15752 1906 15804 1912
rect 16132 800 16160 2994
rect 16224 2310 16252 4111
rect 16302 3904 16358 3913
rect 16302 3839 16358 3848
rect 16316 3126 16344 3839
rect 16304 3120 16356 3126
rect 16304 3062 16356 3068
rect 16408 2774 16436 7103
rect 16776 6458 16804 8026
rect 16868 7954 16896 8434
rect 16856 7948 16908 7954
rect 16856 7890 16908 7896
rect 17224 7404 17276 7410
rect 17224 7346 17276 7352
rect 17236 6866 17264 7346
rect 17420 7041 17448 11766
rect 17604 9994 17632 14214
rect 17696 10470 17724 16526
rect 17788 15162 17816 20266
rect 17960 19372 18012 19378
rect 17960 19314 18012 19320
rect 17972 17746 18000 19314
rect 18236 19304 18288 19310
rect 18236 19246 18288 19252
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 18052 18284 18104 18290
rect 18052 18226 18104 18232
rect 17960 17740 18012 17746
rect 17960 17682 18012 17688
rect 17960 17128 18012 17134
rect 17958 17096 17960 17105
rect 18012 17096 18014 17105
rect 17958 17031 18014 17040
rect 17868 15904 17920 15910
rect 17868 15846 17920 15852
rect 17776 15156 17828 15162
rect 17776 15098 17828 15104
rect 17776 14340 17828 14346
rect 17776 14282 17828 14288
rect 17788 13870 17816 14282
rect 17776 13864 17828 13870
rect 17776 13806 17828 13812
rect 17880 11830 17908 15846
rect 17958 15464 18014 15473
rect 17958 15399 17960 15408
rect 18012 15399 18014 15408
rect 17960 15370 18012 15376
rect 17960 14816 18012 14822
rect 17960 14758 18012 14764
rect 17868 11824 17920 11830
rect 17868 11766 17920 11772
rect 17972 10742 18000 14758
rect 18064 11218 18092 18226
rect 18156 14958 18184 19110
rect 18248 17762 18276 19246
rect 18340 18426 18368 20810
rect 18432 18426 18460 21558
rect 18512 21480 18564 21486
rect 18512 21422 18564 21428
rect 18524 19378 18552 21422
rect 18604 21072 18656 21078
rect 18602 21040 18604 21049
rect 18656 21040 18658 21049
rect 18984 21010 19012 21558
rect 18602 20975 18658 20984
rect 18972 21004 19024 21010
rect 18972 20946 19024 20952
rect 19352 20618 19380 25230
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19984 24812 20036 24818
rect 19984 24754 20036 24760
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19432 22976 19484 22982
rect 19432 22918 19484 22924
rect 19444 22710 19472 22918
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19432 22704 19484 22710
rect 19432 22646 19484 22652
rect 19708 22228 19760 22234
rect 19708 22170 19760 22176
rect 19720 21894 19748 22170
rect 19432 21888 19484 21894
rect 19432 21830 19484 21836
rect 19708 21888 19760 21894
rect 19708 21830 19760 21836
rect 19444 21690 19472 21830
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19432 21684 19484 21690
rect 19432 21626 19484 21632
rect 19524 21616 19576 21622
rect 19524 21558 19576 21564
rect 19536 20942 19564 21558
rect 19616 21480 19668 21486
rect 19616 21422 19668 21428
rect 19628 21010 19656 21422
rect 19616 21004 19668 21010
rect 19616 20946 19668 20952
rect 19524 20936 19576 20942
rect 19524 20878 19576 20884
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19248 20596 19300 20602
rect 19352 20590 19472 20618
rect 19248 20538 19300 20544
rect 19260 19802 19288 20538
rect 19340 20528 19392 20534
rect 19340 20470 19392 20476
rect 19352 19922 19380 20470
rect 19340 19916 19392 19922
rect 19340 19858 19392 19864
rect 19260 19786 19380 19802
rect 18604 19780 18656 19786
rect 19260 19780 19392 19786
rect 19260 19774 19340 19780
rect 18604 19722 18656 19728
rect 19340 19722 19392 19728
rect 18512 19372 18564 19378
rect 18512 19314 18564 19320
rect 18616 19174 18644 19722
rect 19444 19666 19472 20590
rect 19892 20528 19944 20534
rect 19892 20470 19944 20476
rect 19904 19922 19932 20470
rect 19996 20398 20024 24754
rect 20076 24064 20128 24070
rect 20076 24006 20128 24012
rect 20088 23730 20116 24006
rect 20076 23724 20128 23730
rect 20076 23666 20128 23672
rect 20272 22098 20300 26948
rect 20352 26580 20404 26586
rect 20352 26522 20404 26528
rect 20364 23730 20392 26522
rect 20352 23724 20404 23730
rect 20352 23666 20404 23672
rect 20352 22976 20404 22982
rect 20352 22918 20404 22924
rect 20364 22778 20392 22918
rect 20352 22772 20404 22778
rect 20352 22714 20404 22720
rect 20260 22092 20312 22098
rect 20456 22094 20484 31726
rect 21192 29306 21220 37198
rect 21284 37126 21312 39200
rect 22572 37330 22600 39200
rect 22468 37324 22520 37330
rect 22468 37266 22520 37272
rect 22560 37324 22612 37330
rect 22560 37266 22612 37272
rect 21272 37120 21324 37126
rect 21272 37062 21324 37068
rect 22480 35894 22508 37266
rect 22928 37256 22980 37262
rect 22928 37198 22980 37204
rect 22480 35866 22600 35894
rect 21272 31884 21324 31890
rect 21272 31826 21324 31832
rect 21180 29300 21232 29306
rect 21180 29242 21232 29248
rect 21284 28506 21312 31826
rect 21548 31816 21600 31822
rect 21548 31758 21600 31764
rect 21560 29850 21588 31758
rect 21916 30592 21968 30598
rect 21916 30534 21968 30540
rect 21548 29844 21600 29850
rect 21548 29786 21600 29792
rect 21928 29034 21956 30534
rect 22100 29164 22152 29170
rect 22100 29106 22152 29112
rect 21916 29028 21968 29034
rect 21916 28970 21968 28976
rect 21192 28478 21312 28506
rect 20812 26376 20864 26382
rect 20812 26318 20864 26324
rect 20720 24744 20772 24750
rect 20720 24686 20772 24692
rect 20732 23866 20760 24686
rect 20720 23860 20772 23866
rect 20720 23802 20772 23808
rect 20824 23526 20852 26318
rect 21192 25362 21220 28478
rect 22112 27690 22140 29106
rect 21824 27668 21876 27674
rect 21824 27610 21876 27616
rect 22020 27662 22140 27690
rect 21836 25906 21864 27610
rect 21916 26988 21968 26994
rect 21916 26930 21968 26936
rect 21928 26382 21956 26930
rect 21916 26376 21968 26382
rect 21916 26318 21968 26324
rect 21824 25900 21876 25906
rect 21824 25842 21876 25848
rect 21272 25696 21324 25702
rect 21272 25638 21324 25644
rect 21180 25356 21232 25362
rect 21180 25298 21232 25304
rect 21284 25226 21312 25638
rect 21456 25356 21508 25362
rect 21456 25298 21508 25304
rect 21272 25220 21324 25226
rect 21272 25162 21324 25168
rect 20812 23520 20864 23526
rect 20812 23462 20864 23468
rect 21180 23044 21232 23050
rect 21180 22986 21232 22992
rect 21364 23044 21416 23050
rect 21364 22986 21416 22992
rect 20260 22034 20312 22040
rect 20364 22066 20484 22094
rect 20076 20936 20128 20942
rect 20076 20878 20128 20884
rect 19984 20392 20036 20398
rect 19984 20334 20036 20340
rect 20088 20210 20116 20878
rect 20168 20392 20220 20398
rect 20168 20334 20220 20340
rect 19996 20182 20116 20210
rect 19892 19916 19944 19922
rect 19892 19858 19944 19864
rect 19352 19638 19472 19666
rect 18604 19168 18656 19174
rect 18604 19110 18656 19116
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 18420 18420 18472 18426
rect 18420 18362 18472 18368
rect 18788 18284 18840 18290
rect 18788 18226 18840 18232
rect 18248 17734 18368 17762
rect 18236 17672 18288 17678
rect 18236 17614 18288 17620
rect 18248 17066 18276 17614
rect 18236 17060 18288 17066
rect 18236 17002 18288 17008
rect 18236 15632 18288 15638
rect 18236 15574 18288 15580
rect 18144 14952 18196 14958
rect 18144 14894 18196 14900
rect 18156 14249 18184 14894
rect 18248 14482 18276 15574
rect 18236 14476 18288 14482
rect 18236 14418 18288 14424
rect 18340 14362 18368 17734
rect 18420 17740 18472 17746
rect 18420 17682 18472 17688
rect 18432 17241 18460 17682
rect 18418 17232 18474 17241
rect 18418 17167 18474 17176
rect 18512 16176 18564 16182
rect 18512 16118 18564 16124
rect 18420 16040 18472 16046
rect 18420 15982 18472 15988
rect 18432 15638 18460 15982
rect 18420 15632 18472 15638
rect 18420 15574 18472 15580
rect 18340 14334 18460 14362
rect 18328 14272 18380 14278
rect 18142 14240 18198 14249
rect 18328 14214 18380 14220
rect 18142 14175 18198 14184
rect 18234 13832 18290 13841
rect 18234 13767 18290 13776
rect 18248 13530 18276 13767
rect 18236 13524 18288 13530
rect 18236 13466 18288 13472
rect 18236 12368 18288 12374
rect 18236 12310 18288 12316
rect 18248 11898 18276 12310
rect 18236 11892 18288 11898
rect 18236 11834 18288 11840
rect 18052 11212 18104 11218
rect 18052 11154 18104 11160
rect 18236 11212 18288 11218
rect 18236 11154 18288 11160
rect 17960 10736 18012 10742
rect 17960 10678 18012 10684
rect 17868 10600 17920 10606
rect 17868 10542 17920 10548
rect 17684 10464 17736 10470
rect 17684 10406 17736 10412
rect 17880 10169 17908 10542
rect 18248 10538 18276 11154
rect 18340 11082 18368 14214
rect 18432 13802 18460 14334
rect 18420 13796 18472 13802
rect 18420 13738 18472 13744
rect 18524 12442 18552 16118
rect 18696 16040 18748 16046
rect 18696 15982 18748 15988
rect 18708 15745 18736 15982
rect 18694 15736 18750 15745
rect 18694 15671 18750 15680
rect 18696 15496 18748 15502
rect 18696 15438 18748 15444
rect 18512 12436 18564 12442
rect 18512 12378 18564 12384
rect 18420 12232 18472 12238
rect 18420 12174 18472 12180
rect 18328 11076 18380 11082
rect 18328 11018 18380 11024
rect 18236 10532 18288 10538
rect 18236 10474 18288 10480
rect 18236 10192 18288 10198
rect 17866 10160 17922 10169
rect 18236 10134 18288 10140
rect 17866 10095 17868 10104
rect 17920 10095 17922 10104
rect 17868 10066 17920 10072
rect 17592 9988 17644 9994
rect 17592 9930 17644 9936
rect 17776 9648 17828 9654
rect 17776 9590 17828 9596
rect 17788 7478 17816 9590
rect 17960 8900 18012 8906
rect 17960 8842 18012 8848
rect 17972 8634 18000 8842
rect 17960 8628 18012 8634
rect 17960 8570 18012 8576
rect 17776 7472 17828 7478
rect 17776 7414 17828 7420
rect 17788 7342 17816 7414
rect 17776 7336 17828 7342
rect 17776 7278 17828 7284
rect 17500 7268 17552 7274
rect 17500 7210 17552 7216
rect 17406 7032 17462 7041
rect 17406 6967 17462 6976
rect 17512 6866 17540 7210
rect 18144 7200 18196 7206
rect 18144 7142 18196 7148
rect 17224 6860 17276 6866
rect 17224 6802 17276 6808
rect 17500 6860 17552 6866
rect 17500 6802 17552 6808
rect 16764 6452 16816 6458
rect 16764 6394 16816 6400
rect 17236 6322 17264 6802
rect 18156 6730 18184 7142
rect 18144 6724 18196 6730
rect 18144 6666 18196 6672
rect 17408 6656 17460 6662
rect 17408 6598 17460 6604
rect 17224 6316 17276 6322
rect 17224 6258 17276 6264
rect 17132 5772 17184 5778
rect 17236 5760 17264 6258
rect 17184 5732 17264 5760
rect 17132 5714 17184 5720
rect 17420 5642 17448 6598
rect 18248 5681 18276 10134
rect 18432 6089 18460 12174
rect 18602 12064 18658 12073
rect 18602 11999 18658 12008
rect 18512 11212 18564 11218
rect 18512 11154 18564 11160
rect 18524 9518 18552 11154
rect 18616 11150 18644 11999
rect 18604 11144 18656 11150
rect 18604 11086 18656 11092
rect 18604 10804 18656 10810
rect 18604 10746 18656 10752
rect 18512 9512 18564 9518
rect 18512 9454 18564 9460
rect 18418 6080 18474 6089
rect 18418 6015 18474 6024
rect 18234 5672 18290 5681
rect 17408 5636 17460 5642
rect 18234 5607 18290 5616
rect 17408 5578 17460 5584
rect 18052 5568 18104 5574
rect 18052 5510 18104 5516
rect 16948 5160 17000 5166
rect 16948 5102 17000 5108
rect 16960 4622 16988 5102
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 16948 4616 17000 4622
rect 16948 4558 17000 4564
rect 16580 4480 16632 4486
rect 16580 4422 16632 4428
rect 16592 4078 16620 4422
rect 16960 4078 16988 4558
rect 17224 4548 17276 4554
rect 17224 4490 17276 4496
rect 17236 4214 17264 4490
rect 17328 4282 17356 4626
rect 17316 4276 17368 4282
rect 17316 4218 17368 4224
rect 17224 4208 17276 4214
rect 17224 4150 17276 4156
rect 18064 4146 18092 5510
rect 18052 4140 18104 4146
rect 18052 4082 18104 4088
rect 16580 4072 16632 4078
rect 16580 4014 16632 4020
rect 16948 4072 17000 4078
rect 16948 4014 17000 4020
rect 18234 4040 18290 4049
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 16316 2746 16436 2774
rect 16316 2582 16344 2746
rect 16304 2576 16356 2582
rect 16304 2518 16356 2524
rect 16212 2304 16264 2310
rect 16212 2246 16264 2252
rect 16224 1630 16252 2246
rect 16316 1902 16344 2518
rect 16304 1896 16356 1902
rect 16304 1838 16356 1844
rect 16212 1624 16264 1630
rect 16212 1566 16264 1572
rect 16776 800 16804 3878
rect 16960 3602 16988 4014
rect 18234 3975 18236 3984
rect 18288 3975 18290 3984
rect 18236 3946 18288 3952
rect 18418 3632 18474 3641
rect 16948 3596 17000 3602
rect 18418 3567 18420 3576
rect 16948 3538 17000 3544
rect 18472 3567 18474 3576
rect 18420 3538 18472 3544
rect 16960 3058 16988 3538
rect 18512 3528 18564 3534
rect 18512 3470 18564 3476
rect 17408 3460 17460 3466
rect 17408 3402 17460 3408
rect 16948 3052 17000 3058
rect 16948 2994 17000 3000
rect 16960 2514 16988 2994
rect 17420 2854 17448 3402
rect 17408 2848 17460 2854
rect 17408 2790 17460 2796
rect 16948 2508 17000 2514
rect 16948 2450 17000 2456
rect 18524 2106 18552 3470
rect 18616 2394 18644 10746
rect 18708 8022 18736 15438
rect 18800 11218 18828 18226
rect 18880 17536 18932 17542
rect 18880 17478 18932 17484
rect 18892 17270 18920 17478
rect 18880 17264 18932 17270
rect 18880 17206 18932 17212
rect 18972 17264 19024 17270
rect 19156 17264 19208 17270
rect 18972 17206 19024 17212
rect 19076 17224 19156 17252
rect 18984 16794 19012 17206
rect 18972 16788 19024 16794
rect 18972 16730 19024 16736
rect 18972 15020 19024 15026
rect 18972 14962 19024 14968
rect 18984 14414 19012 14962
rect 18972 14408 19024 14414
rect 18972 14350 19024 14356
rect 18878 12472 18934 12481
rect 18878 12407 18934 12416
rect 18892 11626 18920 12407
rect 18972 11824 19024 11830
rect 18972 11766 19024 11772
rect 18880 11620 18932 11626
rect 18880 11562 18932 11568
rect 18984 11558 19012 11766
rect 18972 11552 19024 11558
rect 18972 11494 19024 11500
rect 18880 11280 18932 11286
rect 18880 11222 18932 11228
rect 18788 11212 18840 11218
rect 18788 11154 18840 11160
rect 18788 10600 18840 10606
rect 18788 10542 18840 10548
rect 18800 9625 18828 10542
rect 18786 9616 18842 9625
rect 18786 9551 18842 9560
rect 18696 8016 18748 8022
rect 18696 7958 18748 7964
rect 18892 7562 18920 11222
rect 18972 10124 19024 10130
rect 18972 10066 19024 10072
rect 18984 9926 19012 10066
rect 18972 9920 19024 9926
rect 18972 9862 19024 9868
rect 18984 9518 19012 9862
rect 18972 9512 19024 9518
rect 18972 9454 19024 9460
rect 19076 8090 19104 17224
rect 19156 17206 19208 17212
rect 19352 15609 19380 19638
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19432 19508 19484 19514
rect 19432 19450 19484 19456
rect 19444 17252 19472 19450
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19996 17649 20024 20182
rect 20180 19786 20208 20334
rect 20168 19780 20220 19786
rect 20168 19722 20220 19728
rect 20180 17762 20208 19722
rect 20260 18760 20312 18766
rect 20258 18728 20260 18737
rect 20312 18728 20314 18737
rect 20258 18663 20314 18672
rect 20272 18426 20300 18663
rect 20260 18420 20312 18426
rect 20260 18362 20312 18368
rect 20364 18358 20392 22066
rect 20904 22024 20956 22030
rect 20904 21966 20956 21972
rect 20916 21554 20944 21966
rect 20904 21548 20956 21554
rect 20904 21490 20956 21496
rect 21088 21548 21140 21554
rect 21088 21490 21140 21496
rect 20444 21344 20496 21350
rect 20444 21286 20496 21292
rect 20456 20874 20484 21286
rect 20444 20868 20496 20874
rect 20444 20810 20496 20816
rect 20628 19304 20680 19310
rect 20628 19246 20680 19252
rect 20444 19236 20496 19242
rect 20444 19178 20496 19184
rect 20352 18352 20404 18358
rect 20352 18294 20404 18300
rect 20180 17734 20392 17762
rect 20168 17672 20220 17678
rect 19982 17640 20038 17649
rect 20168 17614 20220 17620
rect 19982 17575 20038 17584
rect 19984 17536 20036 17542
rect 19984 17478 20036 17484
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19444 17224 19564 17252
rect 19536 16697 19564 17224
rect 19616 17128 19668 17134
rect 19614 17096 19616 17105
rect 19668 17096 19670 17105
rect 19614 17031 19670 17040
rect 19522 16688 19578 16697
rect 19522 16623 19578 16632
rect 19536 16522 19564 16623
rect 19996 16522 20024 17478
rect 20076 16992 20128 16998
rect 20076 16934 20128 16940
rect 19524 16516 19576 16522
rect 19524 16458 19576 16464
rect 19984 16516 20036 16522
rect 19984 16458 20036 16464
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19984 16244 20036 16250
rect 19984 16186 20036 16192
rect 19338 15600 19394 15609
rect 19996 15570 20024 16186
rect 20088 16182 20116 16934
rect 20076 16176 20128 16182
rect 20076 16118 20128 16124
rect 20076 15972 20128 15978
rect 20076 15914 20128 15920
rect 19338 15535 19394 15544
rect 19984 15564 20036 15570
rect 19984 15506 20036 15512
rect 19340 15496 19392 15502
rect 19340 15438 19392 15444
rect 19522 15464 19578 15473
rect 19156 14272 19208 14278
rect 19156 14214 19208 14220
rect 19168 9654 19196 14214
rect 19352 14090 19380 15438
rect 19522 15399 19578 15408
rect 19536 15366 19564 15399
rect 19524 15360 19576 15366
rect 19524 15302 19576 15308
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19524 15156 19576 15162
rect 19524 15098 19576 15104
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 19444 14618 19472 14758
rect 19536 14657 19564 15098
rect 19996 14958 20024 15506
rect 20088 15434 20116 15914
rect 20076 15428 20128 15434
rect 20076 15370 20128 15376
rect 20076 15156 20128 15162
rect 20076 15098 20128 15104
rect 20088 15065 20116 15098
rect 20074 15056 20130 15065
rect 20074 14991 20130 15000
rect 20088 14958 20116 14991
rect 19984 14952 20036 14958
rect 19984 14894 20036 14900
rect 20076 14952 20128 14958
rect 20076 14894 20128 14900
rect 19522 14648 19578 14657
rect 19432 14612 19484 14618
rect 19522 14583 19578 14592
rect 19432 14554 19484 14560
rect 19984 14272 20036 14278
rect 19984 14214 20036 14220
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19260 14062 19380 14090
rect 19996 14074 20024 14214
rect 19984 14068 20036 14074
rect 19260 12730 19288 14062
rect 19984 14010 20036 14016
rect 20076 14068 20128 14074
rect 20076 14010 20128 14016
rect 19340 14000 19392 14006
rect 19340 13942 19392 13948
rect 19352 13326 19380 13942
rect 19708 13524 19760 13530
rect 19708 13466 19760 13472
rect 19340 13320 19392 13326
rect 19720 13297 19748 13466
rect 19340 13262 19392 13268
rect 19706 13288 19762 13297
rect 19352 12850 19380 13262
rect 19706 13223 19708 13232
rect 19760 13223 19762 13232
rect 19708 13194 19760 13200
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19982 13016 20038 13025
rect 19524 12980 19576 12986
rect 19982 12951 19984 12960
rect 19524 12922 19576 12928
rect 20036 12951 20038 12960
rect 19984 12922 20036 12928
rect 19340 12844 19392 12850
rect 19392 12804 19472 12832
rect 19340 12786 19392 12792
rect 19260 12702 19380 12730
rect 19352 12186 19380 12702
rect 19444 12306 19472 12804
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 19260 12158 19380 12186
rect 19260 11778 19288 12158
rect 19340 12096 19392 12102
rect 19340 12038 19392 12044
rect 19352 11898 19380 12038
rect 19340 11892 19392 11898
rect 19340 11834 19392 11840
rect 19260 11750 19380 11778
rect 19444 11762 19472 12242
rect 19536 12102 19564 12922
rect 19984 12164 20036 12170
rect 19984 12106 20036 12112
rect 19524 12096 19576 12102
rect 19524 12038 19576 12044
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19248 11212 19300 11218
rect 19248 11154 19300 11160
rect 19260 10674 19288 11154
rect 19352 10810 19380 11750
rect 19432 11756 19484 11762
rect 19432 11698 19484 11704
rect 19444 11218 19472 11698
rect 19432 11212 19484 11218
rect 19432 11154 19484 11160
rect 19432 11076 19484 11082
rect 19432 11018 19484 11024
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 19248 10668 19300 10674
rect 19248 10610 19300 10616
rect 19340 10056 19392 10062
rect 19340 9998 19392 10004
rect 19156 9648 19208 9654
rect 19156 9590 19208 9596
rect 19352 9518 19380 9998
rect 19340 9512 19392 9518
rect 19340 9454 19392 9460
rect 19248 9376 19300 9382
rect 19248 9318 19300 9324
rect 19260 8974 19288 9318
rect 19352 9042 19380 9454
rect 19340 9036 19392 9042
rect 19340 8978 19392 8984
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 19064 8084 19116 8090
rect 19064 8026 19116 8032
rect 18892 7534 19012 7562
rect 18880 7404 18932 7410
rect 18880 7346 18932 7352
rect 18892 7002 18920 7346
rect 18880 6996 18932 7002
rect 18880 6938 18932 6944
rect 18984 5778 19012 7534
rect 19076 6458 19104 8026
rect 19064 6452 19116 6458
rect 19064 6394 19116 6400
rect 18972 5772 19024 5778
rect 18972 5714 19024 5720
rect 18984 5574 19012 5714
rect 18972 5568 19024 5574
rect 18972 5510 19024 5516
rect 18880 5228 18932 5234
rect 18880 5170 18932 5176
rect 18788 5024 18840 5030
rect 18788 4966 18840 4972
rect 18800 4826 18828 4966
rect 18788 4820 18840 4826
rect 18788 4762 18840 4768
rect 18892 4486 18920 5170
rect 19260 4690 19288 8910
rect 19352 8566 19380 8978
rect 19444 8906 19472 11018
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19996 10742 20024 12106
rect 19984 10736 20036 10742
rect 19984 10678 20036 10684
rect 19616 10600 19668 10606
rect 19616 10542 19668 10548
rect 19628 10198 19656 10542
rect 19616 10192 19668 10198
rect 19616 10134 19668 10140
rect 19984 9988 20036 9994
rect 19984 9930 20036 9936
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19432 8900 19484 8906
rect 19432 8842 19484 8848
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19340 8560 19392 8566
rect 19340 8502 19392 8508
rect 19996 8276 20024 9930
rect 20088 8430 20116 14010
rect 20180 10130 20208 17614
rect 20260 17536 20312 17542
rect 20260 17478 20312 17484
rect 20272 17338 20300 17478
rect 20260 17332 20312 17338
rect 20260 17274 20312 17280
rect 20260 17196 20312 17202
rect 20260 17138 20312 17144
rect 20272 16522 20300 17138
rect 20260 16516 20312 16522
rect 20260 16458 20312 16464
rect 20364 16182 20392 17734
rect 20352 16176 20404 16182
rect 20352 16118 20404 16124
rect 20456 15858 20484 19178
rect 20536 19168 20588 19174
rect 20536 19110 20588 19116
rect 20548 18442 20576 19110
rect 20640 18970 20668 19246
rect 20628 18964 20680 18970
rect 20628 18906 20680 18912
rect 20548 18414 20668 18442
rect 20536 18284 20588 18290
rect 20536 18226 20588 18232
rect 20548 18057 20576 18226
rect 20534 18048 20590 18057
rect 20534 17983 20590 17992
rect 20536 17060 20588 17066
rect 20536 17002 20588 17008
rect 20548 15978 20576 17002
rect 20536 15972 20588 15978
rect 20536 15914 20588 15920
rect 20272 15830 20484 15858
rect 20272 10810 20300 15830
rect 20640 15722 20668 18414
rect 20812 17128 20864 17134
rect 20718 17096 20774 17105
rect 20812 17070 20864 17076
rect 20718 17031 20774 17040
rect 20732 16590 20760 17031
rect 20720 16584 20772 16590
rect 20824 16561 20852 17070
rect 20720 16526 20772 16532
rect 20810 16552 20866 16561
rect 20810 16487 20866 16496
rect 20720 16176 20772 16182
rect 20720 16118 20772 16124
rect 20364 15694 20668 15722
rect 20364 14074 20392 15694
rect 20628 15632 20680 15638
rect 20628 15574 20680 15580
rect 20444 15564 20496 15570
rect 20444 15506 20496 15512
rect 20456 14822 20484 15506
rect 20534 15464 20590 15473
rect 20534 15399 20590 15408
rect 20548 15094 20576 15399
rect 20640 15201 20668 15574
rect 20732 15570 20760 16118
rect 20720 15564 20772 15570
rect 20720 15506 20772 15512
rect 20626 15192 20682 15201
rect 20626 15127 20682 15136
rect 20536 15088 20588 15094
rect 20536 15030 20588 15036
rect 20536 14952 20588 14958
rect 20536 14894 20588 14900
rect 20444 14816 20496 14822
rect 20444 14758 20496 14764
rect 20548 14618 20576 14894
rect 20536 14612 20588 14618
rect 20536 14554 20588 14560
rect 20442 14512 20498 14521
rect 20442 14447 20498 14456
rect 20456 14414 20484 14447
rect 20444 14408 20496 14414
rect 20444 14350 20496 14356
rect 20442 14240 20498 14249
rect 20442 14175 20498 14184
rect 20352 14068 20404 14074
rect 20352 14010 20404 14016
rect 20352 13728 20404 13734
rect 20352 13670 20404 13676
rect 20364 12782 20392 13670
rect 20352 12776 20404 12782
rect 20352 12718 20404 12724
rect 20456 10810 20484 14175
rect 20536 13864 20588 13870
rect 20536 13806 20588 13812
rect 20260 10804 20312 10810
rect 20260 10746 20312 10752
rect 20444 10804 20496 10810
rect 20444 10746 20496 10752
rect 20548 10130 20576 13806
rect 20720 12776 20772 12782
rect 20720 12718 20772 12724
rect 20626 12336 20682 12345
rect 20626 12271 20682 12280
rect 20168 10124 20220 10130
rect 20168 10066 20220 10072
rect 20536 10124 20588 10130
rect 20536 10066 20588 10072
rect 20168 9988 20220 9994
rect 20168 9930 20220 9936
rect 20076 8424 20128 8430
rect 20076 8366 20128 8372
rect 19996 8248 20116 8276
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19996 7546 20024 7822
rect 19984 7540 20036 7546
rect 19984 7482 20036 7488
rect 19982 7440 20038 7449
rect 19708 7404 19760 7410
rect 19982 7375 20038 7384
rect 19708 7346 19760 7352
rect 19616 7336 19668 7342
rect 19614 7304 19616 7313
rect 19668 7304 19670 7313
rect 19614 7239 19670 7248
rect 19720 6866 19748 7346
rect 19432 6860 19484 6866
rect 19432 6802 19484 6808
rect 19708 6860 19760 6866
rect 19708 6802 19760 6808
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19352 6322 19380 6394
rect 19444 6322 19472 6802
rect 19616 6792 19668 6798
rect 19614 6760 19616 6769
rect 19668 6760 19670 6769
rect 19996 6730 20024 7375
rect 20088 7018 20116 8248
rect 20180 7206 20208 9930
rect 20272 9166 20484 9194
rect 20272 9042 20300 9166
rect 20260 9036 20312 9042
rect 20260 8978 20312 8984
rect 20352 9036 20404 9042
rect 20352 8978 20404 8984
rect 20364 8294 20392 8978
rect 20456 8362 20484 9166
rect 20640 8922 20668 12271
rect 20732 9518 20760 12718
rect 20720 9512 20772 9518
rect 20720 9454 20772 9460
rect 20548 8894 20668 8922
rect 20718 8936 20774 8945
rect 20444 8356 20496 8362
rect 20444 8298 20496 8304
rect 20352 8288 20404 8294
rect 20352 8230 20404 8236
rect 20364 7342 20392 8230
rect 20352 7336 20404 7342
rect 20352 7278 20404 7284
rect 20168 7200 20220 7206
rect 20168 7142 20220 7148
rect 20088 6990 20208 7018
rect 19614 6695 19670 6704
rect 19984 6724 20036 6730
rect 19984 6666 20036 6672
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19706 6352 19762 6361
rect 19340 6316 19392 6322
rect 19340 6258 19392 6264
rect 19432 6316 19484 6322
rect 19706 6287 19762 6296
rect 19432 6258 19484 6264
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 19352 5166 19380 6054
rect 19444 5778 19472 6258
rect 19720 6186 19748 6287
rect 19708 6180 19760 6186
rect 19708 6122 19760 6128
rect 19432 5772 19484 5778
rect 19432 5714 19484 5720
rect 19444 5234 19472 5714
rect 20074 5536 20130 5545
rect 19574 5468 19882 5477
rect 20074 5471 20130 5480
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 20088 5370 20116 5471
rect 20180 5386 20208 6990
rect 20260 6452 20312 6458
rect 20260 6394 20312 6400
rect 20272 5930 20300 6394
rect 20548 5930 20576 8894
rect 20718 8871 20774 8880
rect 20732 8838 20760 8871
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 20720 8832 20772 8838
rect 20720 8774 20772 8780
rect 20640 7342 20668 8774
rect 20628 7336 20680 7342
rect 20628 7278 20680 7284
rect 20824 6769 20852 16487
rect 20916 12442 20944 21490
rect 20996 21412 21048 21418
rect 20996 21354 21048 21360
rect 21008 20942 21036 21354
rect 20996 20936 21048 20942
rect 20996 20878 21048 20884
rect 20996 20392 21048 20398
rect 20996 20334 21048 20340
rect 21008 13802 21036 20334
rect 21100 19378 21128 21490
rect 21088 19372 21140 19378
rect 21088 19314 21140 19320
rect 21088 18080 21140 18086
rect 21088 18022 21140 18028
rect 21100 17882 21128 18022
rect 21192 17882 21220 22986
rect 21376 22574 21404 22986
rect 21364 22568 21416 22574
rect 21364 22510 21416 22516
rect 21272 21004 21324 21010
rect 21272 20946 21324 20952
rect 21284 19922 21312 20946
rect 21364 20528 21416 20534
rect 21364 20470 21416 20476
rect 21272 19916 21324 19922
rect 21272 19858 21324 19864
rect 21376 19378 21404 20470
rect 21364 19372 21416 19378
rect 21364 19314 21416 19320
rect 21088 17876 21140 17882
rect 21088 17818 21140 17824
rect 21180 17876 21232 17882
rect 21180 17818 21232 17824
rect 21364 17808 21416 17814
rect 21364 17750 21416 17756
rect 21088 16448 21140 16454
rect 21088 16390 21140 16396
rect 21100 16114 21128 16390
rect 21088 16108 21140 16114
rect 21088 16050 21140 16056
rect 21180 15360 21232 15366
rect 21180 15302 21232 15308
rect 21088 14816 21140 14822
rect 21088 14758 21140 14764
rect 20996 13796 21048 13802
rect 20996 13738 21048 13744
rect 21100 13394 21128 14758
rect 21088 13388 21140 13394
rect 21088 13330 21140 13336
rect 20904 12436 20956 12442
rect 20904 12378 20956 12384
rect 21192 11830 21220 15302
rect 21272 14340 21324 14346
rect 21272 14282 21324 14288
rect 21284 13138 21312 14282
rect 21376 13240 21404 17750
rect 21468 14958 21496 25298
rect 21640 23792 21692 23798
rect 21640 23734 21692 23740
rect 21652 20398 21680 23734
rect 21640 20392 21692 20398
rect 21640 20334 21692 20340
rect 21548 20256 21600 20262
rect 21548 20198 21600 20204
rect 21560 19718 21588 20198
rect 21640 19780 21692 19786
rect 21640 19722 21692 19728
rect 21548 19712 21600 19718
rect 21548 19654 21600 19660
rect 21652 17762 21680 19722
rect 21732 19372 21784 19378
rect 21732 19314 21784 19320
rect 21560 17734 21680 17762
rect 21456 14952 21508 14958
rect 21456 14894 21508 14900
rect 21560 14498 21588 17734
rect 21640 17672 21692 17678
rect 21640 17614 21692 17620
rect 21468 14470 21588 14498
rect 21468 13734 21496 14470
rect 21548 14340 21600 14346
rect 21548 14282 21600 14288
rect 21560 14074 21588 14282
rect 21548 14068 21600 14074
rect 21548 14010 21600 14016
rect 21456 13728 21508 13734
rect 21456 13670 21508 13676
rect 21652 13326 21680 17614
rect 21640 13320 21692 13326
rect 21640 13262 21692 13268
rect 21376 13212 21588 13240
rect 21284 13110 21496 13138
rect 21272 12708 21324 12714
rect 21272 12650 21324 12656
rect 21180 11824 21232 11830
rect 21180 11766 21232 11772
rect 21088 11756 21140 11762
rect 21088 11698 21140 11704
rect 21100 9518 21128 11698
rect 21088 9512 21140 9518
rect 21088 9454 21140 9460
rect 20904 9376 20956 9382
rect 20904 9318 20956 9324
rect 20916 9110 20944 9318
rect 20904 9104 20956 9110
rect 20904 9046 20956 9052
rect 21180 8900 21232 8906
rect 21180 8842 21232 8848
rect 21192 8634 21220 8842
rect 21180 8628 21232 8634
rect 21180 8570 21232 8576
rect 20996 8560 21048 8566
rect 20996 8502 21048 8508
rect 21008 8090 21036 8502
rect 21284 8362 21312 12650
rect 21468 12374 21496 13110
rect 21560 12481 21588 13212
rect 21652 12646 21680 13262
rect 21744 12714 21772 19314
rect 21836 14482 21864 25842
rect 21928 24818 21956 26318
rect 21916 24812 21968 24818
rect 21916 24754 21968 24760
rect 21928 23798 21956 24754
rect 21916 23792 21968 23798
rect 21916 23734 21968 23740
rect 21916 22976 21968 22982
rect 21916 22918 21968 22924
rect 21928 17882 21956 22918
rect 22020 21185 22048 27662
rect 22468 26240 22520 26246
rect 22468 26182 22520 26188
rect 22192 25832 22244 25838
rect 22192 25774 22244 25780
rect 22204 24954 22232 25774
rect 22480 25294 22508 26182
rect 22468 25288 22520 25294
rect 22468 25230 22520 25236
rect 22192 24948 22244 24954
rect 22192 24890 22244 24896
rect 22100 24268 22152 24274
rect 22100 24210 22152 24216
rect 22112 23662 22140 24210
rect 22192 23792 22244 23798
rect 22192 23734 22244 23740
rect 22100 23656 22152 23662
rect 22100 23598 22152 23604
rect 22204 22778 22232 23734
rect 22376 23656 22428 23662
rect 22376 23598 22428 23604
rect 22388 22982 22416 23598
rect 22376 22976 22428 22982
rect 22376 22918 22428 22924
rect 22192 22772 22244 22778
rect 22192 22714 22244 22720
rect 22388 21962 22416 22918
rect 22572 22094 22600 35866
rect 22940 25770 22968 37198
rect 23216 36922 23244 39200
rect 24504 37262 24532 39200
rect 25792 37262 25820 39200
rect 24492 37256 24544 37262
rect 24492 37198 24544 37204
rect 25780 37256 25832 37262
rect 25780 37198 25832 37204
rect 25504 37188 25556 37194
rect 25504 37130 25556 37136
rect 24584 37120 24636 37126
rect 24584 37062 24636 37068
rect 23204 36916 23256 36922
rect 23204 36858 23256 36864
rect 23296 36780 23348 36786
rect 23296 36722 23348 36728
rect 23308 32026 23336 36722
rect 23296 32020 23348 32026
rect 23296 31962 23348 31968
rect 23204 31952 23256 31958
rect 23204 31894 23256 31900
rect 23112 26240 23164 26246
rect 23112 26182 23164 26188
rect 23124 25906 23152 26182
rect 23112 25900 23164 25906
rect 23112 25842 23164 25848
rect 22928 25764 22980 25770
rect 22928 25706 22980 25712
rect 22928 24880 22980 24886
rect 22928 24822 22980 24828
rect 22940 24614 22968 24822
rect 22836 24608 22888 24614
rect 22836 24550 22888 24556
rect 22928 24608 22980 24614
rect 22928 24550 22980 24556
rect 22848 23866 22876 24550
rect 23112 24404 23164 24410
rect 23112 24346 23164 24352
rect 22836 23860 22888 23866
rect 22836 23802 22888 23808
rect 22480 22066 22600 22094
rect 22376 21956 22428 21962
rect 22376 21898 22428 21904
rect 22006 21176 22062 21185
rect 22006 21111 22062 21120
rect 21916 17876 21968 17882
rect 21916 17818 21968 17824
rect 22020 17082 22048 21111
rect 22480 20942 22508 22066
rect 22836 21956 22888 21962
rect 22836 21898 22888 21904
rect 22848 21350 22876 21898
rect 22836 21344 22888 21350
rect 22836 21286 22888 21292
rect 22744 21140 22796 21146
rect 22744 21082 22796 21088
rect 22756 21049 22784 21082
rect 22928 21072 22980 21078
rect 22742 21040 22798 21049
rect 22928 21014 22980 21020
rect 22742 20975 22798 20984
rect 22468 20936 22520 20942
rect 22468 20878 22520 20884
rect 22560 20936 22612 20942
rect 22560 20878 22612 20884
rect 22572 20398 22600 20878
rect 22940 20874 22968 21014
rect 22928 20868 22980 20874
rect 22928 20810 22980 20816
rect 23020 20528 23072 20534
rect 23020 20470 23072 20476
rect 22560 20392 22612 20398
rect 22560 20334 22612 20340
rect 22284 20052 22336 20058
rect 22284 19994 22336 20000
rect 22296 19922 22324 19994
rect 22744 19984 22796 19990
rect 22744 19926 22796 19932
rect 22100 19916 22152 19922
rect 22100 19858 22152 19864
rect 22284 19916 22336 19922
rect 22284 19858 22336 19864
rect 21928 17054 22048 17082
rect 22112 17082 22140 19858
rect 22560 19440 22612 19446
rect 22560 19382 22612 19388
rect 22376 18352 22428 18358
rect 22376 18294 22428 18300
rect 22192 17536 22244 17542
rect 22192 17478 22244 17484
rect 22204 17270 22232 17478
rect 22192 17264 22244 17270
rect 22192 17206 22244 17212
rect 22284 17264 22336 17270
rect 22284 17206 22336 17212
rect 22112 17054 22232 17082
rect 21928 16114 21956 17054
rect 21916 16108 21968 16114
rect 21916 16050 21968 16056
rect 22100 16040 22152 16046
rect 22100 15982 22152 15988
rect 22112 15910 22140 15982
rect 22100 15904 22152 15910
rect 22100 15846 22152 15852
rect 22112 15570 22140 15846
rect 22100 15564 22152 15570
rect 22100 15506 22152 15512
rect 22008 15496 22060 15502
rect 22008 15438 22060 15444
rect 21916 14952 21968 14958
rect 21916 14894 21968 14900
rect 21824 14476 21876 14482
rect 21824 14418 21876 14424
rect 21928 14074 21956 14894
rect 22020 14618 22048 15438
rect 22008 14612 22060 14618
rect 22008 14554 22060 14560
rect 21916 14068 21968 14074
rect 21916 14010 21968 14016
rect 21824 14000 21876 14006
rect 21824 13942 21876 13948
rect 21836 13530 21864 13942
rect 21916 13796 21968 13802
rect 21916 13738 21968 13744
rect 21824 13524 21876 13530
rect 21824 13466 21876 13472
rect 21824 13252 21876 13258
rect 21824 13194 21876 13200
rect 21732 12708 21784 12714
rect 21732 12650 21784 12656
rect 21640 12640 21692 12646
rect 21640 12582 21692 12588
rect 21546 12472 21602 12481
rect 21546 12407 21602 12416
rect 21732 12436 21784 12442
rect 21732 12378 21784 12384
rect 21456 12368 21508 12374
rect 21456 12310 21508 12316
rect 21548 12300 21600 12306
rect 21548 12242 21600 12248
rect 21560 11218 21588 12242
rect 21640 12232 21692 12238
rect 21640 12174 21692 12180
rect 21548 11212 21600 11218
rect 21548 11154 21600 11160
rect 21364 9172 21416 9178
rect 21364 9114 21416 9120
rect 21376 8498 21404 9114
rect 21364 8492 21416 8498
rect 21364 8434 21416 8440
rect 21272 8356 21324 8362
rect 21272 8298 21324 8304
rect 20996 8084 21048 8090
rect 20996 8026 21048 8032
rect 21284 7750 21312 8298
rect 21560 8022 21588 11154
rect 21548 8016 21600 8022
rect 21548 7958 21600 7964
rect 21272 7744 21324 7750
rect 21272 7686 21324 7692
rect 21548 7744 21600 7750
rect 21548 7686 21600 7692
rect 21364 7472 21416 7478
rect 21364 7414 21416 7420
rect 21086 7304 21142 7313
rect 20996 7268 21048 7274
rect 21086 7239 21142 7248
rect 20996 7210 21048 7216
rect 20810 6760 20866 6769
rect 20810 6695 20866 6704
rect 20272 5902 20576 5930
rect 20364 5642 20392 5902
rect 20352 5636 20404 5642
rect 20352 5578 20404 5584
rect 20534 5400 20590 5409
rect 20076 5364 20128 5370
rect 20180 5358 20534 5386
rect 20534 5335 20590 5344
rect 20076 5306 20128 5312
rect 19432 5228 19484 5234
rect 19432 5170 19484 5176
rect 19340 5160 19392 5166
rect 19340 5102 19392 5108
rect 19248 4684 19300 4690
rect 19248 4626 19300 4632
rect 19156 4616 19208 4622
rect 19156 4558 19208 4564
rect 18696 4480 18748 4486
rect 18696 4422 18748 4428
rect 18880 4480 18932 4486
rect 18880 4422 18932 4428
rect 18708 4078 18736 4422
rect 18880 4208 18932 4214
rect 18878 4176 18880 4185
rect 18932 4176 18934 4185
rect 18878 4111 18934 4120
rect 18696 4072 18748 4078
rect 18696 4014 18748 4020
rect 19168 3942 19196 4558
rect 19352 4026 19380 5102
rect 19524 5092 19576 5098
rect 19524 5034 19576 5040
rect 19536 4865 19564 5034
rect 19522 4856 19578 4865
rect 19522 4791 19578 4800
rect 19984 4480 20036 4486
rect 19984 4422 20036 4428
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19260 3998 19380 4026
rect 19156 3936 19208 3942
rect 19156 3878 19208 3884
rect 19168 3602 19196 3878
rect 19260 3754 19288 3998
rect 19996 3942 20024 4422
rect 20258 4312 20314 4321
rect 20258 4247 20314 4256
rect 19984 3936 20036 3942
rect 19984 3878 20036 3884
rect 20074 3904 20130 3913
rect 19996 3777 20024 3878
rect 20074 3839 20130 3848
rect 19338 3768 19394 3777
rect 19260 3726 19338 3754
rect 19338 3703 19394 3712
rect 19982 3768 20038 3777
rect 19982 3703 20038 3712
rect 19352 3641 19564 3652
rect 19338 3632 19578 3641
rect 19156 3596 19208 3602
rect 19394 3624 19522 3632
rect 19338 3567 19394 3576
rect 19522 3567 19578 3576
rect 19156 3538 19208 3544
rect 18788 3392 18840 3398
rect 18788 3334 18840 3340
rect 18616 2366 18736 2394
rect 18708 2310 18736 2366
rect 18696 2304 18748 2310
rect 18696 2246 18748 2252
rect 18052 2100 18104 2106
rect 18052 2042 18104 2048
rect 18512 2100 18564 2106
rect 18512 2042 18564 2048
rect 18064 800 18092 2042
rect 18800 1698 18828 3334
rect 19168 3126 19196 3538
rect 19292 3496 19348 3505
rect 19614 3496 19670 3505
rect 19348 3454 19614 3482
rect 19292 3431 19348 3440
rect 19614 3431 19670 3440
rect 19340 3392 19392 3398
rect 19306 3340 19340 3346
rect 19306 3334 19392 3340
rect 19306 3318 19380 3334
rect 19064 3120 19116 3126
rect 19064 3062 19116 3068
rect 19156 3120 19208 3126
rect 19156 3062 19208 3068
rect 18972 3052 19024 3058
rect 18972 2994 19024 3000
rect 18984 2582 19012 2994
rect 18972 2576 19024 2582
rect 18972 2518 19024 2524
rect 19076 2038 19104 3062
rect 19156 2984 19208 2990
rect 19306 2972 19334 3318
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19614 3088 19670 3097
rect 19614 3023 19670 3032
rect 19524 2984 19576 2990
rect 19306 2944 19524 2972
rect 19156 2926 19208 2932
rect 19524 2926 19576 2932
rect 19168 2310 19196 2926
rect 19260 2774 19564 2802
rect 19260 2514 19288 2774
rect 19338 2544 19394 2553
rect 19248 2508 19300 2514
rect 19338 2479 19394 2488
rect 19248 2450 19300 2456
rect 19156 2304 19208 2310
rect 19156 2246 19208 2252
rect 19064 2032 19116 2038
rect 19064 1974 19116 1980
rect 18788 1692 18840 1698
rect 18788 1634 18840 1640
rect 19352 800 19380 2479
rect 19536 2417 19564 2774
rect 19628 2553 19656 3023
rect 20088 2854 20116 3839
rect 20076 2848 20128 2854
rect 20272 2825 20300 4247
rect 20548 4146 20576 5335
rect 20904 5024 20956 5030
rect 20904 4966 20956 4972
rect 20720 4480 20772 4486
rect 20720 4422 20772 4428
rect 20812 4480 20864 4486
rect 20812 4422 20864 4428
rect 20732 4146 20760 4422
rect 20536 4140 20588 4146
rect 20536 4082 20588 4088
rect 20720 4140 20772 4146
rect 20720 4082 20772 4088
rect 20824 4078 20852 4422
rect 20812 4072 20864 4078
rect 20812 4014 20864 4020
rect 20916 3670 20944 4966
rect 21008 4185 21036 7210
rect 21100 7206 21128 7239
rect 21088 7200 21140 7206
rect 21088 7142 21140 7148
rect 21180 6860 21232 6866
rect 21180 6802 21232 6808
rect 21192 6769 21220 6802
rect 21272 6792 21324 6798
rect 21178 6760 21234 6769
rect 21272 6734 21324 6740
rect 21178 6695 21234 6704
rect 21284 6361 21312 6734
rect 21270 6352 21326 6361
rect 21270 6287 21326 6296
rect 21178 6080 21234 6089
rect 21178 6015 21234 6024
rect 21192 4554 21220 6015
rect 21272 5160 21324 5166
rect 21272 5102 21324 5108
rect 21284 4758 21312 5102
rect 21272 4752 21324 4758
rect 21272 4694 21324 4700
rect 21180 4548 21232 4554
rect 21180 4490 21232 4496
rect 20994 4176 21050 4185
rect 21376 4146 21404 7414
rect 21560 6934 21588 7686
rect 21548 6928 21600 6934
rect 21548 6870 21600 6876
rect 21546 6760 21602 6769
rect 21546 6695 21548 6704
rect 21600 6695 21602 6704
rect 21548 6666 21600 6672
rect 21652 6186 21680 12174
rect 21744 8974 21772 12378
rect 21836 10690 21864 13194
rect 21928 12306 21956 13738
rect 22020 12850 22048 14554
rect 22100 13932 22152 13938
rect 22100 13874 22152 13880
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 21916 12300 21968 12306
rect 21916 12242 21968 12248
rect 22020 11082 22048 12786
rect 22112 12442 22140 13874
rect 22100 12436 22152 12442
rect 22100 12378 22152 12384
rect 22100 12300 22152 12306
rect 22100 12242 22152 12248
rect 22112 12209 22140 12242
rect 22098 12200 22154 12209
rect 22098 12135 22154 12144
rect 22100 12096 22152 12102
rect 22100 12038 22152 12044
rect 22112 11354 22140 12038
rect 22100 11348 22152 11354
rect 22100 11290 22152 11296
rect 22008 11076 22060 11082
rect 22008 11018 22060 11024
rect 21836 10662 21956 10690
rect 21824 10600 21876 10606
rect 21824 10542 21876 10548
rect 21836 10130 21864 10542
rect 21928 10470 21956 10662
rect 21916 10464 21968 10470
rect 21916 10406 21968 10412
rect 21824 10124 21876 10130
rect 21824 10066 21876 10072
rect 21732 8968 21784 8974
rect 21732 8910 21784 8916
rect 21824 8832 21876 8838
rect 21824 8774 21876 8780
rect 21836 8022 21864 8774
rect 21824 8016 21876 8022
rect 21824 7958 21876 7964
rect 22008 7812 22060 7818
rect 22008 7754 22060 7760
rect 21916 7268 21968 7274
rect 21916 7210 21968 7216
rect 21822 6488 21878 6497
rect 21822 6423 21878 6432
rect 21640 6180 21692 6186
rect 21640 6122 21692 6128
rect 21456 5704 21508 5710
rect 21456 5646 21508 5652
rect 21546 5672 21602 5681
rect 21468 4457 21496 5646
rect 21546 5607 21602 5616
rect 21560 5574 21588 5607
rect 21548 5568 21600 5574
rect 21548 5510 21600 5516
rect 21652 5386 21680 6122
rect 21730 5536 21786 5545
rect 21730 5471 21786 5480
rect 21560 5358 21680 5386
rect 21560 4554 21588 5358
rect 21744 5302 21772 5471
rect 21640 5296 21692 5302
rect 21640 5238 21692 5244
rect 21732 5296 21784 5302
rect 21732 5238 21784 5244
rect 21548 4548 21600 4554
rect 21548 4490 21600 4496
rect 21454 4448 21510 4457
rect 21454 4383 21510 4392
rect 21652 4185 21680 5238
rect 21732 4616 21784 4622
rect 21732 4558 21784 4564
rect 21454 4176 21510 4185
rect 20994 4111 21050 4120
rect 21088 4140 21140 4146
rect 21088 4082 21140 4088
rect 21364 4140 21416 4146
rect 21454 4111 21510 4120
rect 21638 4176 21694 4185
rect 21638 4111 21694 4120
rect 21364 4082 21416 4088
rect 21100 4010 21128 4082
rect 21088 4004 21140 4010
rect 21088 3946 21140 3952
rect 20904 3664 20956 3670
rect 20534 3632 20590 3641
rect 20904 3606 20956 3612
rect 20534 3567 20590 3576
rect 20548 2990 20576 3567
rect 21468 3466 21496 4111
rect 21456 3460 21508 3466
rect 21456 3402 21508 3408
rect 21744 3058 21772 4558
rect 21836 4049 21864 6423
rect 21928 6118 21956 7210
rect 22020 6866 22048 7754
rect 22008 6860 22060 6866
rect 22008 6802 22060 6808
rect 22204 6662 22232 17054
rect 22296 16522 22324 17206
rect 22284 16516 22336 16522
rect 22284 16458 22336 16464
rect 22388 15502 22416 18294
rect 22468 17740 22520 17746
rect 22468 17682 22520 17688
rect 22480 16590 22508 17682
rect 22572 17218 22600 19382
rect 22756 18766 22784 19926
rect 23032 19514 23060 20470
rect 23020 19508 23072 19514
rect 23020 19450 23072 19456
rect 22928 19440 22980 19446
rect 22928 19382 22980 19388
rect 22744 18760 22796 18766
rect 22744 18702 22796 18708
rect 22572 17190 22692 17218
rect 22560 17060 22612 17066
rect 22560 17002 22612 17008
rect 22572 16590 22600 17002
rect 22468 16584 22520 16590
rect 22468 16526 22520 16532
rect 22560 16584 22612 16590
rect 22560 16526 22612 16532
rect 22466 16144 22522 16153
rect 22466 16079 22522 16088
rect 22376 15496 22428 15502
rect 22376 15438 22428 15444
rect 22480 15042 22508 16079
rect 22296 15014 22508 15042
rect 22296 11778 22324 15014
rect 22664 14464 22692 17190
rect 22756 14822 22784 18702
rect 22836 17264 22888 17270
rect 22836 17206 22888 17212
rect 22848 15162 22876 17206
rect 22940 16046 22968 19382
rect 23124 16658 23152 24346
rect 23216 17270 23244 31894
rect 24596 30802 24624 37062
rect 24676 33516 24728 33522
rect 24676 33458 24728 33464
rect 24584 30796 24636 30802
rect 24584 30738 24636 30744
rect 23572 30048 23624 30054
rect 23572 29990 23624 29996
rect 23296 26784 23348 26790
rect 23296 26726 23348 26732
rect 23308 25906 23336 26726
rect 23296 25900 23348 25906
rect 23296 25842 23348 25848
rect 23296 24336 23348 24342
rect 23296 24278 23348 24284
rect 23308 23186 23336 24278
rect 23480 24064 23532 24070
rect 23480 24006 23532 24012
rect 23388 23792 23440 23798
rect 23388 23734 23440 23740
rect 23400 23322 23428 23734
rect 23492 23662 23520 24006
rect 23480 23656 23532 23662
rect 23480 23598 23532 23604
rect 23388 23316 23440 23322
rect 23388 23258 23440 23264
rect 23492 23202 23520 23598
rect 23296 23180 23348 23186
rect 23296 23122 23348 23128
rect 23400 23174 23520 23202
rect 23296 21480 23348 21486
rect 23296 21422 23348 21428
rect 23308 20398 23336 21422
rect 23296 20392 23348 20398
rect 23296 20334 23348 20340
rect 23400 20058 23428 23174
rect 23584 22094 23612 29990
rect 24216 25968 24268 25974
rect 24216 25910 24268 25916
rect 23492 22066 23612 22094
rect 24228 22094 24256 25910
rect 24400 25696 24452 25702
rect 24400 25638 24452 25644
rect 24308 24812 24360 24818
rect 24308 24754 24360 24760
rect 24320 24070 24348 24754
rect 24308 24064 24360 24070
rect 24308 24006 24360 24012
rect 24228 22066 24348 22094
rect 23492 21894 23520 22066
rect 23480 21888 23532 21894
rect 23480 21830 23532 21836
rect 23572 21888 23624 21894
rect 23572 21830 23624 21836
rect 23584 21622 23612 21830
rect 23572 21616 23624 21622
rect 23572 21558 23624 21564
rect 23572 21072 23624 21078
rect 23756 21072 23808 21078
rect 23572 21014 23624 21020
rect 23754 21040 23756 21049
rect 23808 21040 23810 21049
rect 23388 20052 23440 20058
rect 23388 19994 23440 20000
rect 23584 18358 23612 21014
rect 23754 20975 23810 20984
rect 23848 18964 23900 18970
rect 23848 18906 23900 18912
rect 23572 18352 23624 18358
rect 23572 18294 23624 18300
rect 23664 18284 23716 18290
rect 23664 18226 23716 18232
rect 23388 18216 23440 18222
rect 23388 18158 23440 18164
rect 23296 17740 23348 17746
rect 23296 17682 23348 17688
rect 23308 17338 23336 17682
rect 23400 17338 23428 18158
rect 23296 17332 23348 17338
rect 23296 17274 23348 17280
rect 23388 17332 23440 17338
rect 23388 17274 23440 17280
rect 23204 17264 23256 17270
rect 23204 17206 23256 17212
rect 23112 16652 23164 16658
rect 23112 16594 23164 16600
rect 23124 16046 23152 16594
rect 23388 16584 23440 16590
rect 23386 16552 23388 16561
rect 23440 16552 23442 16561
rect 23386 16487 23442 16496
rect 23676 16114 23704 18226
rect 23860 17610 23888 18906
rect 23848 17604 23900 17610
rect 23848 17546 23900 17552
rect 23860 16266 23888 17546
rect 24216 17264 24268 17270
rect 24216 17206 24268 17212
rect 24228 16794 24256 17206
rect 24216 16788 24268 16794
rect 24216 16730 24268 16736
rect 23768 16238 23888 16266
rect 23664 16108 23716 16114
rect 23664 16050 23716 16056
rect 22928 16040 22980 16046
rect 23112 16040 23164 16046
rect 22980 15988 23060 15994
rect 22928 15982 23060 15988
rect 23112 15982 23164 15988
rect 22940 15966 23060 15982
rect 22836 15156 22888 15162
rect 22836 15098 22888 15104
rect 22744 14816 22796 14822
rect 22744 14758 22796 14764
rect 22572 14436 22692 14464
rect 22572 13410 22600 14436
rect 22652 14340 22704 14346
rect 22652 14282 22704 14288
rect 22480 13382 22600 13410
rect 22480 13002 22508 13382
rect 22388 12974 22508 13002
rect 22664 12986 22692 14282
rect 22928 13796 22980 13802
rect 22928 13738 22980 13744
rect 22836 13456 22888 13462
rect 22836 13398 22888 13404
rect 22652 12980 22704 12986
rect 22388 12714 22416 12974
rect 22652 12922 22704 12928
rect 22664 12889 22692 12922
rect 22650 12880 22706 12889
rect 22468 12844 22520 12850
rect 22650 12815 22706 12824
rect 22468 12786 22520 12792
rect 22376 12708 22428 12714
rect 22376 12650 22428 12656
rect 22376 12164 22428 12170
rect 22376 12106 22428 12112
rect 22388 11898 22416 12106
rect 22376 11892 22428 11898
rect 22376 11834 22428 11840
rect 22296 11750 22416 11778
rect 22284 11620 22336 11626
rect 22284 11562 22336 11568
rect 22296 11286 22324 11562
rect 22284 11280 22336 11286
rect 22284 11222 22336 11228
rect 22388 7993 22416 11750
rect 22374 7984 22430 7993
rect 22374 7919 22430 7928
rect 22376 7880 22428 7886
rect 22376 7822 22428 7828
rect 22388 6798 22416 7822
rect 22376 6792 22428 6798
rect 22376 6734 22428 6740
rect 22008 6656 22060 6662
rect 22006 6624 22008 6633
rect 22192 6656 22244 6662
rect 22060 6624 22062 6633
rect 22192 6598 22244 6604
rect 22006 6559 22062 6568
rect 22008 6384 22060 6390
rect 22008 6326 22060 6332
rect 21916 6112 21968 6118
rect 21916 6054 21968 6060
rect 22020 5817 22048 6326
rect 22100 6316 22152 6322
rect 22100 6258 22152 6264
rect 22006 5808 22062 5817
rect 21916 5772 21968 5778
rect 22006 5743 22062 5752
rect 21916 5714 21968 5720
rect 21928 5545 21956 5714
rect 21914 5536 21970 5545
rect 21914 5471 21970 5480
rect 21916 5364 21968 5370
rect 21916 5306 21968 5312
rect 21928 5250 21956 5306
rect 21928 5222 22048 5250
rect 22020 5098 22048 5222
rect 21916 5092 21968 5098
rect 21916 5034 21968 5040
rect 22008 5092 22060 5098
rect 22008 5034 22060 5040
rect 21928 5001 21956 5034
rect 21914 4992 21970 5001
rect 21914 4927 21970 4936
rect 21914 4856 21970 4865
rect 21970 4826 22048 4842
rect 21970 4820 22060 4826
rect 21970 4814 22008 4820
rect 21914 4791 21970 4800
rect 22008 4762 22060 4768
rect 21916 4480 21968 4486
rect 21916 4422 21968 4428
rect 21928 4146 21956 4422
rect 21916 4140 21968 4146
rect 21916 4082 21968 4088
rect 21822 4040 21878 4049
rect 21822 3975 21878 3984
rect 21732 3052 21784 3058
rect 21732 2994 21784 3000
rect 20536 2984 20588 2990
rect 20720 2984 20772 2990
rect 20536 2926 20588 2932
rect 20640 2944 20720 2972
rect 20076 2790 20128 2796
rect 20258 2816 20314 2825
rect 20258 2751 20314 2760
rect 20444 2644 20496 2650
rect 20640 2632 20668 2944
rect 20720 2926 20772 2932
rect 21836 2854 21864 3975
rect 21916 3528 21968 3534
rect 21916 3470 21968 3476
rect 21824 2848 21876 2854
rect 21824 2790 21876 2796
rect 20496 2604 20668 2632
rect 20444 2586 20496 2592
rect 19614 2544 19670 2553
rect 19614 2479 19670 2488
rect 21272 2440 21324 2446
rect 19522 2408 19578 2417
rect 19432 2372 19484 2378
rect 19522 2343 19578 2352
rect 19706 2408 19762 2417
rect 21928 2417 21956 3470
rect 22112 2774 22140 6258
rect 22284 6180 22336 6186
rect 22284 6122 22336 6128
rect 22296 5914 22324 6122
rect 22480 6066 22508 12786
rect 22848 12714 22876 13398
rect 22940 13326 22968 13738
rect 22928 13320 22980 13326
rect 22928 13262 22980 13268
rect 22836 12708 22888 12714
rect 22836 12650 22888 12656
rect 22848 12434 22876 12650
rect 22664 12406 22876 12434
rect 22560 10668 22612 10674
rect 22560 10610 22612 10616
rect 22572 9722 22600 10610
rect 22560 9716 22612 9722
rect 22560 9658 22612 9664
rect 22480 6038 22600 6066
rect 22284 5908 22336 5914
rect 22468 5908 22520 5914
rect 22284 5850 22336 5856
rect 22388 5868 22468 5896
rect 22192 5704 22244 5710
rect 22192 5646 22244 5652
rect 22204 3738 22232 5646
rect 22388 5030 22416 5868
rect 22468 5850 22520 5856
rect 22468 5568 22520 5574
rect 22466 5536 22468 5545
rect 22520 5536 22522 5545
rect 22466 5471 22522 5480
rect 22572 5386 22600 6038
rect 22480 5358 22600 5386
rect 22376 5024 22428 5030
rect 22376 4966 22428 4972
rect 22284 4480 22336 4486
rect 22284 4422 22336 4428
rect 22192 3732 22244 3738
rect 22192 3674 22244 3680
rect 22296 3534 22324 4422
rect 22480 3777 22508 5358
rect 22560 5296 22612 5302
rect 22560 5238 22612 5244
rect 22572 4146 22600 5238
rect 22560 4140 22612 4146
rect 22560 4082 22612 4088
rect 22664 3942 22692 12406
rect 22836 10464 22888 10470
rect 22836 10406 22888 10412
rect 22744 9988 22796 9994
rect 22744 9930 22796 9936
rect 22756 9178 22784 9930
rect 22744 9172 22796 9178
rect 22744 9114 22796 9120
rect 22848 8378 22876 10406
rect 22756 8350 22876 8378
rect 22756 6066 22784 8350
rect 22940 8242 22968 13262
rect 23032 12209 23060 15966
rect 23204 15972 23256 15978
rect 23204 15914 23256 15920
rect 23112 15700 23164 15706
rect 23112 15642 23164 15648
rect 23124 14958 23152 15642
rect 23216 15162 23244 15914
rect 23664 15428 23716 15434
rect 23664 15370 23716 15376
rect 23296 15360 23348 15366
rect 23296 15302 23348 15308
rect 23204 15156 23256 15162
rect 23204 15098 23256 15104
rect 23112 14952 23164 14958
rect 23112 14894 23164 14900
rect 23124 14822 23152 14894
rect 23112 14816 23164 14822
rect 23112 14758 23164 14764
rect 23202 14648 23258 14657
rect 23202 14583 23258 14592
rect 23216 14550 23244 14583
rect 23204 14544 23256 14550
rect 23204 14486 23256 14492
rect 23308 13852 23336 15302
rect 23572 14408 23624 14414
rect 23572 14350 23624 14356
rect 23388 13864 23440 13870
rect 23308 13824 23388 13852
rect 23308 13394 23336 13824
rect 23388 13806 23440 13812
rect 23296 13388 23348 13394
rect 23296 13330 23348 13336
rect 23110 12880 23166 12889
rect 23110 12815 23166 12824
rect 23018 12200 23074 12209
rect 23018 12135 23074 12144
rect 23020 11144 23072 11150
rect 23020 11086 23072 11092
rect 23032 8974 23060 11086
rect 23020 8968 23072 8974
rect 23020 8910 23072 8916
rect 22848 8214 22968 8242
rect 22848 6254 22876 8214
rect 22928 7812 22980 7818
rect 22928 7754 22980 7760
rect 22836 6248 22888 6254
rect 22836 6190 22888 6196
rect 22756 6038 22876 6066
rect 22742 5808 22798 5817
rect 22742 5743 22798 5752
rect 22756 4282 22784 5743
rect 22744 4276 22796 4282
rect 22744 4218 22796 4224
rect 22652 3936 22704 3942
rect 22652 3878 22704 3884
rect 22466 3768 22522 3777
rect 22466 3703 22522 3712
rect 22664 3602 22692 3878
rect 22652 3596 22704 3602
rect 22652 3538 22704 3544
rect 22744 3596 22796 3602
rect 22744 3538 22796 3544
rect 22284 3528 22336 3534
rect 22284 3470 22336 3476
rect 22756 3466 22784 3538
rect 22744 3460 22796 3466
rect 22744 3402 22796 3408
rect 22112 2746 22416 2774
rect 22388 2582 22416 2746
rect 22376 2576 22428 2582
rect 22376 2518 22428 2524
rect 22742 2544 22798 2553
rect 22742 2479 22798 2488
rect 21272 2382 21324 2388
rect 21914 2408 21970 2417
rect 19706 2343 19708 2352
rect 19432 2314 19484 2320
rect 19760 2343 19762 2352
rect 19708 2314 19760 2320
rect 19444 1562 19472 2314
rect 21180 2304 21232 2310
rect 21180 2246 21232 2252
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 21192 1834 21220 2246
rect 21180 1828 21232 1834
rect 21180 1770 21232 1776
rect 19984 1692 20036 1698
rect 19984 1634 20036 1640
rect 19432 1556 19484 1562
rect 19432 1498 19484 1504
rect 19996 800 20024 1634
rect 21284 800 21312 2382
rect 21914 2343 21970 2352
rect 22560 2304 22612 2310
rect 22560 2246 22612 2252
rect 22572 800 22600 2246
rect 22756 2106 22784 2479
rect 22744 2100 22796 2106
rect 22744 2042 22796 2048
rect 22848 1902 22876 6038
rect 22940 5166 22968 7754
rect 23124 7478 23152 12815
rect 23478 12472 23534 12481
rect 23204 12436 23256 12442
rect 23478 12407 23534 12416
rect 23204 12378 23256 12384
rect 23216 11354 23244 12378
rect 23388 12300 23440 12306
rect 23388 12242 23440 12248
rect 23294 12200 23350 12209
rect 23294 12135 23296 12144
rect 23348 12135 23350 12144
rect 23296 12106 23348 12112
rect 23400 12073 23428 12242
rect 23386 12064 23442 12073
rect 23386 11999 23442 12008
rect 23296 11824 23348 11830
rect 23296 11766 23348 11772
rect 23388 11824 23440 11830
rect 23388 11766 23440 11772
rect 23204 11348 23256 11354
rect 23204 11290 23256 11296
rect 23308 10266 23336 11766
rect 23296 10260 23348 10266
rect 23296 10202 23348 10208
rect 23400 10146 23428 11766
rect 23492 10606 23520 12407
rect 23584 12102 23612 14350
rect 23572 12096 23624 12102
rect 23572 12038 23624 12044
rect 23676 11694 23704 15370
rect 23664 11688 23716 11694
rect 23664 11630 23716 11636
rect 23572 11280 23624 11286
rect 23572 11222 23624 11228
rect 23480 10600 23532 10606
rect 23480 10542 23532 10548
rect 23308 10118 23428 10146
rect 23112 7472 23164 7478
rect 23112 7414 23164 7420
rect 23020 6792 23072 6798
rect 23020 6734 23072 6740
rect 23032 6390 23060 6734
rect 23112 6656 23164 6662
rect 23112 6598 23164 6604
rect 23020 6384 23072 6390
rect 23020 6326 23072 6332
rect 23020 6112 23072 6118
rect 23020 6054 23072 6060
rect 23032 5778 23060 6054
rect 23020 5772 23072 5778
rect 23020 5714 23072 5720
rect 23124 5642 23152 6598
rect 23308 6497 23336 10118
rect 23480 8968 23532 8974
rect 23480 8910 23532 8916
rect 23388 8424 23440 8430
rect 23388 8366 23440 8372
rect 23400 7546 23428 8366
rect 23388 7540 23440 7546
rect 23388 7482 23440 7488
rect 23492 6633 23520 8910
rect 23584 8634 23612 11222
rect 23768 10826 23796 16238
rect 24216 15904 24268 15910
rect 24216 15846 24268 15852
rect 24228 15638 24256 15846
rect 24216 15632 24268 15638
rect 24216 15574 24268 15580
rect 24320 14414 24348 22066
rect 24412 20466 24440 25638
rect 24688 25498 24716 33458
rect 25516 27606 25544 37130
rect 26436 37126 26464 39200
rect 27724 37262 27752 39200
rect 29012 37262 29040 39200
rect 29656 37330 29684 39200
rect 29644 37324 29696 37330
rect 29644 37266 29696 37272
rect 27160 37256 27212 37262
rect 27160 37198 27212 37204
rect 27712 37256 27764 37262
rect 27712 37198 27764 37204
rect 29000 37256 29052 37262
rect 29000 37198 29052 37204
rect 25872 37120 25924 37126
rect 25872 37062 25924 37068
rect 26424 37120 26476 37126
rect 26424 37062 26476 37068
rect 25688 32292 25740 32298
rect 25688 32234 25740 32240
rect 25700 31822 25728 32234
rect 25688 31816 25740 31822
rect 25688 31758 25740 31764
rect 25884 30734 25912 37062
rect 27172 36922 27200 37198
rect 30944 37126 30972 39200
rect 32232 37262 32260 39200
rect 31024 37256 31076 37262
rect 31024 37198 31076 37204
rect 32220 37256 32272 37262
rect 32220 37198 32272 37204
rect 27436 37120 27488 37126
rect 27436 37062 27488 37068
rect 29736 37120 29788 37126
rect 29736 37062 29788 37068
rect 30380 37120 30432 37126
rect 30380 37062 30432 37068
rect 30932 37120 30984 37126
rect 30932 37062 30984 37068
rect 27160 36916 27212 36922
rect 27160 36858 27212 36864
rect 27252 31884 27304 31890
rect 27252 31826 27304 31832
rect 26884 31816 26936 31822
rect 26884 31758 26936 31764
rect 25872 30728 25924 30734
rect 25872 30670 25924 30676
rect 25504 27600 25556 27606
rect 25504 27542 25556 27548
rect 24768 25696 24820 25702
rect 24768 25638 24820 25644
rect 24676 25492 24728 25498
rect 24676 25434 24728 25440
rect 24780 25242 24808 25638
rect 24688 25214 24808 25242
rect 24584 24268 24636 24274
rect 24584 24210 24636 24216
rect 24596 23730 24624 24210
rect 24584 23724 24636 23730
rect 24584 23666 24636 23672
rect 24688 23594 24716 25214
rect 24768 25152 24820 25158
rect 24768 25094 24820 25100
rect 24780 24274 24808 25094
rect 26896 24818 26924 31758
rect 27160 29640 27212 29646
rect 27160 29582 27212 29588
rect 25780 24812 25832 24818
rect 25780 24754 25832 24760
rect 26884 24812 26936 24818
rect 26884 24754 26936 24760
rect 25792 24410 25820 24754
rect 27172 24682 27200 29582
rect 27160 24676 27212 24682
rect 27160 24618 27212 24624
rect 25780 24404 25832 24410
rect 25780 24346 25832 24352
rect 24860 24336 24912 24342
rect 24860 24278 24912 24284
rect 24768 24268 24820 24274
rect 24768 24210 24820 24216
rect 24768 24064 24820 24070
rect 24768 24006 24820 24012
rect 24676 23588 24728 23594
rect 24676 23530 24728 23536
rect 24688 23254 24716 23530
rect 24676 23248 24728 23254
rect 24676 23190 24728 23196
rect 24780 22574 24808 24006
rect 24872 22710 24900 24278
rect 27160 23588 27212 23594
rect 27160 23530 27212 23536
rect 25136 23520 25188 23526
rect 25136 23462 25188 23468
rect 25044 23044 25096 23050
rect 25044 22986 25096 22992
rect 25056 22778 25084 22986
rect 25044 22772 25096 22778
rect 25044 22714 25096 22720
rect 24860 22704 24912 22710
rect 24860 22646 24912 22652
rect 24768 22568 24820 22574
rect 24768 22510 24820 22516
rect 24780 22094 24808 22510
rect 24872 22250 24900 22646
rect 25044 22636 25096 22642
rect 25044 22578 25096 22584
rect 24872 22222 24992 22250
rect 24596 22066 24808 22094
rect 24400 20460 24452 20466
rect 24400 20402 24452 20408
rect 24492 19848 24544 19854
rect 24492 19790 24544 19796
rect 24504 19378 24532 19790
rect 24492 19372 24544 19378
rect 24492 19314 24544 19320
rect 24596 19242 24624 22066
rect 24768 21344 24820 21350
rect 24768 21286 24820 21292
rect 24676 19848 24728 19854
rect 24676 19790 24728 19796
rect 24688 19514 24716 19790
rect 24676 19508 24728 19514
rect 24676 19450 24728 19456
rect 24584 19236 24636 19242
rect 24584 19178 24636 19184
rect 24676 18692 24728 18698
rect 24676 18634 24728 18640
rect 24688 18222 24716 18634
rect 24780 18290 24808 21286
rect 24964 19922 24992 22222
rect 25056 22166 25084 22578
rect 25044 22160 25096 22166
rect 25044 22102 25096 22108
rect 25044 20800 25096 20806
rect 25044 20742 25096 20748
rect 25056 20466 25084 20742
rect 25148 20602 25176 23462
rect 26884 22568 26936 22574
rect 26884 22510 26936 22516
rect 25412 22160 25464 22166
rect 25412 22102 25464 22108
rect 25228 20936 25280 20942
rect 25228 20878 25280 20884
rect 25136 20596 25188 20602
rect 25136 20538 25188 20544
rect 25044 20460 25096 20466
rect 25044 20402 25096 20408
rect 25136 20256 25188 20262
rect 25136 20198 25188 20204
rect 25148 19990 25176 20198
rect 25240 20058 25268 20878
rect 25228 20052 25280 20058
rect 25228 19994 25280 20000
rect 25136 19984 25188 19990
rect 25136 19926 25188 19932
rect 25424 19922 25452 22102
rect 25780 21004 25832 21010
rect 25780 20946 25832 20952
rect 25792 20466 25820 20946
rect 25780 20460 25832 20466
rect 25780 20402 25832 20408
rect 24952 19916 25004 19922
rect 24952 19858 25004 19864
rect 25412 19916 25464 19922
rect 25412 19858 25464 19864
rect 25504 19780 25556 19786
rect 25504 19722 25556 19728
rect 25320 19712 25372 19718
rect 25320 19654 25372 19660
rect 25332 18698 25360 19654
rect 25516 19378 25544 19722
rect 25792 19514 25820 20402
rect 26792 20324 26844 20330
rect 26792 20266 26844 20272
rect 26700 19848 26752 19854
rect 26700 19790 26752 19796
rect 26516 19712 26568 19718
rect 26516 19654 26568 19660
rect 25780 19508 25832 19514
rect 25780 19450 25832 19456
rect 25504 19372 25556 19378
rect 25504 19314 25556 19320
rect 26056 19304 26108 19310
rect 26056 19246 26108 19252
rect 26068 18970 26096 19246
rect 26056 18964 26108 18970
rect 26056 18906 26108 18912
rect 25688 18896 25740 18902
rect 25688 18838 25740 18844
rect 25320 18692 25372 18698
rect 25320 18634 25372 18640
rect 24768 18284 24820 18290
rect 24768 18226 24820 18232
rect 25700 18222 25728 18838
rect 26528 18698 26556 19654
rect 26608 19372 26660 19378
rect 26608 19314 26660 19320
rect 26620 18834 26648 19314
rect 26608 18828 26660 18834
rect 26608 18770 26660 18776
rect 26516 18692 26568 18698
rect 26516 18634 26568 18640
rect 25964 18624 26016 18630
rect 25964 18566 26016 18572
rect 24676 18216 24728 18222
rect 24676 18158 24728 18164
rect 25688 18216 25740 18222
rect 25688 18158 25740 18164
rect 25976 17610 26004 18566
rect 25964 17604 26016 17610
rect 25964 17546 26016 17552
rect 24768 17536 24820 17542
rect 24768 17478 24820 17484
rect 24400 17128 24452 17134
rect 24400 17070 24452 17076
rect 24412 16726 24440 17070
rect 24780 16998 24808 17478
rect 24952 17060 25004 17066
rect 24952 17002 25004 17008
rect 24584 16992 24636 16998
rect 24584 16934 24636 16940
rect 24768 16992 24820 16998
rect 24768 16934 24820 16940
rect 24400 16720 24452 16726
rect 24400 16662 24452 16668
rect 24492 16448 24544 16454
rect 24492 16390 24544 16396
rect 24400 15700 24452 15706
rect 24400 15642 24452 15648
rect 24412 15434 24440 15642
rect 24400 15428 24452 15434
rect 24400 15370 24452 15376
rect 24308 14408 24360 14414
rect 24308 14350 24360 14356
rect 24308 14272 24360 14278
rect 24308 14214 24360 14220
rect 24032 14000 24084 14006
rect 24032 13942 24084 13948
rect 23940 13184 23992 13190
rect 23940 13126 23992 13132
rect 23848 12912 23900 12918
rect 23848 12854 23900 12860
rect 23860 11354 23888 12854
rect 23952 12782 23980 13126
rect 23940 12776 23992 12782
rect 23940 12718 23992 12724
rect 23848 11348 23900 11354
rect 23848 11290 23900 11296
rect 23768 10798 23980 10826
rect 23756 10736 23808 10742
rect 23756 10678 23808 10684
rect 23664 9648 23716 9654
rect 23664 9590 23716 9596
rect 23676 9178 23704 9590
rect 23664 9172 23716 9178
rect 23664 9114 23716 9120
rect 23572 8628 23624 8634
rect 23572 8570 23624 8576
rect 23664 8492 23716 8498
rect 23664 8434 23716 8440
rect 23676 7886 23704 8434
rect 23768 8090 23796 10678
rect 23848 10600 23900 10606
rect 23848 10542 23900 10548
rect 23756 8084 23808 8090
rect 23756 8026 23808 8032
rect 23754 7984 23810 7993
rect 23754 7919 23810 7928
rect 23664 7880 23716 7886
rect 23664 7822 23716 7828
rect 23478 6624 23534 6633
rect 23478 6559 23534 6568
rect 23294 6488 23350 6497
rect 23294 6423 23350 6432
rect 23388 6452 23440 6458
rect 23388 6394 23440 6400
rect 23204 6112 23256 6118
rect 23204 6054 23256 6060
rect 23020 5636 23072 5642
rect 23020 5578 23072 5584
rect 23112 5636 23164 5642
rect 23112 5578 23164 5584
rect 23032 5522 23060 5578
rect 23216 5522 23244 6054
rect 23032 5494 23244 5522
rect 22928 5160 22980 5166
rect 22928 5102 22980 5108
rect 23204 5160 23256 5166
rect 23204 5102 23256 5108
rect 23216 4078 23244 5102
rect 23400 5030 23428 6394
rect 23768 6254 23796 7919
rect 23664 6248 23716 6254
rect 23664 6190 23716 6196
rect 23756 6248 23808 6254
rect 23756 6190 23808 6196
rect 23676 5778 23704 6190
rect 23860 6186 23888 10542
rect 23952 9518 23980 10798
rect 24044 10198 24072 13942
rect 24320 12918 24348 14214
rect 24412 13462 24440 13493
rect 24400 13456 24452 13462
rect 24398 13424 24400 13433
rect 24452 13424 24454 13433
rect 24398 13359 24454 13368
rect 24308 12912 24360 12918
rect 24308 12854 24360 12860
rect 24412 12434 24440 13359
rect 24504 13258 24532 16390
rect 24596 14006 24624 16934
rect 24676 15360 24728 15366
rect 24676 15302 24728 15308
rect 24768 15360 24820 15366
rect 24768 15302 24820 15308
rect 24688 15094 24716 15302
rect 24676 15088 24728 15094
rect 24676 15030 24728 15036
rect 24780 14958 24808 15302
rect 24768 14952 24820 14958
rect 24768 14894 24820 14900
rect 24676 14272 24728 14278
rect 24676 14214 24728 14220
rect 24768 14272 24820 14278
rect 24768 14214 24820 14220
rect 24584 14000 24636 14006
rect 24584 13942 24636 13948
rect 24688 13394 24716 14214
rect 24780 14006 24808 14214
rect 24768 14000 24820 14006
rect 24768 13942 24820 13948
rect 24676 13388 24728 13394
rect 24676 13330 24728 13336
rect 24492 13252 24544 13258
rect 24492 13194 24544 13200
rect 24688 12782 24716 13330
rect 24676 12776 24728 12782
rect 24676 12718 24728 12724
rect 24320 12406 24440 12434
rect 24584 12436 24636 12442
rect 24216 11688 24268 11694
rect 24214 11656 24216 11665
rect 24268 11656 24270 11665
rect 24214 11591 24270 11600
rect 24216 11144 24268 11150
rect 24216 11086 24268 11092
rect 24032 10192 24084 10198
rect 24032 10134 24084 10140
rect 23940 9512 23992 9518
rect 24032 9512 24084 9518
rect 23940 9454 23992 9460
rect 24030 9480 24032 9489
rect 24084 9480 24086 9489
rect 23848 6180 23900 6186
rect 23848 6122 23900 6128
rect 23664 5772 23716 5778
rect 23664 5714 23716 5720
rect 23296 5024 23348 5030
rect 23296 4966 23348 4972
rect 23388 5024 23440 5030
rect 23388 4966 23440 4972
rect 23308 4214 23336 4966
rect 23846 4448 23902 4457
rect 23846 4383 23902 4392
rect 23296 4208 23348 4214
rect 23296 4150 23348 4156
rect 23204 4072 23256 4078
rect 23204 4014 23256 4020
rect 23216 3194 23244 4014
rect 23756 4004 23808 4010
rect 23756 3946 23808 3952
rect 23386 3768 23442 3777
rect 23386 3703 23442 3712
rect 23296 3528 23348 3534
rect 23296 3470 23348 3476
rect 23308 3369 23336 3470
rect 23294 3360 23350 3369
rect 23294 3295 23350 3304
rect 23204 3188 23256 3194
rect 23204 3130 23256 3136
rect 23400 3058 23428 3703
rect 23768 3534 23796 3946
rect 23860 3738 23888 4383
rect 23848 3732 23900 3738
rect 23848 3674 23900 3680
rect 23756 3528 23808 3534
rect 23756 3470 23808 3476
rect 23388 3052 23440 3058
rect 23388 2994 23440 3000
rect 22928 2644 22980 2650
rect 22928 2586 22980 2592
rect 22940 2106 22968 2586
rect 23952 2514 23980 9454
rect 24030 9415 24086 9424
rect 24032 8628 24084 8634
rect 24032 8570 24084 8576
rect 24044 6390 24072 8570
rect 24124 8560 24176 8566
rect 24124 8502 24176 8508
rect 24032 6384 24084 6390
rect 24032 6326 24084 6332
rect 24030 5536 24086 5545
rect 24030 5471 24086 5480
rect 24044 5166 24072 5471
rect 24032 5160 24084 5166
rect 24032 5102 24084 5108
rect 24136 4690 24164 8502
rect 24228 8498 24256 11086
rect 24216 8492 24268 8498
rect 24216 8434 24268 8440
rect 24228 7954 24256 8434
rect 24216 7948 24268 7954
rect 24216 7890 24268 7896
rect 24216 7336 24268 7342
rect 24216 7278 24268 7284
rect 24228 7177 24256 7278
rect 24214 7168 24270 7177
rect 24214 7103 24270 7112
rect 24320 5642 24348 12406
rect 24780 12434 24808 13942
rect 24584 12378 24636 12384
rect 24688 12406 24808 12434
rect 24492 12096 24544 12102
rect 24490 12064 24492 12073
rect 24544 12064 24546 12073
rect 24490 11999 24546 12008
rect 24492 7880 24544 7886
rect 24492 7822 24544 7828
rect 24504 7274 24532 7822
rect 24492 7268 24544 7274
rect 24492 7210 24544 7216
rect 24308 5636 24360 5642
rect 24308 5578 24360 5584
rect 24400 5568 24452 5574
rect 24400 5510 24452 5516
rect 24124 4684 24176 4690
rect 24124 4626 24176 4632
rect 24136 4162 24164 4626
rect 24044 4134 24164 4162
rect 24044 3194 24072 4134
rect 24412 4078 24440 5510
rect 24596 5234 24624 12378
rect 24688 11626 24716 12406
rect 24768 12232 24820 12238
rect 24768 12174 24820 12180
rect 24780 11898 24808 12174
rect 24768 11892 24820 11898
rect 24768 11834 24820 11840
rect 24676 11620 24728 11626
rect 24676 11562 24728 11568
rect 24964 10690 24992 17002
rect 26332 16584 26384 16590
rect 26332 16526 26384 16532
rect 26148 15632 26200 15638
rect 26148 15574 26200 15580
rect 26056 15496 26108 15502
rect 26056 15438 26108 15444
rect 26068 15162 26096 15438
rect 26056 15156 26108 15162
rect 26056 15098 26108 15104
rect 25228 14884 25280 14890
rect 25228 14826 25280 14832
rect 25136 12164 25188 12170
rect 25136 12106 25188 12112
rect 25148 11286 25176 12106
rect 25136 11280 25188 11286
rect 25136 11222 25188 11228
rect 25148 11082 25176 11222
rect 25136 11076 25188 11082
rect 25136 11018 25188 11024
rect 24964 10662 25176 10690
rect 24952 10532 25004 10538
rect 24952 10474 25004 10480
rect 24674 10160 24730 10169
rect 24674 10095 24676 10104
rect 24728 10095 24730 10104
rect 24676 10066 24728 10072
rect 24768 9988 24820 9994
rect 24768 9930 24820 9936
rect 24780 8090 24808 9930
rect 24964 8906 24992 10474
rect 24952 8900 25004 8906
rect 24952 8842 25004 8848
rect 25044 8900 25096 8906
rect 25044 8842 25096 8848
rect 25056 8634 25084 8842
rect 25044 8628 25096 8634
rect 25044 8570 25096 8576
rect 24768 8084 24820 8090
rect 24768 8026 24820 8032
rect 24768 7948 24820 7954
rect 24768 7890 24820 7896
rect 24780 7410 24808 7890
rect 24952 7880 25004 7886
rect 24952 7822 25004 7828
rect 24768 7404 24820 7410
rect 24768 7346 24820 7352
rect 24964 7342 24992 7822
rect 24952 7336 25004 7342
rect 24952 7278 25004 7284
rect 24858 7168 24914 7177
rect 25148 7154 25176 10662
rect 24858 7103 24914 7112
rect 24964 7126 25176 7154
rect 24584 5228 24636 5234
rect 24584 5170 24636 5176
rect 24596 5001 24624 5170
rect 24582 4992 24638 5001
rect 24582 4927 24638 4936
rect 24766 4584 24822 4593
rect 24766 4519 24768 4528
rect 24820 4519 24822 4528
rect 24768 4490 24820 4496
rect 24768 4276 24820 4282
rect 24768 4218 24820 4224
rect 24124 4072 24176 4078
rect 24122 4040 24124 4049
rect 24400 4072 24452 4078
rect 24176 4040 24178 4049
rect 24780 4049 24808 4218
rect 24872 4078 24900 7103
rect 24964 6730 24992 7126
rect 25240 6866 25268 14826
rect 25412 14476 25464 14482
rect 25412 14418 25464 14424
rect 25688 14476 25740 14482
rect 25688 14418 25740 14424
rect 25320 12096 25372 12102
rect 25320 12038 25372 12044
rect 25332 11082 25360 12038
rect 25424 11082 25452 14418
rect 25596 13932 25648 13938
rect 25596 13874 25648 13880
rect 25608 13297 25636 13874
rect 25594 13288 25650 13297
rect 25594 13223 25650 13232
rect 25700 12850 25728 14418
rect 25780 14340 25832 14346
rect 25780 14282 25832 14288
rect 25792 14074 25820 14282
rect 25780 14068 25832 14074
rect 25780 14010 25832 14016
rect 25872 13932 25924 13938
rect 25872 13874 25924 13880
rect 25688 12844 25740 12850
rect 25688 12786 25740 12792
rect 25884 12434 25912 13874
rect 25964 13796 26016 13802
rect 25964 13738 26016 13744
rect 25700 12406 25912 12434
rect 25504 11824 25556 11830
rect 25504 11766 25556 11772
rect 25320 11076 25372 11082
rect 25320 11018 25372 11024
rect 25412 11076 25464 11082
rect 25412 11018 25464 11024
rect 25516 10810 25544 11766
rect 25504 10804 25556 10810
rect 25504 10746 25556 10752
rect 25700 9110 25728 12406
rect 25872 11076 25924 11082
rect 25872 11018 25924 11024
rect 25780 9444 25832 9450
rect 25780 9386 25832 9392
rect 25688 9104 25740 9110
rect 25688 9046 25740 9052
rect 25596 8832 25648 8838
rect 25596 8774 25648 8780
rect 25688 8832 25740 8838
rect 25688 8774 25740 8780
rect 25228 6860 25280 6866
rect 25228 6802 25280 6808
rect 24952 6724 25004 6730
rect 24952 6666 25004 6672
rect 24964 6633 24992 6666
rect 24950 6624 25006 6633
rect 24950 6559 25006 6568
rect 25320 6384 25372 6390
rect 25320 6326 25372 6332
rect 24952 6248 25004 6254
rect 24952 6190 25004 6196
rect 24964 4690 24992 6190
rect 25332 6186 25360 6326
rect 25320 6180 25372 6186
rect 25320 6122 25372 6128
rect 25608 5710 25636 8774
rect 25700 7324 25728 8774
rect 25792 7546 25820 9386
rect 25780 7540 25832 7546
rect 25780 7482 25832 7488
rect 25780 7336 25832 7342
rect 25700 7296 25780 7324
rect 25700 6984 25728 7296
rect 25780 7278 25832 7284
rect 25700 6956 25820 6984
rect 25596 5704 25648 5710
rect 25596 5646 25648 5652
rect 25686 5672 25742 5681
rect 25042 4856 25098 4865
rect 25042 4791 25098 4800
rect 24952 4684 25004 4690
rect 24952 4626 25004 4632
rect 25056 4214 25084 4791
rect 25504 4548 25556 4554
rect 25504 4490 25556 4496
rect 25516 4457 25544 4490
rect 25502 4448 25558 4457
rect 25502 4383 25558 4392
rect 25044 4208 25096 4214
rect 25044 4150 25096 4156
rect 24860 4072 24912 4078
rect 24400 4014 24452 4020
rect 24766 4040 24822 4049
rect 24122 3975 24178 3984
rect 24860 4014 24912 4020
rect 25608 4010 25636 5646
rect 25686 5607 25688 5616
rect 25740 5607 25742 5616
rect 25688 5578 25740 5584
rect 25688 5160 25740 5166
rect 25688 5102 25740 5108
rect 25700 4758 25728 5102
rect 25688 4752 25740 4758
rect 25688 4694 25740 4700
rect 24766 3975 24822 3984
rect 25596 4004 25648 4010
rect 25596 3946 25648 3952
rect 25320 3936 25372 3942
rect 25320 3878 25372 3884
rect 24492 3732 24544 3738
rect 24492 3674 24544 3680
rect 24032 3188 24084 3194
rect 24032 3130 24084 3136
rect 23940 2508 23992 2514
rect 23940 2450 23992 2456
rect 23112 2372 23164 2378
rect 23112 2314 23164 2320
rect 23204 2372 23256 2378
rect 23204 2314 23256 2320
rect 22928 2100 22980 2106
rect 22928 2042 22980 2048
rect 23124 2038 23152 2314
rect 23020 2032 23072 2038
rect 23020 1974 23072 1980
rect 23112 2032 23164 2038
rect 23112 1974 23164 1980
rect 22836 1896 22888 1902
rect 22836 1838 22888 1844
rect 23032 1698 23060 1974
rect 23020 1692 23072 1698
rect 23020 1634 23072 1640
rect 23216 800 23244 2314
rect 24504 800 24532 3674
rect 25332 3534 25360 3878
rect 25320 3528 25372 3534
rect 24674 3496 24730 3505
rect 25320 3470 25372 3476
rect 24674 3431 24676 3440
rect 24728 3431 24730 3440
rect 24676 3402 24728 3408
rect 24860 3392 24912 3398
rect 24860 3334 24912 3340
rect 24872 2990 24900 3334
rect 24860 2984 24912 2990
rect 24860 2926 24912 2932
rect 25136 2984 25188 2990
rect 25136 2926 25188 2932
rect 24952 2916 25004 2922
rect 24952 2858 25004 2864
rect 24860 2440 24912 2446
rect 24860 2382 24912 2388
rect 24872 1766 24900 2382
rect 24964 1902 24992 2858
rect 25148 2514 25176 2926
rect 25136 2508 25188 2514
rect 25700 2496 25728 4694
rect 25792 4690 25820 6956
rect 25780 4684 25832 4690
rect 25780 4626 25832 4632
rect 25792 4282 25820 4626
rect 25780 4276 25832 4282
rect 25780 4218 25832 4224
rect 25884 3466 25912 11018
rect 25976 10742 26004 13738
rect 26160 12434 26188 15574
rect 26240 15360 26292 15366
rect 26240 15302 26292 15308
rect 26252 15026 26280 15302
rect 26240 15020 26292 15026
rect 26240 14962 26292 14968
rect 26344 14362 26372 16526
rect 26424 15564 26476 15570
rect 26424 15506 26476 15512
rect 26252 14334 26372 14362
rect 26252 12986 26280 14334
rect 26332 14272 26384 14278
rect 26332 14214 26384 14220
rect 26344 14074 26372 14214
rect 26332 14068 26384 14074
rect 26332 14010 26384 14016
rect 26436 12986 26464 15506
rect 26516 15496 26568 15502
rect 26516 15438 26568 15444
rect 26240 12980 26292 12986
rect 26240 12922 26292 12928
rect 26424 12980 26476 12986
rect 26424 12922 26476 12928
rect 26424 12776 26476 12782
rect 26424 12718 26476 12724
rect 26436 12442 26464 12718
rect 26424 12436 26476 12442
rect 26160 12406 26280 12434
rect 26252 11778 26280 12406
rect 26424 12378 26476 12384
rect 26332 12232 26384 12238
rect 26528 12220 26556 15438
rect 26384 12192 26556 12220
rect 26332 12174 26384 12180
rect 26344 11898 26372 12174
rect 26332 11892 26384 11898
rect 26332 11834 26384 11840
rect 26252 11750 26556 11778
rect 26240 11688 26292 11694
rect 26240 11630 26292 11636
rect 26252 11218 26280 11630
rect 26240 11212 26292 11218
rect 26240 11154 26292 11160
rect 25964 10736 26016 10742
rect 25964 10678 26016 10684
rect 25964 9988 26016 9994
rect 25964 9930 26016 9936
rect 25976 8906 26004 9930
rect 25964 8900 26016 8906
rect 25964 8842 26016 8848
rect 25964 8492 26016 8498
rect 25964 8434 26016 8440
rect 25976 8090 26004 8434
rect 25964 8084 26016 8090
rect 25964 8026 26016 8032
rect 25976 6934 26004 8026
rect 26240 7812 26292 7818
rect 26240 7754 26292 7760
rect 26252 7546 26280 7754
rect 26240 7540 26292 7546
rect 26240 7482 26292 7488
rect 26528 7410 26556 11750
rect 26620 8634 26648 18770
rect 26712 13530 26740 19790
rect 26700 13524 26752 13530
rect 26700 13466 26752 13472
rect 26700 12980 26752 12986
rect 26700 12922 26752 12928
rect 26712 8906 26740 12922
rect 26804 11830 26832 20266
rect 26896 18698 26924 22510
rect 27068 22432 27120 22438
rect 27068 22374 27120 22380
rect 27080 21962 27108 22374
rect 26976 21956 27028 21962
rect 26976 21898 27028 21904
rect 27068 21956 27120 21962
rect 27068 21898 27120 21904
rect 26988 20602 27016 21898
rect 26976 20596 27028 20602
rect 26976 20538 27028 20544
rect 26988 19514 27016 20538
rect 27172 20466 27200 23530
rect 27264 22710 27292 31826
rect 27448 30326 27476 37062
rect 27988 36916 28040 36922
rect 27988 36858 28040 36864
rect 27528 36712 27580 36718
rect 27528 36654 27580 36660
rect 27436 30320 27488 30326
rect 27436 30262 27488 30268
rect 27540 28558 27568 36654
rect 28000 32026 28028 36858
rect 29644 32428 29696 32434
rect 29644 32370 29696 32376
rect 27988 32020 28040 32026
rect 27988 31962 28040 31968
rect 28080 30592 28132 30598
rect 28080 30534 28132 30540
rect 28092 30394 28120 30534
rect 28080 30388 28132 30394
rect 28080 30330 28132 30336
rect 29656 30326 29684 32370
rect 29748 32298 29776 37062
rect 29736 32292 29788 32298
rect 29736 32234 29788 32240
rect 30392 31890 30420 37062
rect 31036 36922 31064 37198
rect 31300 37120 31352 37126
rect 32876 37108 32904 39200
rect 34164 39114 34192 39200
rect 34256 39114 34284 39222
rect 34164 39086 34284 39114
rect 33232 37256 33284 37262
rect 33232 37198 33284 37204
rect 33140 37120 33192 37126
rect 32876 37080 33140 37108
rect 31300 37062 31352 37068
rect 33140 37062 33192 37068
rect 31024 36916 31076 36922
rect 31024 36858 31076 36864
rect 31116 32904 31168 32910
rect 31116 32846 31168 32852
rect 31128 32026 31156 32846
rect 31116 32020 31168 32026
rect 31116 31962 31168 31968
rect 30380 31884 30432 31890
rect 30380 31826 30432 31832
rect 30380 31340 30432 31346
rect 30380 31282 30432 31288
rect 29644 30320 29696 30326
rect 29644 30262 29696 30268
rect 29552 30252 29604 30258
rect 29552 30194 29604 30200
rect 27528 28552 27580 28558
rect 27528 28494 27580 28500
rect 27804 28416 27856 28422
rect 27804 28358 27856 28364
rect 27436 25288 27488 25294
rect 27436 25230 27488 25236
rect 27252 22704 27304 22710
rect 27252 22646 27304 22652
rect 27344 22704 27396 22710
rect 27344 22646 27396 22652
rect 27356 22234 27384 22646
rect 27344 22228 27396 22234
rect 27344 22170 27396 22176
rect 27160 20460 27212 20466
rect 27160 20402 27212 20408
rect 26976 19508 27028 19514
rect 26976 19450 27028 19456
rect 27172 19378 27200 20402
rect 27160 19372 27212 19378
rect 27160 19314 27212 19320
rect 27068 19168 27120 19174
rect 27068 19110 27120 19116
rect 27080 18834 27108 19110
rect 27068 18828 27120 18834
rect 27068 18770 27120 18776
rect 26884 18692 26936 18698
rect 26884 18634 26936 18640
rect 26976 18692 27028 18698
rect 26976 18634 27028 18640
rect 26988 18086 27016 18634
rect 26976 18080 27028 18086
rect 26976 18022 27028 18028
rect 27448 16658 27476 25230
rect 27528 24676 27580 24682
rect 27528 24618 27580 24624
rect 27540 22166 27568 24618
rect 27528 22160 27580 22166
rect 27528 22102 27580 22108
rect 27620 19984 27672 19990
rect 27620 19926 27672 19932
rect 27528 19168 27580 19174
rect 27528 19110 27580 19116
rect 27540 18766 27568 19110
rect 27528 18760 27580 18766
rect 27528 18702 27580 18708
rect 27632 17678 27660 19926
rect 27816 18358 27844 28358
rect 27988 24064 28040 24070
rect 27988 24006 28040 24012
rect 28000 23730 28028 24006
rect 27988 23724 28040 23730
rect 27988 23666 28040 23672
rect 29564 23322 29592 30194
rect 30392 29850 30420 31282
rect 31312 30190 31340 37062
rect 32128 36576 32180 36582
rect 32128 36518 32180 36524
rect 32140 30734 32168 36518
rect 32404 35624 32456 35630
rect 32404 35566 32456 35572
rect 32128 30728 32180 30734
rect 32128 30670 32180 30676
rect 31300 30184 31352 30190
rect 31300 30126 31352 30132
rect 30380 29844 30432 29850
rect 30380 29786 30432 29792
rect 31208 25152 31260 25158
rect 31208 25094 31260 25100
rect 31220 24750 31248 25094
rect 31208 24744 31260 24750
rect 31208 24686 31260 24692
rect 30656 24608 30708 24614
rect 30656 24550 30708 24556
rect 30472 24132 30524 24138
rect 30472 24074 30524 24080
rect 30484 23866 30512 24074
rect 30472 23860 30524 23866
rect 30472 23802 30524 23808
rect 29552 23316 29604 23322
rect 29552 23258 29604 23264
rect 28264 22092 28316 22098
rect 28264 22034 28316 22040
rect 28276 21690 28304 22034
rect 28264 21684 28316 21690
rect 28264 21626 28316 21632
rect 28540 21140 28592 21146
rect 28540 21082 28592 21088
rect 28552 19360 28580 21082
rect 28632 19848 28684 19854
rect 28632 19790 28684 19796
rect 28644 19514 28672 19790
rect 29920 19712 29972 19718
rect 29920 19654 29972 19660
rect 28632 19508 28684 19514
rect 28632 19450 28684 19456
rect 28724 19508 28776 19514
rect 28724 19450 28776 19456
rect 28552 19332 28672 19360
rect 27804 18352 27856 18358
rect 27804 18294 27856 18300
rect 27816 17746 27844 18294
rect 27988 18148 28040 18154
rect 27988 18090 28040 18096
rect 27804 17740 27856 17746
rect 27804 17682 27856 17688
rect 27620 17672 27672 17678
rect 27620 17614 27672 17620
rect 27436 16652 27488 16658
rect 27436 16594 27488 16600
rect 27160 16040 27212 16046
rect 27160 15982 27212 15988
rect 26884 14816 26936 14822
rect 26884 14758 26936 14764
rect 26896 12753 26924 14758
rect 27172 13938 27200 15982
rect 27436 15972 27488 15978
rect 27436 15914 27488 15920
rect 27448 15502 27476 15914
rect 27436 15496 27488 15502
rect 27436 15438 27488 15444
rect 27344 14952 27396 14958
rect 27344 14894 27396 14900
rect 27252 14340 27304 14346
rect 27252 14282 27304 14288
rect 27264 14074 27292 14282
rect 27252 14068 27304 14074
rect 27252 14010 27304 14016
rect 27356 13938 27384 14894
rect 27160 13932 27212 13938
rect 27160 13874 27212 13880
rect 27344 13932 27396 13938
rect 27344 13874 27396 13880
rect 26882 12744 26938 12753
rect 26882 12679 26938 12688
rect 26792 11824 26844 11830
rect 26792 11766 26844 11772
rect 26974 10296 27030 10305
rect 26974 10231 27030 10240
rect 26700 8900 26752 8906
rect 26700 8842 26752 8848
rect 26608 8628 26660 8634
rect 26608 8570 26660 8576
rect 26240 7404 26292 7410
rect 26240 7346 26292 7352
rect 26516 7404 26568 7410
rect 26516 7346 26568 7352
rect 26252 7206 26280 7346
rect 26240 7200 26292 7206
rect 26238 7168 26240 7177
rect 26332 7200 26384 7206
rect 26292 7168 26294 7177
rect 26332 7142 26384 7148
rect 26238 7103 26294 7112
rect 26240 6996 26292 7002
rect 26240 6938 26292 6944
rect 25964 6928 26016 6934
rect 25964 6870 26016 6876
rect 26148 6860 26200 6866
rect 26148 6802 26200 6808
rect 25964 6112 26016 6118
rect 25964 6054 26016 6060
rect 25976 4026 26004 6054
rect 26056 4072 26108 4078
rect 25976 4020 26056 4026
rect 25976 4014 26108 4020
rect 25976 3998 26096 4014
rect 25964 3936 26016 3942
rect 25964 3878 26016 3884
rect 25976 3466 26004 3878
rect 25872 3460 25924 3466
rect 25872 3402 25924 3408
rect 25964 3460 26016 3466
rect 25964 3402 26016 3408
rect 26160 2990 26188 6802
rect 26252 5710 26280 6938
rect 26344 6798 26372 7142
rect 26988 6934 27016 10231
rect 27172 9926 27200 13874
rect 27448 13462 27476 15438
rect 27620 13728 27672 13734
rect 27620 13670 27672 13676
rect 27632 13530 27660 13670
rect 27620 13524 27672 13530
rect 27620 13466 27672 13472
rect 27436 13456 27488 13462
rect 27436 13398 27488 13404
rect 27620 13320 27672 13326
rect 27620 13262 27672 13268
rect 27250 12744 27306 12753
rect 27250 12679 27306 12688
rect 27160 9920 27212 9926
rect 27160 9862 27212 9868
rect 27264 7954 27292 12679
rect 27632 12434 27660 13262
rect 28000 12782 28028 18090
rect 28540 18080 28592 18086
rect 28540 18022 28592 18028
rect 28172 17536 28224 17542
rect 28172 17478 28224 17484
rect 28184 17202 28212 17478
rect 28172 17196 28224 17202
rect 28172 17138 28224 17144
rect 28552 16522 28580 18022
rect 28172 16516 28224 16522
rect 28172 16458 28224 16464
rect 28540 16516 28592 16522
rect 28540 16458 28592 16464
rect 28184 16250 28212 16458
rect 28172 16244 28224 16250
rect 28172 16186 28224 16192
rect 28264 16244 28316 16250
rect 28264 16186 28316 16192
rect 28184 15706 28212 16186
rect 28276 15910 28304 16186
rect 28540 16040 28592 16046
rect 28540 15982 28592 15988
rect 28356 15972 28408 15978
rect 28356 15914 28408 15920
rect 28264 15904 28316 15910
rect 28264 15846 28316 15852
rect 28172 15700 28224 15706
rect 28172 15642 28224 15648
rect 28368 15502 28396 15914
rect 28552 15706 28580 15982
rect 28540 15700 28592 15706
rect 28540 15642 28592 15648
rect 28356 15496 28408 15502
rect 28356 15438 28408 15444
rect 28264 14340 28316 14346
rect 28264 14282 28316 14288
rect 28276 14074 28304 14282
rect 28264 14068 28316 14074
rect 28264 14010 28316 14016
rect 27988 12776 28040 12782
rect 27988 12718 28040 12724
rect 28172 12776 28224 12782
rect 28172 12718 28224 12724
rect 28184 12442 28212 12718
rect 28172 12436 28224 12442
rect 27632 12406 27844 12434
rect 27620 11688 27672 11694
rect 27620 11630 27672 11636
rect 27344 8492 27396 8498
rect 27344 8434 27396 8440
rect 27252 7948 27304 7954
rect 27252 7890 27304 7896
rect 26976 6928 27028 6934
rect 26976 6870 27028 6876
rect 26700 6860 26752 6866
rect 26700 6802 26752 6808
rect 26332 6792 26384 6798
rect 26332 6734 26384 6740
rect 26606 6760 26662 6769
rect 26606 6695 26662 6704
rect 26330 6624 26386 6633
rect 26330 6559 26386 6568
rect 26344 6118 26372 6559
rect 26516 6248 26568 6254
rect 26516 6190 26568 6196
rect 26332 6112 26384 6118
rect 26332 6054 26384 6060
rect 26332 5908 26384 5914
rect 26332 5850 26384 5856
rect 26240 5704 26292 5710
rect 26240 5646 26292 5652
rect 26240 5568 26292 5574
rect 26344 5545 26372 5850
rect 26424 5704 26476 5710
rect 26424 5646 26476 5652
rect 26240 5510 26292 5516
rect 26330 5536 26386 5545
rect 26252 4690 26280 5510
rect 26330 5471 26386 5480
rect 26436 5409 26464 5646
rect 26422 5400 26478 5409
rect 26422 5335 26478 5344
rect 26240 4684 26292 4690
rect 26240 4626 26292 4632
rect 26424 4616 26476 4622
rect 26238 4584 26294 4593
rect 26238 4519 26294 4528
rect 26422 4584 26424 4593
rect 26476 4584 26478 4593
rect 26422 4519 26478 4528
rect 26252 4486 26280 4519
rect 26240 4480 26292 4486
rect 26240 4422 26292 4428
rect 26424 4004 26476 4010
rect 26424 3946 26476 3952
rect 26240 3460 26292 3466
rect 26240 3402 26292 3408
rect 26252 3369 26280 3402
rect 26238 3360 26294 3369
rect 26238 3295 26294 3304
rect 26238 3224 26294 3233
rect 26238 3159 26240 3168
rect 26292 3159 26294 3168
rect 26240 3130 26292 3136
rect 26148 2984 26200 2990
rect 26148 2926 26200 2932
rect 26436 2922 26464 3946
rect 26528 2961 26556 6190
rect 26620 5914 26648 6695
rect 26608 5908 26660 5914
rect 26608 5850 26660 5856
rect 26712 4758 26740 6802
rect 26790 6488 26846 6497
rect 26790 6423 26846 6432
rect 26804 5234 26832 6423
rect 27158 6352 27214 6361
rect 27356 6338 27384 8434
rect 27436 7744 27488 7750
rect 27436 7686 27488 7692
rect 27264 6322 27384 6338
rect 27158 6287 27160 6296
rect 27212 6287 27214 6296
rect 27252 6316 27384 6322
rect 27160 6258 27212 6264
rect 27304 6310 27384 6316
rect 27252 6258 27304 6264
rect 27448 5710 27476 7686
rect 27528 6384 27580 6390
rect 27632 6361 27660 11630
rect 27816 11286 27844 12406
rect 28172 12378 28224 12384
rect 28276 12170 28304 14010
rect 28368 12345 28396 15438
rect 28448 13728 28500 13734
rect 28448 13670 28500 13676
rect 28354 12336 28410 12345
rect 28354 12271 28410 12280
rect 28356 12232 28408 12238
rect 28356 12174 28408 12180
rect 28264 12164 28316 12170
rect 28264 12106 28316 12112
rect 27896 11824 27948 11830
rect 27896 11766 27948 11772
rect 27908 11354 27936 11766
rect 28368 11558 28396 12174
rect 28356 11552 28408 11558
rect 28356 11494 28408 11500
rect 27896 11348 27948 11354
rect 27896 11290 27948 11296
rect 27804 11280 27856 11286
rect 27804 11222 27856 11228
rect 27712 8356 27764 8362
rect 27712 8298 27764 8304
rect 27528 6326 27580 6332
rect 27618 6352 27674 6361
rect 27540 5914 27568 6326
rect 27618 6287 27674 6296
rect 27528 5908 27580 5914
rect 27528 5850 27580 5856
rect 27160 5704 27212 5710
rect 27160 5646 27212 5652
rect 27436 5704 27488 5710
rect 27436 5646 27488 5652
rect 26792 5228 26844 5234
rect 26792 5170 26844 5176
rect 26792 5024 26844 5030
rect 26792 4966 26844 4972
rect 26700 4752 26752 4758
rect 26700 4694 26752 4700
rect 26804 4690 26832 4966
rect 26884 4752 26936 4758
rect 26884 4694 26936 4700
rect 26792 4684 26844 4690
rect 26792 4626 26844 4632
rect 26896 4282 26924 4694
rect 26884 4276 26936 4282
rect 26884 4218 26936 4224
rect 26976 4276 27028 4282
rect 26976 4218 27028 4224
rect 26792 3936 26844 3942
rect 26792 3878 26844 3884
rect 26700 3664 26752 3670
rect 26700 3606 26752 3612
rect 26514 2952 26570 2961
rect 26424 2916 26476 2922
rect 26514 2887 26570 2896
rect 26424 2858 26476 2864
rect 26436 2825 26464 2858
rect 26422 2816 26478 2825
rect 26422 2751 26478 2760
rect 26436 2514 26464 2751
rect 26712 2650 26740 3606
rect 26804 3602 26832 3878
rect 26792 3596 26844 3602
rect 26792 3538 26844 3544
rect 26882 3496 26938 3505
rect 26988 3482 27016 4218
rect 27172 4146 27200 5646
rect 27528 5024 27580 5030
rect 27528 4966 27580 4972
rect 27540 4214 27568 4966
rect 27528 4208 27580 4214
rect 27528 4150 27580 4156
rect 27618 4176 27674 4185
rect 27160 4140 27212 4146
rect 27618 4111 27674 4120
rect 27160 4082 27212 4088
rect 27632 4078 27660 4111
rect 27620 4072 27672 4078
rect 27620 4014 27672 4020
rect 27528 3732 27580 3738
rect 27528 3674 27580 3680
rect 27252 3664 27304 3670
rect 27080 3612 27252 3618
rect 27080 3606 27304 3612
rect 27080 3602 27292 3606
rect 27068 3596 27292 3602
rect 27120 3590 27292 3596
rect 27068 3538 27120 3544
rect 26938 3454 27016 3482
rect 27066 3496 27122 3505
rect 26882 3431 26938 3440
rect 27066 3431 27068 3440
rect 27120 3431 27122 3440
rect 27344 3460 27396 3466
rect 27068 3402 27120 3408
rect 27396 3420 27476 3448
rect 27344 3402 27396 3408
rect 26976 3120 27028 3126
rect 26976 3062 27028 3068
rect 26988 2922 27016 3062
rect 26976 2916 27028 2922
rect 26976 2858 27028 2864
rect 27080 2836 27108 3402
rect 27250 3360 27306 3369
rect 27250 3295 27306 3304
rect 27264 2990 27292 3295
rect 27448 3194 27476 3420
rect 27436 3188 27488 3194
rect 27436 3130 27488 3136
rect 27344 3120 27396 3126
rect 27342 3088 27344 3097
rect 27396 3088 27398 3097
rect 27342 3023 27398 3032
rect 27252 2984 27304 2990
rect 27252 2926 27304 2932
rect 27344 2984 27396 2990
rect 27344 2926 27396 2932
rect 27356 2836 27384 2926
rect 27080 2808 27384 2836
rect 27540 2774 27568 3674
rect 27620 3120 27672 3126
rect 27620 3062 27672 3068
rect 27448 2746 27568 2774
rect 26608 2644 26660 2650
rect 26608 2586 26660 2592
rect 26700 2644 26752 2650
rect 26700 2586 26752 2592
rect 26620 2514 26648 2586
rect 25964 2508 26016 2514
rect 25700 2468 25964 2496
rect 25136 2450 25188 2456
rect 25964 2450 26016 2456
rect 26424 2508 26476 2514
rect 26424 2450 26476 2456
rect 26608 2508 26660 2514
rect 26608 2450 26660 2456
rect 27160 2440 27212 2446
rect 27160 2382 27212 2388
rect 27172 1970 27200 2382
rect 27160 1964 27212 1970
rect 27160 1906 27212 1912
rect 24952 1896 25004 1902
rect 24952 1838 25004 1844
rect 24860 1760 24912 1766
rect 24860 1702 24912 1708
rect 25780 1760 25832 1766
rect 25780 1702 25832 1708
rect 25792 800 25820 1702
rect 27080 870 27200 898
rect 27080 800 27108 870
rect 13188 734 13492 762
rect 13542 200 13598 800
rect 14830 200 14886 800
rect 16118 200 16174 800
rect 16762 200 16818 800
rect 18050 200 18106 800
rect 19338 200 19394 800
rect 19982 200 20038 800
rect 21270 200 21326 800
rect 22558 200 22614 800
rect 23202 200 23258 800
rect 24490 200 24546 800
rect 25778 200 25834 800
rect 27066 200 27122 800
rect 27172 762 27200 870
rect 27448 762 27476 2746
rect 27632 1766 27660 3062
rect 27724 2446 27752 8298
rect 27816 6458 27844 11222
rect 28460 11218 28488 13670
rect 28644 12434 28672 19332
rect 28736 17202 28764 19450
rect 28908 19372 28960 19378
rect 28908 19314 28960 19320
rect 29092 19372 29144 19378
rect 29092 19314 29144 19320
rect 28920 18290 28948 19314
rect 29000 18760 29052 18766
rect 29000 18702 29052 18708
rect 29012 18290 29040 18702
rect 28908 18284 28960 18290
rect 28908 18226 28960 18232
rect 29000 18284 29052 18290
rect 29000 18226 29052 18232
rect 28920 18193 28948 18226
rect 28906 18184 28962 18193
rect 28906 18119 28962 18128
rect 28724 17196 28776 17202
rect 28724 17138 28776 17144
rect 29000 15360 29052 15366
rect 29000 15302 29052 15308
rect 29012 15026 29040 15302
rect 29104 15026 29132 19314
rect 29368 19168 29420 19174
rect 29368 19110 29420 19116
rect 29380 18358 29408 19110
rect 29368 18352 29420 18358
rect 29368 18294 29420 18300
rect 29828 17128 29880 17134
rect 29828 17070 29880 17076
rect 29840 16658 29868 17070
rect 29828 16652 29880 16658
rect 29828 16594 29880 16600
rect 29932 16522 29960 19654
rect 30104 19372 30156 19378
rect 30104 19314 30156 19320
rect 30116 18426 30144 19314
rect 30196 18624 30248 18630
rect 30196 18566 30248 18572
rect 30104 18420 30156 18426
rect 30104 18362 30156 18368
rect 30208 18290 30236 18566
rect 30196 18284 30248 18290
rect 30196 18226 30248 18232
rect 30208 17338 30236 18226
rect 30564 17808 30616 17814
rect 30564 17750 30616 17756
rect 30196 17332 30248 17338
rect 30196 17274 30248 17280
rect 29920 16516 29972 16522
rect 29920 16458 29972 16464
rect 29276 16040 29328 16046
rect 29276 15982 29328 15988
rect 29000 15020 29052 15026
rect 29000 14962 29052 14968
rect 29092 15020 29144 15026
rect 29092 14962 29144 14968
rect 28816 14816 28868 14822
rect 28816 14758 28868 14764
rect 28828 14414 28856 14758
rect 28816 14408 28868 14414
rect 28816 14350 28868 14356
rect 29104 13258 29132 14962
rect 29288 14958 29316 15982
rect 30196 15972 30248 15978
rect 30196 15914 30248 15920
rect 29920 15904 29972 15910
rect 29920 15846 29972 15852
rect 29932 15502 29960 15846
rect 30208 15638 30236 15914
rect 30196 15632 30248 15638
rect 30196 15574 30248 15580
rect 29920 15496 29972 15502
rect 29920 15438 29972 15444
rect 30472 15020 30524 15026
rect 30472 14962 30524 14968
rect 29276 14952 29328 14958
rect 29276 14894 29328 14900
rect 29920 14816 29972 14822
rect 29920 14758 29972 14764
rect 29736 13864 29788 13870
rect 29736 13806 29788 13812
rect 29748 13530 29776 13806
rect 29736 13524 29788 13530
rect 29736 13466 29788 13472
rect 29932 13326 29960 14758
rect 29184 13320 29236 13326
rect 29184 13262 29236 13268
rect 29920 13320 29972 13326
rect 29920 13262 29972 13268
rect 29092 13252 29144 13258
rect 29092 13194 29144 13200
rect 29196 12986 29224 13262
rect 29368 13184 29420 13190
rect 29368 13126 29420 13132
rect 29184 12980 29236 12986
rect 29184 12922 29236 12928
rect 29380 12714 29408 13126
rect 30484 12850 30512 14962
rect 30472 12844 30524 12850
rect 30472 12786 30524 12792
rect 29368 12708 29420 12714
rect 29368 12650 29420 12656
rect 29000 12640 29052 12646
rect 29000 12582 29052 12588
rect 29012 12434 29040 12582
rect 28644 12406 28856 12434
rect 29012 12406 29132 12434
rect 28448 11212 28500 11218
rect 28448 11154 28500 11160
rect 28448 8492 28500 8498
rect 28448 8434 28500 8440
rect 27896 7404 27948 7410
rect 27896 7346 27948 7352
rect 27804 6452 27856 6458
rect 27804 6394 27856 6400
rect 27908 4729 27936 7346
rect 27986 7168 28042 7177
rect 27986 7103 28042 7112
rect 28000 6798 28028 7103
rect 28460 6798 28488 8434
rect 28630 8392 28686 8401
rect 28630 8327 28632 8336
rect 28684 8327 28686 8336
rect 28632 8298 28684 8304
rect 27988 6792 28040 6798
rect 27988 6734 28040 6740
rect 28448 6792 28500 6798
rect 28448 6734 28500 6740
rect 28000 5710 28028 6734
rect 28264 6112 28316 6118
rect 28264 6054 28316 6060
rect 27988 5704 28040 5710
rect 27988 5646 28040 5652
rect 27988 5568 28040 5574
rect 28172 5568 28224 5574
rect 28040 5528 28120 5556
rect 27988 5510 28040 5516
rect 27894 4720 27950 4729
rect 27804 4684 27856 4690
rect 27894 4655 27950 4664
rect 27804 4626 27856 4632
rect 27816 4554 27844 4626
rect 27804 4548 27856 4554
rect 27804 4490 27856 4496
rect 27988 4208 28040 4214
rect 27988 4150 28040 4156
rect 27896 4140 27948 4146
rect 27896 4082 27948 4088
rect 27712 2440 27764 2446
rect 27712 2382 27764 2388
rect 27712 2304 27764 2310
rect 27712 2246 27764 2252
rect 27620 1760 27672 1766
rect 27620 1702 27672 1708
rect 27724 800 27752 2246
rect 27908 1834 27936 4082
rect 28000 4049 28028 4150
rect 27986 4040 28042 4049
rect 27986 3975 28042 3984
rect 27988 3936 28040 3942
rect 27988 3878 28040 3884
rect 28000 3398 28028 3878
rect 28092 3466 28120 5528
rect 28172 5510 28224 5516
rect 28184 5302 28212 5510
rect 28172 5296 28224 5302
rect 28172 5238 28224 5244
rect 28276 5098 28304 6054
rect 28356 5228 28408 5234
rect 28356 5170 28408 5176
rect 28368 5137 28396 5170
rect 28354 5128 28410 5137
rect 28264 5092 28316 5098
rect 28354 5063 28410 5072
rect 28264 5034 28316 5040
rect 28170 4992 28226 5001
rect 28170 4927 28226 4936
rect 28184 4622 28212 4927
rect 28354 4720 28410 4729
rect 28354 4655 28410 4664
rect 28368 4622 28396 4655
rect 28172 4616 28224 4622
rect 28172 4558 28224 4564
rect 28356 4616 28408 4622
rect 28356 4558 28408 4564
rect 28184 4146 28212 4558
rect 28264 4548 28316 4554
rect 28264 4490 28316 4496
rect 28172 4140 28224 4146
rect 28172 4082 28224 4088
rect 28276 3505 28304 4490
rect 28356 4140 28408 4146
rect 28356 4082 28408 4088
rect 28368 3534 28396 4082
rect 28460 3602 28488 6734
rect 28724 6656 28776 6662
rect 28724 6598 28776 6604
rect 28538 5944 28594 5953
rect 28538 5879 28594 5888
rect 28448 3596 28500 3602
rect 28448 3538 28500 3544
rect 28356 3528 28408 3534
rect 28262 3496 28318 3505
rect 28080 3460 28132 3466
rect 28356 3470 28408 3476
rect 28262 3431 28318 3440
rect 28080 3402 28132 3408
rect 28552 3398 28580 5879
rect 28736 5778 28764 6598
rect 28828 5778 28856 12406
rect 29104 11082 29132 12406
rect 29380 11830 29408 12650
rect 30472 12232 30524 12238
rect 30472 12174 30524 12180
rect 29460 12096 29512 12102
rect 29460 12038 29512 12044
rect 29472 11830 29500 12038
rect 30484 11898 30512 12174
rect 30472 11892 30524 11898
rect 30472 11834 30524 11840
rect 29368 11824 29420 11830
rect 29368 11766 29420 11772
rect 29460 11824 29512 11830
rect 29460 11766 29512 11772
rect 29920 11552 29972 11558
rect 29920 11494 29972 11500
rect 29932 11150 29960 11494
rect 29276 11144 29328 11150
rect 29276 11086 29328 11092
rect 29920 11144 29972 11150
rect 29920 11086 29972 11092
rect 29092 11076 29144 11082
rect 29092 11018 29144 11024
rect 29000 11008 29052 11014
rect 29000 10950 29052 10956
rect 29012 8022 29040 10950
rect 29104 8974 29132 11018
rect 29288 10810 29316 11086
rect 29460 11008 29512 11014
rect 29460 10950 29512 10956
rect 29276 10804 29328 10810
rect 29276 10746 29328 10752
rect 29472 10674 29500 10950
rect 29460 10668 29512 10674
rect 29460 10610 29512 10616
rect 30380 9580 30432 9586
rect 30380 9522 30432 9528
rect 29276 9512 29328 9518
rect 29276 9454 29328 9460
rect 29092 8968 29144 8974
rect 29092 8910 29144 8916
rect 29288 8498 29316 9454
rect 29460 9376 29512 9382
rect 29460 9318 29512 9324
rect 29472 8498 29500 9318
rect 30392 8838 30420 9522
rect 30576 9194 30604 17750
rect 30668 16250 30696 24550
rect 32416 22778 32444 35566
rect 33244 32570 33272 37198
rect 34440 37108 34468 39222
rect 35438 39200 35494 39800
rect 36082 39200 36138 39800
rect 37370 39200 37426 39800
rect 38658 39200 38714 39800
rect 39302 39200 39358 39800
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34520 37120 34572 37126
rect 34440 37080 34520 37108
rect 34520 37062 34572 37068
rect 35452 36786 35480 39200
rect 35992 37256 36044 37262
rect 35992 37198 36044 37204
rect 35440 36780 35492 36786
rect 35440 36722 35492 36728
rect 35900 36780 35952 36786
rect 35900 36722 35952 36728
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 33232 32564 33284 32570
rect 33232 32506 33284 32512
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 35912 31482 35940 36722
rect 36004 33114 36032 37198
rect 36096 37126 36124 39200
rect 37186 38856 37242 38865
rect 37186 38791 37242 38800
rect 36174 37496 36230 37505
rect 36174 37431 36230 37440
rect 36084 37120 36136 37126
rect 36084 37062 36136 37068
rect 36188 36922 36216 37431
rect 36820 37392 36872 37398
rect 36820 37334 36872 37340
rect 36832 36922 36860 37334
rect 36176 36916 36228 36922
rect 36176 36858 36228 36864
rect 36820 36916 36872 36922
rect 36820 36858 36872 36864
rect 36636 36780 36688 36786
rect 36636 36722 36688 36728
rect 36648 36378 36676 36722
rect 36636 36372 36688 36378
rect 36636 36314 36688 36320
rect 37200 36174 37228 38791
rect 37384 36922 37412 39200
rect 38672 37330 38700 39200
rect 39316 37398 39344 39200
rect 39304 37392 39356 37398
rect 39304 37334 39356 37340
rect 38660 37324 38712 37330
rect 38660 37266 38712 37272
rect 37740 37256 37792 37262
rect 37740 37198 37792 37204
rect 37372 36916 37424 36922
rect 37372 36858 37424 36864
rect 37372 36780 37424 36786
rect 37372 36722 37424 36728
rect 36820 36168 36872 36174
rect 36820 36110 36872 36116
rect 37188 36168 37240 36174
rect 37188 36110 37240 36116
rect 36832 35834 36860 36110
rect 37280 36032 37332 36038
rect 37280 35974 37332 35980
rect 36820 35828 36872 35834
rect 36820 35770 36872 35776
rect 35992 33108 36044 33114
rect 35992 33050 36044 33056
rect 37096 31816 37148 31822
rect 37096 31758 37148 31764
rect 35900 31476 35952 31482
rect 35900 31418 35952 31424
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 37108 30938 37136 31758
rect 37096 30932 37148 30938
rect 37096 30874 37148 30880
rect 36176 30728 36228 30734
rect 36176 30670 36228 30676
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34612 27328 34664 27334
rect 34612 27270 34664 27276
rect 33784 26580 33836 26586
rect 33784 26522 33836 26528
rect 32404 22772 32456 22778
rect 32404 22714 32456 22720
rect 30932 22636 30984 22642
rect 30932 22578 30984 22584
rect 30656 16244 30708 16250
rect 30656 16186 30708 16192
rect 30748 15904 30800 15910
rect 30748 15846 30800 15852
rect 30760 15570 30788 15846
rect 30748 15564 30800 15570
rect 30748 15506 30800 15512
rect 30840 13388 30892 13394
rect 30840 13330 30892 13336
rect 30656 13184 30708 13190
rect 30656 13126 30708 13132
rect 30668 12850 30696 13126
rect 30656 12844 30708 12850
rect 30656 12786 30708 12792
rect 30852 11898 30880 13330
rect 30840 11892 30892 11898
rect 30840 11834 30892 11840
rect 30656 11756 30708 11762
rect 30656 11698 30708 11704
rect 30668 11218 30696 11698
rect 30656 11212 30708 11218
rect 30656 11154 30708 11160
rect 30840 9580 30892 9586
rect 30840 9522 30892 9528
rect 30484 9166 30604 9194
rect 30196 8832 30248 8838
rect 30196 8774 30248 8780
rect 30380 8832 30432 8838
rect 30380 8774 30432 8780
rect 29276 8492 29328 8498
rect 29276 8434 29328 8440
rect 29460 8492 29512 8498
rect 29460 8434 29512 8440
rect 29000 8016 29052 8022
rect 29000 7958 29052 7964
rect 29552 7268 29604 7274
rect 29552 7210 29604 7216
rect 28724 5772 28776 5778
rect 28724 5714 28776 5720
rect 28816 5772 28868 5778
rect 28816 5714 28868 5720
rect 29366 5672 29422 5681
rect 29366 5607 29422 5616
rect 28724 5568 28776 5574
rect 28630 5536 28686 5545
rect 28724 5510 28776 5516
rect 28630 5471 28686 5480
rect 28644 5302 28672 5471
rect 28632 5296 28684 5302
rect 28632 5238 28684 5244
rect 28736 4593 28764 5510
rect 29000 5228 29052 5234
rect 29000 5170 29052 5176
rect 29184 5228 29236 5234
rect 29184 5170 29236 5176
rect 28814 4856 28870 4865
rect 28814 4791 28870 4800
rect 28828 4758 28856 4791
rect 28816 4752 28868 4758
rect 28816 4694 28868 4700
rect 28722 4584 28778 4593
rect 28722 4519 28778 4528
rect 28908 4480 28960 4486
rect 28908 4422 28960 4428
rect 28816 3528 28868 3534
rect 28816 3470 28868 3476
rect 28828 3398 28856 3470
rect 27988 3392 28040 3398
rect 27988 3334 28040 3340
rect 28540 3392 28592 3398
rect 28540 3334 28592 3340
rect 28816 3392 28868 3398
rect 28816 3334 28868 3340
rect 28356 3052 28408 3058
rect 28356 2994 28408 3000
rect 28368 2650 28396 2994
rect 28920 2990 28948 4422
rect 29012 4282 29040 5170
rect 29000 4276 29052 4282
rect 29000 4218 29052 4224
rect 29012 4146 29040 4218
rect 29000 4140 29052 4146
rect 29000 4082 29052 4088
rect 29012 3534 29040 4082
rect 29000 3528 29052 3534
rect 29000 3470 29052 3476
rect 29092 3052 29144 3058
rect 29092 2994 29144 3000
rect 28908 2984 28960 2990
rect 28908 2926 28960 2932
rect 28448 2848 28500 2854
rect 28448 2790 28500 2796
rect 28356 2644 28408 2650
rect 28356 2586 28408 2592
rect 28460 2514 28488 2790
rect 28448 2508 28500 2514
rect 28448 2450 28500 2456
rect 29000 2304 29052 2310
rect 29000 2246 29052 2252
rect 27896 1828 27948 1834
rect 27896 1770 27948 1776
rect 29012 800 29040 2246
rect 29104 1630 29132 2994
rect 29196 2689 29224 5170
rect 29276 5024 29328 5030
rect 29276 4966 29328 4972
rect 29288 4690 29316 4966
rect 29276 4684 29328 4690
rect 29276 4626 29328 4632
rect 29274 4040 29330 4049
rect 29274 3975 29330 3984
rect 29288 3738 29316 3975
rect 29276 3732 29328 3738
rect 29276 3674 29328 3680
rect 29182 2680 29238 2689
rect 29182 2615 29238 2624
rect 29380 2446 29408 5607
rect 29460 3732 29512 3738
rect 29460 3674 29512 3680
rect 29472 3398 29500 3674
rect 29460 3392 29512 3398
rect 29460 3334 29512 3340
rect 29564 3058 29592 7210
rect 30208 6322 30236 8774
rect 30392 8634 30420 8774
rect 30380 8628 30432 8634
rect 30380 8570 30432 8576
rect 30484 8362 30512 9166
rect 30852 8974 30880 9522
rect 30840 8968 30892 8974
rect 30840 8910 30892 8916
rect 30472 8356 30524 8362
rect 30472 8298 30524 8304
rect 30484 6866 30512 8298
rect 30472 6860 30524 6866
rect 30472 6802 30524 6808
rect 30196 6316 30248 6322
rect 30196 6258 30248 6264
rect 29734 6216 29790 6225
rect 29734 6151 29790 6160
rect 29642 6080 29698 6089
rect 29642 6015 29698 6024
rect 29656 3398 29684 6015
rect 29748 5710 29776 6151
rect 29918 5808 29974 5817
rect 29918 5743 29974 5752
rect 29736 5704 29788 5710
rect 29736 5646 29788 5652
rect 29828 5568 29880 5574
rect 29828 5510 29880 5516
rect 29736 4140 29788 4146
rect 29736 4082 29788 4088
rect 29748 3913 29776 4082
rect 29734 3904 29790 3913
rect 29734 3839 29790 3848
rect 29840 3670 29868 5510
rect 29828 3664 29880 3670
rect 29828 3606 29880 3612
rect 29644 3392 29696 3398
rect 29644 3334 29696 3340
rect 29932 3058 29960 5743
rect 30378 5264 30434 5273
rect 30378 5199 30380 5208
rect 30432 5199 30434 5208
rect 30380 5170 30432 5176
rect 30012 5092 30064 5098
rect 30012 5034 30064 5040
rect 30024 4826 30052 5034
rect 30564 5024 30616 5030
rect 30564 4966 30616 4972
rect 30012 4820 30064 4826
rect 30012 4762 30064 4768
rect 30380 4616 30432 4622
rect 30380 4558 30432 4564
rect 30392 4321 30420 4558
rect 30470 4448 30526 4457
rect 30470 4383 30526 4392
rect 30378 4312 30434 4321
rect 30378 4247 30434 4256
rect 30484 4146 30512 4383
rect 30012 4140 30064 4146
rect 30012 4082 30064 4088
rect 30472 4140 30524 4146
rect 30472 4082 30524 4088
rect 30024 3942 30052 4082
rect 30012 3936 30064 3942
rect 30012 3878 30064 3884
rect 30288 3936 30340 3942
rect 30288 3878 30340 3884
rect 30300 3777 30328 3878
rect 30286 3768 30342 3777
rect 30286 3703 30342 3712
rect 30472 3392 30524 3398
rect 30472 3334 30524 3340
rect 30484 3233 30512 3334
rect 30470 3224 30526 3233
rect 30470 3159 30526 3168
rect 30380 3120 30432 3126
rect 30378 3088 30380 3097
rect 30432 3088 30434 3097
rect 29552 3052 29604 3058
rect 29552 2994 29604 3000
rect 29920 3052 29972 3058
rect 30378 3023 30434 3032
rect 29920 2994 29972 3000
rect 29736 2848 29788 2854
rect 29736 2790 29788 2796
rect 30380 2848 30432 2854
rect 30380 2790 30432 2796
rect 30472 2848 30524 2854
rect 30472 2790 30524 2796
rect 29748 2553 29776 2790
rect 29734 2544 29790 2553
rect 29734 2479 29790 2488
rect 29368 2440 29420 2446
rect 29368 2382 29420 2388
rect 30288 2304 30340 2310
rect 30288 2246 30340 2252
rect 29092 1624 29144 1630
rect 29092 1566 29144 1572
rect 30300 800 30328 2246
rect 30392 2038 30420 2790
rect 30380 2032 30432 2038
rect 30380 1974 30432 1980
rect 30484 1698 30512 2790
rect 30576 2582 30604 4966
rect 30944 4298 30972 22578
rect 33600 18624 33652 18630
rect 33600 18566 33652 18572
rect 31300 17536 31352 17542
rect 31300 17478 31352 17484
rect 31312 15026 31340 17478
rect 32588 17196 32640 17202
rect 32588 17138 32640 17144
rect 31300 15020 31352 15026
rect 31300 14962 31352 14968
rect 31484 14816 31536 14822
rect 31484 14758 31536 14764
rect 31496 13938 31524 14758
rect 32600 14346 32628 17138
rect 33612 16182 33640 18566
rect 33600 16176 33652 16182
rect 33600 16118 33652 16124
rect 32588 14340 32640 14346
rect 32588 14282 32640 14288
rect 31484 13932 31536 13938
rect 31484 13874 31536 13880
rect 31300 13728 31352 13734
rect 31300 13670 31352 13676
rect 31312 12850 31340 13670
rect 31300 12844 31352 12850
rect 31300 12786 31352 12792
rect 31760 10736 31812 10742
rect 31760 10678 31812 10684
rect 31668 8016 31720 8022
rect 31668 7958 31720 7964
rect 31484 6384 31536 6390
rect 31484 6326 31536 6332
rect 31024 4480 31076 4486
rect 31024 4422 31076 4428
rect 30656 4276 30708 4282
rect 30656 4218 30708 4224
rect 30852 4270 30972 4298
rect 30668 4146 30696 4218
rect 30656 4140 30708 4146
rect 30656 4082 30708 4088
rect 30748 3732 30800 3738
rect 30748 3674 30800 3680
rect 30654 3632 30710 3641
rect 30654 3567 30710 3576
rect 30668 2990 30696 3567
rect 30760 3534 30788 3674
rect 30748 3528 30800 3534
rect 30748 3470 30800 3476
rect 30656 2984 30708 2990
rect 30852 2961 30880 4270
rect 30932 4004 30984 4010
rect 30932 3946 30984 3952
rect 30656 2926 30708 2932
rect 30838 2952 30894 2961
rect 30838 2887 30894 2896
rect 30564 2576 30616 2582
rect 30564 2518 30616 2524
rect 30472 1692 30524 1698
rect 30472 1634 30524 1640
rect 30944 800 30972 3946
rect 31036 2446 31064 4422
rect 31300 3528 31352 3534
rect 31300 3470 31352 3476
rect 31116 3392 31168 3398
rect 31116 3334 31168 3340
rect 31024 2440 31076 2446
rect 31024 2382 31076 2388
rect 31128 2106 31156 3334
rect 31312 2446 31340 3470
rect 31496 3398 31524 6326
rect 31680 4622 31708 7958
rect 31772 4826 31800 10678
rect 31852 5840 31904 5846
rect 31852 5782 31904 5788
rect 31760 4820 31812 4826
rect 31760 4762 31812 4768
rect 31668 4616 31720 4622
rect 31668 4558 31720 4564
rect 31576 4140 31628 4146
rect 31576 4082 31628 4088
rect 31484 3392 31536 3398
rect 31484 3334 31536 3340
rect 31588 3058 31616 4082
rect 31760 3392 31812 3398
rect 31666 3360 31722 3369
rect 31722 3340 31760 3346
rect 31722 3334 31812 3340
rect 31722 3318 31800 3334
rect 31666 3295 31722 3304
rect 31864 3058 31892 5782
rect 32496 4140 32548 4146
rect 32496 4082 32548 4088
rect 32508 4049 32536 4082
rect 32494 4040 32550 4049
rect 32494 3975 32550 3984
rect 32312 3936 32364 3942
rect 32312 3878 32364 3884
rect 32324 3602 32352 3878
rect 32312 3596 32364 3602
rect 32312 3538 32364 3544
rect 31944 3528 31996 3534
rect 31944 3470 31996 3476
rect 31576 3052 31628 3058
rect 31576 2994 31628 3000
rect 31852 3052 31904 3058
rect 31852 2994 31904 3000
rect 31956 2922 31984 3470
rect 32404 3052 32456 3058
rect 32404 2994 32456 3000
rect 31944 2916 31996 2922
rect 31944 2858 31996 2864
rect 31668 2848 31720 2854
rect 32416 2825 32444 2994
rect 31668 2790 31720 2796
rect 32402 2816 32458 2825
rect 31300 2440 31352 2446
rect 31300 2382 31352 2388
rect 31300 2304 31352 2310
rect 31300 2246 31352 2252
rect 31116 2100 31168 2106
rect 31116 2042 31168 2048
rect 31312 1902 31340 2246
rect 31300 1896 31352 1902
rect 31300 1838 31352 1844
rect 31680 1562 31708 2790
rect 32402 2751 32458 2760
rect 32600 2514 32628 14282
rect 33796 12442 33824 26522
rect 34520 26512 34572 26518
rect 34520 26454 34572 26460
rect 34532 25294 34560 26454
rect 34520 25288 34572 25294
rect 34520 25230 34572 25236
rect 34624 23730 34652 27270
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34612 23724 34664 23730
rect 34612 23666 34664 23672
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34796 22024 34848 22030
rect 34796 21966 34848 21972
rect 34704 20256 34756 20262
rect 34704 20198 34756 20204
rect 34716 18766 34744 20198
rect 34704 18760 34756 18766
rect 34704 18702 34756 18708
rect 34808 15978 34836 21966
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35164 18760 35216 18766
rect 35164 18702 35216 18708
rect 35176 18426 35204 18702
rect 35164 18420 35216 18426
rect 35164 18362 35216 18368
rect 35348 18352 35400 18358
rect 35348 18294 35400 18300
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34796 15972 34848 15978
rect 34796 15914 34848 15920
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34428 14816 34480 14822
rect 34428 14758 34480 14764
rect 34440 12850 34468 14758
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34428 12844 34480 12850
rect 34428 12786 34480 12792
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 33784 12436 33836 12442
rect 33784 12378 33836 12384
rect 34520 12436 34572 12442
rect 34520 12378 34572 12384
rect 34060 11756 34112 11762
rect 34060 11698 34112 11704
rect 33140 10600 33192 10606
rect 33140 10542 33192 10548
rect 33152 9654 33180 10542
rect 33140 9648 33192 9654
rect 33140 9590 33192 9596
rect 34072 7546 34100 11698
rect 34532 10674 34560 12378
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34520 10668 34572 10674
rect 34520 10610 34572 10616
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34060 7540 34112 7546
rect 34060 7482 34112 7488
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34612 6248 34664 6254
rect 34612 6190 34664 6196
rect 33416 6112 33468 6118
rect 33416 6054 33468 6060
rect 32956 5160 33008 5166
rect 32956 5102 33008 5108
rect 32968 3738 32996 5102
rect 33048 4548 33100 4554
rect 33048 4490 33100 4496
rect 32956 3732 33008 3738
rect 32956 3674 33008 3680
rect 33060 3194 33088 4490
rect 33048 3188 33100 3194
rect 33048 3130 33100 3136
rect 32588 2508 32640 2514
rect 32588 2450 32640 2456
rect 33428 2446 33456 6054
rect 33508 4480 33560 4486
rect 33508 4422 33560 4428
rect 33600 4480 33652 4486
rect 33600 4422 33652 4428
rect 33520 4146 33548 4422
rect 33612 4214 33640 4422
rect 33600 4208 33652 4214
rect 33600 4150 33652 4156
rect 33508 4140 33560 4146
rect 33508 4082 33560 4088
rect 33784 4004 33836 4010
rect 33784 3946 33836 3952
rect 33796 3534 33824 3946
rect 33784 3528 33836 3534
rect 33784 3470 33836 3476
rect 34624 2922 34652 6190
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34704 4616 34756 4622
rect 34704 4558 34756 4564
rect 34716 3194 34744 4558
rect 34796 3936 34848 3942
rect 34796 3878 34848 3884
rect 34704 3188 34756 3194
rect 34704 3130 34756 3136
rect 34612 2916 34664 2922
rect 34612 2858 34664 2864
rect 34808 2446 34836 3878
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35360 2514 35388 18294
rect 36188 14074 36216 30670
rect 37292 19417 37320 35974
rect 37384 21622 37412 36722
rect 37752 36718 37780 37198
rect 37740 36712 37792 36718
rect 37740 36654 37792 36660
rect 37832 36168 37884 36174
rect 37832 36110 37884 36116
rect 38198 36136 38254 36145
rect 37464 32904 37516 32910
rect 37464 32846 37516 32852
rect 37476 32745 37504 32846
rect 37462 32736 37518 32745
rect 37462 32671 37518 32680
rect 37648 32224 37700 32230
rect 37648 32166 37700 32172
rect 37660 24818 37688 32166
rect 37740 30252 37792 30258
rect 37740 30194 37792 30200
rect 37648 24812 37700 24818
rect 37648 24754 37700 24760
rect 37752 24274 37780 30194
rect 37844 30122 37872 36110
rect 38198 36071 38254 36080
rect 38212 36038 38240 36071
rect 38200 36032 38252 36038
rect 38200 35974 38252 35980
rect 38200 35488 38252 35494
rect 38198 35456 38200 35465
rect 38252 35456 38254 35465
rect 38198 35391 38254 35400
rect 38016 34604 38068 34610
rect 38016 34546 38068 34552
rect 38028 32026 38056 34546
rect 38200 34400 38252 34406
rect 38200 34342 38252 34348
rect 38212 34105 38240 34342
rect 38198 34096 38254 34105
rect 38198 34031 38254 34040
rect 38384 32904 38436 32910
rect 38384 32846 38436 32852
rect 38292 32428 38344 32434
rect 38292 32370 38344 32376
rect 38304 32065 38332 32370
rect 38290 32056 38346 32065
rect 38016 32020 38068 32026
rect 38290 31991 38346 32000
rect 38016 31962 38068 31968
rect 38292 30728 38344 30734
rect 38290 30696 38292 30705
rect 38344 30696 38346 30705
rect 38290 30631 38346 30640
rect 38016 30592 38068 30598
rect 38016 30534 38068 30540
rect 37832 30116 37884 30122
rect 37832 30058 37884 30064
rect 37924 29028 37976 29034
rect 37924 28970 37976 28976
rect 37740 24268 37792 24274
rect 37740 24210 37792 24216
rect 37464 24200 37516 24206
rect 37464 24142 37516 24148
rect 37476 23905 37504 24142
rect 37462 23896 37518 23905
rect 37462 23831 37518 23840
rect 37936 23662 37964 28970
rect 38028 26234 38056 30534
rect 38108 29572 38160 29578
rect 38108 29514 38160 29520
rect 38120 29345 38148 29514
rect 38200 29504 38252 29510
rect 38200 29446 38252 29452
rect 38106 29336 38162 29345
rect 38106 29271 38162 29280
rect 38212 27538 38240 29446
rect 38292 29164 38344 29170
rect 38292 29106 38344 29112
rect 38304 28665 38332 29106
rect 38290 28656 38346 28665
rect 38290 28591 38346 28600
rect 38200 27532 38252 27538
rect 38200 27474 38252 27480
rect 38292 27464 38344 27470
rect 38292 27406 38344 27412
rect 38304 27305 38332 27406
rect 38290 27296 38346 27305
rect 38290 27231 38346 27240
rect 38292 26376 38344 26382
rect 38292 26318 38344 26324
rect 38028 26206 38148 26234
rect 38120 25906 38148 26206
rect 38304 25945 38332 26318
rect 38290 25936 38346 25945
rect 38108 25900 38160 25906
rect 38290 25871 38346 25880
rect 38108 25842 38160 25848
rect 38016 25288 38068 25294
rect 38016 25230 38068 25236
rect 38198 25256 38254 25265
rect 38028 23798 38056 25230
rect 38198 25191 38254 25200
rect 38212 25158 38240 25191
rect 38200 25152 38252 25158
rect 38200 25094 38252 25100
rect 38016 23792 38068 23798
rect 38016 23734 38068 23740
rect 37924 23656 37976 23662
rect 37924 23598 37976 23604
rect 38016 22636 38068 22642
rect 38016 22578 38068 22584
rect 37372 21616 37424 21622
rect 37372 21558 37424 21564
rect 37740 21548 37792 21554
rect 37740 21490 37792 21496
rect 37278 19408 37334 19417
rect 36912 19372 36964 19378
rect 37278 19343 37334 19352
rect 36912 19314 36964 19320
rect 36924 18970 36952 19314
rect 36912 18964 36964 18970
rect 36912 18906 36964 18912
rect 36176 14068 36228 14074
rect 36176 14010 36228 14016
rect 37370 12744 37426 12753
rect 37370 12679 37426 12688
rect 37384 11150 37412 12679
rect 37372 11144 37424 11150
rect 37372 11086 37424 11092
rect 36912 11076 36964 11082
rect 36912 11018 36964 11024
rect 36924 10810 36952 11018
rect 37464 11008 37516 11014
rect 37464 10950 37516 10956
rect 36912 10804 36964 10810
rect 36912 10746 36964 10752
rect 35532 10464 35584 10470
rect 35532 10406 35584 10412
rect 35440 3052 35492 3058
rect 35440 2994 35492 3000
rect 35348 2508 35400 2514
rect 35348 2450 35400 2456
rect 32220 2440 32272 2446
rect 32220 2382 32272 2388
rect 33416 2440 33468 2446
rect 33416 2382 33468 2388
rect 34796 2440 34848 2446
rect 34796 2382 34848 2388
rect 31668 1556 31720 1562
rect 31668 1498 31720 1504
rect 32232 800 32260 2382
rect 33508 2304 33560 2310
rect 33508 2246 33560 2252
rect 34152 2304 34204 2310
rect 34152 2246 34204 2252
rect 33520 800 33548 2246
rect 34164 800 34192 2246
rect 35452 800 35480 2994
rect 35544 2446 35572 10406
rect 37476 10062 37504 10950
rect 37464 10056 37516 10062
rect 37464 9998 37516 10004
rect 37464 7880 37516 7886
rect 37464 7822 37516 7828
rect 37476 7585 37504 7822
rect 37462 7576 37518 7585
rect 37462 7511 37518 7520
rect 35808 7200 35860 7206
rect 35808 7142 35860 7148
rect 35820 6322 35848 7142
rect 35808 6316 35860 6322
rect 35808 6258 35860 6264
rect 37188 3936 37240 3942
rect 37188 3878 37240 3884
rect 37096 2576 37148 2582
rect 37096 2518 37148 2524
rect 35532 2440 35584 2446
rect 35532 2382 35584 2388
rect 36728 2304 36780 2310
rect 36728 2246 36780 2252
rect 36740 800 36768 2246
rect 27172 734 27476 762
rect 27710 200 27766 800
rect 28998 200 29054 800
rect 30286 200 30342 800
rect 30930 200 30986 800
rect 32218 200 32274 800
rect 33506 200 33562 800
rect 34150 200 34206 800
rect 35438 200 35494 800
rect 36726 200 36782 800
rect 37108 105 37136 2518
rect 37200 2145 37228 3878
rect 37752 2514 37780 21490
rect 38028 21146 38056 22578
rect 38198 22536 38254 22545
rect 38198 22471 38200 22480
rect 38252 22471 38254 22480
rect 38200 22442 38252 22448
rect 38200 21888 38252 21894
rect 38198 21856 38200 21865
rect 38252 21856 38254 21865
rect 38198 21791 38254 21800
rect 38016 21140 38068 21146
rect 38016 21082 38068 21088
rect 38396 20942 38424 32846
rect 38384 20936 38436 20942
rect 38384 20878 38436 20884
rect 38290 20496 38346 20505
rect 38290 20431 38292 20440
rect 38344 20431 38346 20440
rect 38292 20402 38344 20408
rect 37832 19780 37884 19786
rect 37832 19722 37884 19728
rect 37844 4826 37872 19722
rect 38200 19168 38252 19174
rect 38198 19136 38200 19145
rect 38252 19136 38254 19145
rect 38198 19071 38254 19080
rect 38396 18902 38424 20878
rect 38384 18896 38436 18902
rect 38384 18838 38436 18844
rect 37924 17264 37976 17270
rect 37924 17206 37976 17212
rect 37832 4820 37884 4826
rect 37832 4762 37884 4768
rect 37936 3058 37964 17206
rect 38198 17096 38254 17105
rect 38198 17031 38200 17040
rect 38252 17031 38254 17040
rect 38200 17002 38252 17008
rect 38016 16448 38068 16454
rect 38016 16390 38068 16396
rect 38028 16114 38056 16390
rect 38016 16108 38068 16114
rect 38016 16050 38068 16056
rect 38200 15904 38252 15910
rect 38200 15846 38252 15852
rect 38212 15745 38240 15846
rect 38198 15736 38254 15745
rect 38198 15671 38254 15680
rect 38108 15428 38160 15434
rect 38108 15370 38160 15376
rect 38120 15065 38148 15370
rect 38200 15360 38252 15366
rect 38200 15302 38252 15308
rect 38106 15056 38162 15065
rect 38106 14991 38162 15000
rect 38212 14482 38240 15302
rect 38200 14476 38252 14482
rect 38200 14418 38252 14424
rect 38016 14272 38068 14278
rect 38016 14214 38068 14220
rect 38028 13938 38056 14214
rect 38016 13932 38068 13938
rect 38016 13874 38068 13880
rect 38200 13728 38252 13734
rect 38198 13696 38200 13705
rect 38252 13696 38254 13705
rect 38198 13631 38254 13640
rect 38200 12640 38252 12646
rect 38200 12582 38252 12588
rect 38212 12345 38240 12582
rect 38198 12336 38254 12345
rect 38198 12271 38254 12280
rect 38200 11280 38252 11286
rect 38200 11222 38252 11228
rect 38212 10985 38240 11222
rect 38198 10976 38254 10985
rect 38198 10911 38254 10920
rect 38016 10668 38068 10674
rect 38016 10610 38068 10616
rect 38028 10266 38056 10610
rect 38200 10464 38252 10470
rect 38200 10406 38252 10412
rect 38212 10305 38240 10406
rect 38198 10296 38254 10305
rect 38016 10260 38068 10266
rect 38198 10231 38254 10240
rect 38016 10202 38068 10208
rect 38292 8968 38344 8974
rect 38290 8936 38292 8945
rect 38344 8936 38346 8945
rect 38290 8871 38346 8880
rect 38108 8832 38160 8838
rect 38108 8774 38160 8780
rect 38120 8498 38148 8774
rect 38108 8492 38160 8498
rect 38108 8434 38160 8440
rect 38292 7404 38344 7410
rect 38292 7346 38344 7352
rect 38304 6905 38332 7346
rect 38290 6896 38346 6905
rect 38290 6831 38346 6840
rect 38016 6112 38068 6118
rect 38016 6054 38068 6060
rect 38028 3534 38056 6054
rect 38200 5568 38252 5574
rect 38198 5536 38200 5545
rect 38252 5536 38254 5545
rect 38198 5471 38254 5480
rect 38108 4548 38160 4554
rect 38108 4490 38160 4496
rect 38120 4185 38148 4490
rect 38106 4176 38162 4185
rect 38106 4111 38162 4120
rect 38016 3528 38068 3534
rect 38016 3470 38068 3476
rect 38198 3496 38254 3505
rect 38198 3431 38254 3440
rect 38212 3398 38240 3431
rect 38200 3392 38252 3398
rect 38200 3334 38252 3340
rect 37832 3052 37884 3058
rect 37832 2994 37884 3000
rect 37924 3052 37976 3058
rect 37924 2994 37976 3000
rect 37740 2508 37792 2514
rect 37740 2450 37792 2456
rect 37372 2440 37424 2446
rect 37372 2382 37424 2388
rect 37186 2136 37242 2145
rect 37186 2071 37242 2080
rect 37384 800 37412 2382
rect 37370 200 37426 800
rect 37844 785 37872 2994
rect 38660 2848 38712 2854
rect 38660 2790 38712 2796
rect 38672 800 38700 2790
rect 37830 776 37886 785
rect 37830 711 37886 720
rect 38658 200 38714 800
rect 37094 96 37150 105
rect 37094 31 37150 40
<< via2 >>
rect 2962 39480 3018 39536
rect 1766 37440 1822 37496
rect 1766 36080 1822 36136
rect 1766 34040 1822 34096
rect 1766 32716 1768 32736
rect 1768 32716 1820 32736
rect 1820 32716 1822 32736
rect 1766 32680 1822 32716
rect 1766 32000 1822 32056
rect 1766 30640 1822 30696
rect 1766 29280 1822 29336
rect 1766 28600 1822 28656
rect 1582 27240 1638 27296
rect 1674 25880 1730 25936
rect 1766 24556 1768 24576
rect 1768 24556 1820 24576
rect 1820 24556 1822 24576
rect 1766 24520 1822 24556
rect 1582 23840 1638 23896
rect 1950 23468 1952 23488
rect 1952 23468 2004 23488
rect 2004 23468 2006 23488
rect 1950 23432 2006 23468
rect 1766 22480 1822 22536
rect 1674 21120 1730 21176
rect 2870 38800 2926 38856
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4526 20712 4582 20768
rect 1582 20440 1638 20496
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 1766 19080 1822 19136
rect 1582 17720 1638 17776
rect 1766 17040 1822 17096
rect 1398 6840 1454 6896
rect 1766 15680 1822 15736
rect 1582 8336 1638 8392
rect 1766 14356 1768 14376
rect 1768 14356 1820 14376
rect 1820 14356 1822 14376
rect 1766 14320 1822 14356
rect 1766 13676 1768 13696
rect 1768 13676 1820 13696
rect 1820 13676 1822 13696
rect 1766 13640 1822 13676
rect 1766 12280 1822 12336
rect 1766 10920 1822 10976
rect 1766 10240 1822 10296
rect 1766 8880 1822 8936
rect 1766 7520 1822 7576
rect 1674 6704 1730 6760
rect 1582 5480 1638 5536
rect 1582 5344 1638 5400
rect 1766 4120 1822 4176
rect 1766 3440 1822 3496
rect 1674 2624 1730 2680
rect 3330 9444 3386 9480
rect 3330 9424 3332 9444
rect 3332 9424 3384 9444
rect 3384 9424 3386 9444
rect 2226 3596 2282 3632
rect 2226 3576 2228 3596
rect 2228 3576 2280 3596
rect 2280 3576 2282 3596
rect 1858 2080 1914 2136
rect 2410 3068 2412 3088
rect 2412 3068 2464 3088
rect 2464 3068 2466 3088
rect 2410 3032 2466 3068
rect 3330 5480 3386 5536
rect 3238 4664 3294 4720
rect 3146 3304 3202 3360
rect 3146 3188 3202 3224
rect 3146 3168 3148 3188
rect 3148 3168 3200 3188
rect 3200 3168 3202 3188
rect 3146 2624 3202 2680
rect 3054 856 3110 912
rect 3698 13776 3754 13832
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4250 17620 4252 17640
rect 4252 17620 4304 17640
rect 4304 17620 4306 17640
rect 4250 17584 4306 17620
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4710 14356 4712 14376
rect 4712 14356 4764 14376
rect 4764 14356 4766 14376
rect 4710 14320 4766 14356
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 3790 9696 3846 9752
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4526 9560 4582 9616
rect 3698 7404 3754 7440
rect 3698 7384 3700 7404
rect 3700 7384 3752 7404
rect 3752 7384 3754 7404
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4066 9016 4122 9072
rect 3790 5208 3846 5264
rect 3790 4120 3846 4176
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4066 7964 4068 7984
rect 4068 7964 4120 7984
rect 4120 7964 4122 7984
rect 4066 7928 4122 7964
rect 4526 7656 4582 7712
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4342 6840 4398 6896
rect 4066 6332 4068 6352
rect 4068 6332 4120 6352
rect 4120 6332 4122 6352
rect 4066 6296 4122 6332
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4894 12824 4950 12880
rect 4802 9716 4858 9752
rect 4802 9696 4804 9716
rect 4804 9696 4856 9716
rect 4856 9696 4858 9716
rect 4526 5108 4528 5128
rect 4528 5108 4580 5128
rect 4580 5108 4582 5128
rect 4526 5072 4582 5108
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 3974 4120 4030 4176
rect 4158 3984 4214 4040
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 5078 13912 5134 13968
rect 5538 12552 5594 12608
rect 5078 7268 5134 7304
rect 5078 7248 5080 7268
rect 5080 7248 5132 7268
rect 5132 7248 5134 7268
rect 5078 6568 5134 6624
rect 5354 7520 5410 7576
rect 6090 14456 6146 14512
rect 6182 12552 6238 12608
rect 5078 4800 5134 4856
rect 4802 4392 4858 4448
rect 4526 3440 4582 3496
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 5722 4528 5778 4584
rect 5998 4664 6054 4720
rect 6274 5908 6330 5944
rect 6274 5888 6276 5908
rect 6276 5888 6328 5908
rect 6328 5888 6330 5908
rect 6182 4256 6238 4312
rect 6458 11228 6460 11248
rect 6460 11228 6512 11248
rect 6512 11228 6514 11248
rect 6458 11192 6514 11228
rect 6550 9696 6606 9752
rect 6918 13932 6974 13968
rect 6918 13912 6920 13932
rect 6920 13912 6972 13932
rect 6972 13912 6974 13932
rect 6826 13504 6882 13560
rect 6826 13368 6882 13424
rect 6642 6024 6698 6080
rect 6550 5616 6606 5672
rect 6918 5752 6974 5808
rect 6826 5344 6882 5400
rect 6918 5208 6974 5264
rect 7010 4120 7066 4176
rect 7194 5344 7250 5400
rect 7194 5244 7196 5264
rect 7196 5244 7248 5264
rect 7248 5244 7250 5264
rect 7194 5208 7250 5244
rect 7562 15428 7618 15464
rect 7562 15408 7564 15428
rect 7564 15408 7616 15428
rect 7616 15408 7618 15428
rect 7838 16632 7894 16688
rect 7838 14320 7894 14376
rect 7378 12708 7434 12744
rect 7378 12688 7380 12708
rect 7380 12688 7432 12708
rect 7432 12688 7434 12708
rect 8022 16360 8078 16416
rect 8022 15564 8078 15600
rect 8022 15544 8024 15564
rect 8024 15544 8076 15564
rect 8076 15544 8078 15564
rect 7562 12416 7618 12472
rect 7930 9152 7986 9208
rect 7562 6840 7618 6896
rect 7470 5344 7526 5400
rect 7838 7420 7840 7440
rect 7840 7420 7892 7440
rect 7892 7420 7894 7440
rect 7838 7384 7894 7420
rect 10506 25744 10562 25800
rect 8482 17448 8538 17504
rect 8298 15544 8354 15600
rect 8482 15580 8484 15600
rect 8484 15580 8536 15600
rect 8536 15580 8538 15600
rect 8482 15544 8538 15580
rect 8482 14492 8484 14512
rect 8484 14492 8536 14512
rect 8536 14492 8538 14512
rect 8114 12416 8170 12472
rect 8482 14456 8538 14492
rect 8574 11192 8630 11248
rect 8390 9152 8446 9208
rect 9126 14320 9182 14376
rect 9126 13524 9182 13560
rect 9126 13504 9128 13524
rect 9128 13504 9180 13524
rect 9180 13504 9182 13524
rect 9586 20712 9642 20768
rect 11058 24248 11114 24304
rect 9770 17196 9826 17232
rect 9770 17176 9772 17196
rect 9772 17176 9824 17196
rect 9824 17176 9826 17196
rect 9678 16904 9734 16960
rect 9770 15680 9826 15736
rect 9126 13096 9182 13152
rect 8850 8608 8906 8664
rect 8298 7656 8354 7712
rect 8390 6704 8446 6760
rect 7930 5752 7986 5808
rect 8390 6432 8446 6488
rect 7930 3848 7986 3904
rect 8666 6568 8722 6624
rect 8666 6180 8722 6216
rect 8666 6160 8668 6180
rect 8668 6160 8720 6180
rect 8720 6160 8722 6180
rect 8482 5788 8484 5808
rect 8484 5788 8536 5808
rect 8536 5788 8538 5808
rect 8482 5752 8538 5788
rect 8298 4120 8354 4176
rect 8390 3440 8446 3496
rect 8574 3304 8630 3360
rect 9586 15580 9588 15600
rect 9588 15580 9640 15600
rect 9640 15580 9642 15600
rect 9586 15544 9642 15580
rect 9770 15428 9826 15464
rect 9770 15408 9772 15428
rect 9772 15408 9824 15428
rect 9824 15408 9826 15428
rect 9770 14456 9826 14512
rect 9586 13096 9642 13152
rect 9678 12824 9734 12880
rect 9770 12416 9826 12472
rect 9678 12144 9734 12200
rect 9494 11736 9550 11792
rect 9862 11620 9918 11656
rect 9862 11600 9864 11620
rect 9864 11600 9916 11620
rect 9916 11600 9918 11620
rect 10230 17040 10286 17096
rect 9586 9716 9642 9752
rect 9586 9696 9588 9716
rect 9588 9696 9640 9716
rect 9640 9696 9642 9716
rect 9494 9036 9550 9072
rect 9494 9016 9496 9036
rect 9496 9016 9548 9036
rect 9548 9016 9550 9036
rect 9586 8880 9642 8936
rect 9770 9868 9772 9888
rect 9772 9868 9824 9888
rect 9824 9868 9826 9888
rect 9770 9832 9826 9868
rect 9770 9560 9826 9616
rect 9402 7248 9458 7304
rect 9586 6160 9642 6216
rect 9218 5480 9274 5536
rect 9126 5072 9182 5128
rect 9126 4664 9182 4720
rect 8850 3848 8906 3904
rect 9494 4256 9550 4312
rect 9494 3732 9550 3768
rect 9494 3712 9496 3732
rect 9496 3712 9548 3732
rect 9548 3712 9550 3732
rect 9402 3460 9458 3496
rect 9402 3440 9404 3460
rect 9404 3440 9456 3460
rect 9456 3440 9458 3460
rect 9954 9988 10010 10024
rect 9954 9968 9956 9988
rect 9956 9968 10008 9988
rect 10008 9968 10010 9988
rect 10230 12688 10286 12744
rect 10874 19372 10930 19408
rect 10874 19352 10876 19372
rect 10876 19352 10928 19372
rect 10928 19352 10930 19372
rect 10598 16768 10654 16824
rect 10414 12316 10416 12336
rect 10416 12316 10468 12336
rect 10468 12316 10470 12336
rect 10414 12280 10470 12316
rect 10230 9832 10286 9888
rect 10414 9560 10470 9616
rect 10874 17040 10930 17096
rect 10874 16652 10930 16688
rect 10874 16632 10876 16652
rect 10876 16632 10928 16652
rect 10928 16632 10930 16652
rect 10966 15000 11022 15056
rect 10690 12552 10746 12608
rect 10966 14456 11022 14512
rect 11242 18944 11298 19000
rect 11334 18400 11390 18456
rect 12070 19236 12126 19272
rect 12070 19216 12072 19236
rect 12072 19216 12124 19236
rect 12124 19216 12126 19236
rect 11702 18708 11704 18728
rect 11704 18708 11756 18728
rect 11756 18708 11758 18728
rect 11702 18672 11758 18708
rect 11794 18420 11850 18456
rect 11794 18400 11796 18420
rect 11796 18400 11848 18420
rect 11848 18400 11850 18420
rect 11702 18128 11758 18184
rect 11334 17584 11390 17640
rect 11610 16904 11666 16960
rect 10782 10784 10838 10840
rect 10598 9968 10654 10024
rect 10230 7520 10286 7576
rect 10322 6432 10378 6488
rect 9954 6024 10010 6080
rect 9954 4392 10010 4448
rect 10230 6160 10286 6216
rect 11518 13912 11574 13968
rect 11426 12552 11482 12608
rect 11426 12280 11482 12336
rect 11978 15544 12034 15600
rect 11886 14864 11942 14920
rect 11794 13912 11850 13968
rect 11886 13776 11942 13832
rect 11518 11872 11574 11928
rect 10598 5480 10654 5536
rect 10506 5208 10562 5264
rect 10690 3732 10746 3768
rect 10690 3712 10692 3732
rect 10692 3712 10744 3732
rect 10744 3712 10746 3732
rect 11150 6840 11206 6896
rect 11150 5616 11206 5672
rect 12622 19352 12678 19408
rect 12622 19216 12678 19272
rect 12346 17312 12402 17368
rect 12254 17040 12310 17096
rect 12990 20984 13046 21040
rect 12346 15408 12402 15464
rect 12346 13912 12402 13968
rect 11794 11736 11850 11792
rect 11334 6024 11390 6080
rect 11886 6976 11942 7032
rect 13174 21256 13230 21312
rect 13266 20712 13322 20768
rect 12990 19080 13046 19136
rect 12530 15036 12532 15056
rect 12532 15036 12584 15056
rect 12584 15036 12586 15056
rect 12530 15000 12586 15036
rect 12530 13368 12586 13424
rect 12806 15272 12862 15328
rect 12806 12688 12862 12744
rect 12530 12144 12586 12200
rect 12438 11600 12494 11656
rect 12990 15408 13046 15464
rect 13082 15136 13138 15192
rect 12990 13640 13046 13696
rect 12898 11464 12954 11520
rect 12438 10920 12494 10976
rect 12254 9016 12310 9072
rect 12438 8744 12494 8800
rect 12346 8508 12348 8528
rect 12348 8508 12400 8528
rect 12400 8508 12402 8528
rect 12346 8472 12402 8508
rect 12162 7112 12218 7168
rect 12162 6840 12218 6896
rect 12070 6704 12126 6760
rect 12254 5888 12310 5944
rect 12346 5616 12402 5672
rect 12070 4936 12126 4992
rect 13174 12416 13230 12472
rect 13082 9596 13084 9616
rect 13084 9596 13136 9616
rect 13136 9596 13138 9616
rect 13082 9560 13138 9596
rect 13726 17312 13782 17368
rect 13450 15988 13452 16008
rect 13452 15988 13504 16008
rect 13504 15988 13506 16008
rect 13450 15952 13506 15988
rect 13542 15136 13598 15192
rect 13634 13640 13690 13696
rect 13818 15408 13874 15464
rect 14370 21120 14426 21176
rect 14278 20304 14334 20360
rect 14094 16088 14150 16144
rect 14094 15544 14150 15600
rect 13818 14864 13874 14920
rect 13450 11736 13506 11792
rect 12806 5344 12862 5400
rect 13266 4936 13322 4992
rect 12990 4800 13046 4856
rect 12530 4256 12586 4312
rect 12622 3304 12678 3360
rect 11886 3032 11942 3088
rect 11978 2916 12034 2952
rect 11978 2896 11980 2916
rect 11980 2896 12032 2916
rect 12032 2896 12034 2916
rect 11058 2216 11114 2272
rect 12622 2760 12678 2816
rect 14278 17448 14334 17504
rect 15382 21972 15384 21992
rect 15384 21972 15436 21992
rect 15436 21972 15438 21992
rect 15382 21936 15438 21972
rect 14094 11228 14096 11248
rect 14096 11228 14148 11248
rect 14148 11228 14150 11248
rect 14094 11192 14150 11228
rect 13542 9424 13598 9480
rect 15658 23432 15714 23488
rect 15750 21936 15806 21992
rect 15842 21800 15898 21856
rect 14830 15272 14886 15328
rect 15014 13912 15070 13968
rect 13634 8508 13636 8528
rect 13636 8508 13688 8528
rect 13688 8508 13690 8528
rect 13634 8472 13690 8508
rect 13358 2796 13360 2816
rect 13360 2796 13412 2816
rect 13412 2796 13414 2816
rect 13358 2760 13414 2796
rect 14370 6704 14426 6760
rect 14646 5752 14702 5808
rect 14646 5072 14702 5128
rect 14646 4528 14702 4584
rect 14830 4548 14886 4584
rect 14830 4528 14832 4548
rect 14832 4528 14884 4548
rect 14884 4528 14886 4548
rect 13634 3032 13690 3088
rect 14554 3984 14610 4040
rect 14830 3032 14886 3088
rect 15382 15408 15438 15464
rect 15290 11192 15346 11248
rect 15106 8608 15162 8664
rect 15934 19372 15990 19408
rect 15934 19352 15936 19372
rect 15936 19352 15988 19372
rect 15988 19352 15990 19372
rect 15842 18264 15898 18320
rect 16118 17584 16174 17640
rect 15658 13504 15714 13560
rect 15566 12008 15622 12064
rect 15750 8744 15806 8800
rect 15658 7384 15714 7440
rect 15106 5480 15162 5536
rect 15106 3168 15162 3224
rect 14462 2624 14518 2680
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 16946 21004 17002 21040
rect 16946 20984 16948 21004
rect 16948 20984 17000 21004
rect 17000 20984 17002 21004
rect 16118 14320 16174 14376
rect 17406 20984 17462 21040
rect 16670 18944 16726 19000
rect 16578 16088 16634 16144
rect 16302 14320 16358 14376
rect 16302 10784 16358 10840
rect 16302 9016 16358 9072
rect 16578 9016 16634 9072
rect 17130 15544 17186 15600
rect 16946 12688 17002 12744
rect 17958 21292 17960 21312
rect 17960 21292 18012 21312
rect 18012 21292 18014 21312
rect 17958 21256 18014 21292
rect 18326 23976 18382 24032
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 18602 21800 18658 21856
rect 16394 7112 16450 7168
rect 16026 5208 16082 5264
rect 16026 4528 16082 4584
rect 16210 4120 16266 4176
rect 16302 3848 16358 3904
rect 17958 17076 17960 17096
rect 17960 17076 18012 17096
rect 18012 17076 18014 17096
rect 17958 17040 18014 17076
rect 17958 15428 18014 15464
rect 17958 15408 17960 15428
rect 17960 15408 18012 15428
rect 18012 15408 18014 15428
rect 18602 21020 18604 21040
rect 18604 21020 18656 21040
rect 18656 21020 18658 21040
rect 18602 20984 18658 21020
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 18418 17176 18474 17232
rect 18142 14184 18198 14240
rect 18234 13776 18290 13832
rect 18694 15680 18750 15736
rect 17866 10124 17922 10160
rect 17866 10104 17868 10124
rect 17868 10104 17920 10124
rect 17920 10104 17922 10124
rect 17406 6976 17462 7032
rect 18602 12008 18658 12064
rect 18418 6024 18474 6080
rect 18234 5616 18290 5672
rect 18234 4004 18290 4040
rect 18234 3984 18236 4004
rect 18236 3984 18288 4004
rect 18288 3984 18290 4004
rect 18418 3596 18474 3632
rect 18418 3576 18420 3596
rect 18420 3576 18472 3596
rect 18472 3576 18474 3596
rect 18878 12416 18934 12472
rect 18786 9560 18842 9616
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 20258 18708 20260 18728
rect 20260 18708 20312 18728
rect 20312 18708 20314 18728
rect 20258 18672 20314 18708
rect 19982 17584 20038 17640
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19614 17076 19616 17096
rect 19616 17076 19668 17096
rect 19668 17076 19670 17096
rect 19614 17040 19670 17076
rect 19522 16632 19578 16688
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19338 15544 19394 15600
rect 19522 15408 19578 15464
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 20074 15000 20130 15056
rect 19522 14592 19578 14648
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19706 13252 19762 13288
rect 19706 13232 19708 13252
rect 19708 13232 19760 13252
rect 19760 13232 19762 13252
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19982 12980 20038 13016
rect 19982 12960 19984 12980
rect 19984 12960 20036 12980
rect 20036 12960 20038 12980
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 20534 17992 20590 18048
rect 20718 17040 20774 17096
rect 20810 16496 20866 16552
rect 20534 15408 20590 15464
rect 20626 15136 20682 15192
rect 20442 14456 20498 14512
rect 20442 14184 20498 14240
rect 20626 12280 20682 12336
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19982 7384 20038 7440
rect 19614 7284 19616 7304
rect 19616 7284 19668 7304
rect 19668 7284 19670 7304
rect 19614 7248 19670 7284
rect 19614 6740 19616 6760
rect 19616 6740 19668 6760
rect 19668 6740 19670 6760
rect 19614 6704 19670 6740
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19706 6296 19762 6352
rect 20074 5480 20130 5536
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 20718 8880 20774 8936
rect 22006 21120 22062 21176
rect 22742 20984 22798 21040
rect 21546 12416 21602 12472
rect 21086 7248 21142 7304
rect 20810 6704 20866 6760
rect 20534 5344 20590 5400
rect 18878 4156 18880 4176
rect 18880 4156 18932 4176
rect 18932 4156 18934 4176
rect 18878 4120 18934 4156
rect 19522 4800 19578 4856
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 20258 4256 20314 4312
rect 20074 3848 20130 3904
rect 19338 3712 19394 3768
rect 19982 3712 20038 3768
rect 19338 3576 19394 3632
rect 19522 3576 19578 3632
rect 19292 3440 19348 3496
rect 19614 3440 19670 3496
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19614 3032 19670 3088
rect 19338 2488 19394 2544
rect 21178 6704 21234 6760
rect 21270 6296 21326 6352
rect 21178 6024 21234 6080
rect 20994 4120 21050 4176
rect 21546 6724 21602 6760
rect 21546 6704 21548 6724
rect 21548 6704 21600 6724
rect 21600 6704 21602 6724
rect 22098 12144 22154 12200
rect 21822 6432 21878 6488
rect 21546 5616 21602 5672
rect 21730 5480 21786 5536
rect 21454 4392 21510 4448
rect 21454 4120 21510 4176
rect 21638 4120 21694 4176
rect 20534 3576 20590 3632
rect 22466 16088 22522 16144
rect 23754 21020 23756 21040
rect 23756 21020 23808 21040
rect 23808 21020 23810 21040
rect 23754 20984 23810 21020
rect 23386 16532 23388 16552
rect 23388 16532 23440 16552
rect 23440 16532 23442 16552
rect 23386 16496 23442 16532
rect 22650 12824 22706 12880
rect 22374 7928 22430 7984
rect 22006 6604 22008 6624
rect 22008 6604 22060 6624
rect 22060 6604 22062 6624
rect 22006 6568 22062 6604
rect 22006 5752 22062 5808
rect 21914 5480 21970 5536
rect 21914 4936 21970 4992
rect 21914 4800 21970 4856
rect 21822 3984 21878 4040
rect 20258 2760 20314 2816
rect 19614 2488 19670 2544
rect 19522 2352 19578 2408
rect 19706 2372 19762 2408
rect 22466 5516 22468 5536
rect 22468 5516 22520 5536
rect 22520 5516 22522 5536
rect 22466 5480 22522 5516
rect 23202 14592 23258 14648
rect 23110 12824 23166 12880
rect 23018 12144 23074 12200
rect 22742 5752 22798 5808
rect 22466 3712 22522 3768
rect 22742 2488 22798 2544
rect 19706 2352 19708 2372
rect 19708 2352 19760 2372
rect 19760 2352 19762 2372
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 21914 2352 21970 2408
rect 23478 12416 23534 12472
rect 23294 12164 23350 12200
rect 23294 12144 23296 12164
rect 23296 12144 23348 12164
rect 23348 12144 23350 12164
rect 23386 12008 23442 12064
rect 23754 7928 23810 7984
rect 23478 6568 23534 6624
rect 23294 6432 23350 6488
rect 24398 13404 24400 13424
rect 24400 13404 24452 13424
rect 24452 13404 24454 13424
rect 24398 13368 24454 13404
rect 24214 11636 24216 11656
rect 24216 11636 24268 11656
rect 24268 11636 24270 11656
rect 24214 11600 24270 11636
rect 24030 9460 24032 9480
rect 24032 9460 24084 9480
rect 24084 9460 24086 9480
rect 23846 4392 23902 4448
rect 23386 3712 23442 3768
rect 23294 3304 23350 3360
rect 24030 9424 24086 9460
rect 24030 5480 24086 5536
rect 24214 7112 24270 7168
rect 24490 12044 24492 12064
rect 24492 12044 24544 12064
rect 24544 12044 24546 12064
rect 24490 12008 24546 12044
rect 24674 10124 24730 10160
rect 24674 10104 24676 10124
rect 24676 10104 24728 10124
rect 24728 10104 24730 10124
rect 24858 7112 24914 7168
rect 24582 4936 24638 4992
rect 24766 4548 24822 4584
rect 24766 4528 24768 4548
rect 24768 4528 24820 4548
rect 24820 4528 24822 4548
rect 24122 4020 24124 4040
rect 24124 4020 24176 4040
rect 24176 4020 24178 4040
rect 24122 3984 24178 4020
rect 25594 13232 25650 13288
rect 24950 6568 25006 6624
rect 25042 4800 25098 4856
rect 25502 4392 25558 4448
rect 24766 3984 24822 4040
rect 25686 5636 25742 5672
rect 25686 5616 25688 5636
rect 25688 5616 25740 5636
rect 25740 5616 25742 5636
rect 24674 3460 24730 3496
rect 24674 3440 24676 3460
rect 24676 3440 24728 3460
rect 24728 3440 24730 3460
rect 26882 12688 26938 12744
rect 26974 10240 27030 10296
rect 26238 7148 26240 7168
rect 26240 7148 26292 7168
rect 26292 7148 26294 7168
rect 26238 7112 26294 7148
rect 27250 12688 27306 12744
rect 26606 6704 26662 6760
rect 26330 6568 26386 6624
rect 26330 5480 26386 5536
rect 26422 5344 26478 5400
rect 26238 4528 26294 4584
rect 26422 4564 26424 4584
rect 26424 4564 26476 4584
rect 26476 4564 26478 4584
rect 26422 4528 26478 4564
rect 26238 3304 26294 3360
rect 26238 3188 26294 3224
rect 26238 3168 26240 3188
rect 26240 3168 26292 3188
rect 26292 3168 26294 3188
rect 26790 6432 26846 6488
rect 27158 6316 27214 6352
rect 27158 6296 27160 6316
rect 27160 6296 27212 6316
rect 27212 6296 27214 6316
rect 28354 12280 28410 12336
rect 27618 6296 27674 6352
rect 26514 2896 26570 2952
rect 26422 2760 26478 2816
rect 26882 3440 26938 3496
rect 27618 4120 27674 4176
rect 27066 3460 27122 3496
rect 27066 3440 27068 3460
rect 27068 3440 27120 3460
rect 27120 3440 27122 3460
rect 27250 3304 27306 3360
rect 27342 3068 27344 3088
rect 27344 3068 27396 3088
rect 27396 3068 27398 3088
rect 27342 3032 27398 3068
rect 28906 18128 28962 18184
rect 27986 7112 28042 7168
rect 28630 8356 28686 8392
rect 28630 8336 28632 8356
rect 28632 8336 28684 8356
rect 28684 8336 28686 8356
rect 27894 4664 27950 4720
rect 27986 3984 28042 4040
rect 28354 5072 28410 5128
rect 28170 4936 28226 4992
rect 28354 4664 28410 4720
rect 28538 5888 28594 5944
rect 28262 3440 28318 3496
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 37186 38800 37242 38856
rect 36174 37440 36230 37496
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 29366 5616 29422 5672
rect 28630 5480 28686 5536
rect 28814 4800 28870 4856
rect 28722 4528 28778 4584
rect 29274 3984 29330 4040
rect 29182 2624 29238 2680
rect 29734 6160 29790 6216
rect 29642 6024 29698 6080
rect 29918 5752 29974 5808
rect 29734 3848 29790 3904
rect 30378 5228 30434 5264
rect 30378 5208 30380 5228
rect 30380 5208 30432 5228
rect 30432 5208 30434 5228
rect 30470 4392 30526 4448
rect 30378 4256 30434 4312
rect 30286 3712 30342 3768
rect 30470 3168 30526 3224
rect 30378 3068 30380 3088
rect 30380 3068 30432 3088
rect 30432 3068 30434 3088
rect 30378 3032 30434 3068
rect 29734 2488 29790 2544
rect 30654 3576 30710 3632
rect 30838 2896 30894 2952
rect 31666 3304 31722 3360
rect 32494 3984 32550 4040
rect 32402 2760 32458 2816
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 37462 32680 37518 32736
rect 38198 36080 38254 36136
rect 38198 35436 38200 35456
rect 38200 35436 38252 35456
rect 38252 35436 38254 35456
rect 38198 35400 38254 35436
rect 38198 34040 38254 34096
rect 38290 32000 38346 32056
rect 38290 30676 38292 30696
rect 38292 30676 38344 30696
rect 38344 30676 38346 30696
rect 38290 30640 38346 30676
rect 37462 23840 37518 23896
rect 38106 29280 38162 29336
rect 38290 28600 38346 28656
rect 38290 27240 38346 27296
rect 38290 25880 38346 25936
rect 38198 25200 38254 25256
rect 37278 19352 37334 19408
rect 37370 12688 37426 12744
rect 37462 7520 37518 7576
rect 38198 22500 38254 22536
rect 38198 22480 38200 22500
rect 38200 22480 38252 22500
rect 38252 22480 38254 22500
rect 38198 21836 38200 21856
rect 38200 21836 38252 21856
rect 38252 21836 38254 21856
rect 38198 21800 38254 21836
rect 38290 20460 38346 20496
rect 38290 20440 38292 20460
rect 38292 20440 38344 20460
rect 38344 20440 38346 20460
rect 38198 19116 38200 19136
rect 38200 19116 38252 19136
rect 38252 19116 38254 19136
rect 38198 19080 38254 19116
rect 38198 17060 38254 17096
rect 38198 17040 38200 17060
rect 38200 17040 38252 17060
rect 38252 17040 38254 17060
rect 38198 15680 38254 15736
rect 38106 15000 38162 15056
rect 38198 13676 38200 13696
rect 38200 13676 38252 13696
rect 38252 13676 38254 13696
rect 38198 13640 38254 13676
rect 38198 12280 38254 12336
rect 38198 10920 38254 10976
rect 38198 10240 38254 10296
rect 38290 8916 38292 8936
rect 38292 8916 38344 8936
rect 38344 8916 38346 8936
rect 38290 8880 38346 8916
rect 38290 6840 38346 6896
rect 38198 5516 38200 5536
rect 38200 5516 38252 5536
rect 38252 5516 38254 5536
rect 38198 5480 38254 5516
rect 38106 4120 38162 4176
rect 38198 3440 38254 3496
rect 37186 2080 37242 2136
rect 37830 720 37886 776
rect 37094 40 37150 96
<< metal3 >>
rect 200 39538 800 39568
rect 2957 39538 3023 39541
rect 200 39536 3023 39538
rect 200 39480 2962 39536
rect 3018 39480 3023 39536
rect 200 39478 3023 39480
rect 200 39448 800 39478
rect 2957 39475 3023 39478
rect 200 38858 800 38888
rect 2865 38858 2931 38861
rect 200 38856 2931 38858
rect 200 38800 2870 38856
rect 2926 38800 2931 38856
rect 200 38798 2931 38800
rect 200 38768 800 38798
rect 2865 38795 2931 38798
rect 37181 38858 37247 38861
rect 39200 38858 39800 38888
rect 37181 38856 39800 38858
rect 37181 38800 37186 38856
rect 37242 38800 39800 38856
rect 37181 38798 39800 38800
rect 37181 38795 37247 38798
rect 39200 38768 39800 38798
rect 4210 37568 4526 37569
rect 200 37498 800 37528
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 1761 37498 1827 37501
rect 200 37496 1827 37498
rect 200 37440 1766 37496
rect 1822 37440 1827 37496
rect 200 37438 1827 37440
rect 200 37408 800 37438
rect 1761 37435 1827 37438
rect 36169 37498 36235 37501
rect 39200 37498 39800 37528
rect 36169 37496 39800 37498
rect 36169 37440 36174 37496
rect 36230 37440 39800 37496
rect 36169 37438 39800 37440
rect 36169 37435 36235 37438
rect 39200 37408 39800 37438
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 200 36138 800 36168
rect 1761 36138 1827 36141
rect 200 36136 1827 36138
rect 200 36080 1766 36136
rect 1822 36080 1827 36136
rect 200 36078 1827 36080
rect 200 36048 800 36078
rect 1761 36075 1827 36078
rect 38193 36138 38259 36141
rect 39200 36138 39800 36168
rect 38193 36136 39800 36138
rect 38193 36080 38198 36136
rect 38254 36080 39800 36136
rect 38193 36078 39800 36080
rect 38193 36075 38259 36078
rect 39200 36048 39800 36078
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 200 35368 800 35488
rect 38193 35458 38259 35461
rect 39200 35458 39800 35488
rect 38193 35456 39800 35458
rect 38193 35400 38198 35456
rect 38254 35400 39800 35456
rect 38193 35398 39800 35400
rect 38193 35395 38259 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 39200 35368 39800 35398
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 200 34098 800 34128
rect 1761 34098 1827 34101
rect 200 34096 1827 34098
rect 200 34040 1766 34096
rect 1822 34040 1827 34096
rect 200 34038 1827 34040
rect 200 34008 800 34038
rect 1761 34035 1827 34038
rect 38193 34098 38259 34101
rect 39200 34098 39800 34128
rect 38193 34096 39800 34098
rect 38193 34040 38198 34096
rect 38254 34040 39800 34096
rect 38193 34038 39800 34040
rect 38193 34035 38259 34038
rect 39200 34008 39800 34038
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 200 32738 800 32768
rect 1761 32738 1827 32741
rect 200 32736 1827 32738
rect 200 32680 1766 32736
rect 1822 32680 1827 32736
rect 200 32678 1827 32680
rect 200 32648 800 32678
rect 1761 32675 1827 32678
rect 37457 32738 37523 32741
rect 39200 32738 39800 32768
rect 37457 32736 39800 32738
rect 37457 32680 37462 32736
rect 37518 32680 39800 32736
rect 37457 32678 39800 32680
rect 37457 32675 37523 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 39200 32648 39800 32678
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 200 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 1761 32058 1827 32061
rect 200 32056 1827 32058
rect 200 32000 1766 32056
rect 1822 32000 1827 32056
rect 200 31998 1827 32000
rect 200 31968 800 31998
rect 1761 31995 1827 31998
rect 38285 32058 38351 32061
rect 39200 32058 39800 32088
rect 38285 32056 39800 32058
rect 38285 32000 38290 32056
rect 38346 32000 39800 32056
rect 38285 31998 39800 32000
rect 38285 31995 38351 31998
rect 39200 31968 39800 31998
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 200 30698 800 30728
rect 1761 30698 1827 30701
rect 200 30696 1827 30698
rect 200 30640 1766 30696
rect 1822 30640 1827 30696
rect 200 30638 1827 30640
rect 200 30608 800 30638
rect 1761 30635 1827 30638
rect 38285 30698 38351 30701
rect 39200 30698 39800 30728
rect 38285 30696 39800 30698
rect 38285 30640 38290 30696
rect 38346 30640 39800 30696
rect 38285 30638 39800 30640
rect 38285 30635 38351 30638
rect 39200 30608 39800 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 200 29338 800 29368
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 1761 29338 1827 29341
rect 200 29336 1827 29338
rect 200 29280 1766 29336
rect 1822 29280 1827 29336
rect 200 29278 1827 29280
rect 200 29248 800 29278
rect 1761 29275 1827 29278
rect 38101 29338 38167 29341
rect 39200 29338 39800 29368
rect 38101 29336 39800 29338
rect 38101 29280 38106 29336
rect 38162 29280 39800 29336
rect 38101 29278 39800 29280
rect 38101 29275 38167 29278
rect 39200 29248 39800 29278
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 200 28658 800 28688
rect 1761 28658 1827 28661
rect 200 28656 1827 28658
rect 200 28600 1766 28656
rect 1822 28600 1827 28656
rect 200 28598 1827 28600
rect 200 28568 800 28598
rect 1761 28595 1827 28598
rect 38285 28658 38351 28661
rect 39200 28658 39800 28688
rect 38285 28656 39800 28658
rect 38285 28600 38290 28656
rect 38346 28600 39800 28656
rect 38285 28598 39800 28600
rect 38285 28595 38351 28598
rect 39200 28568 39800 28598
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 200 27298 800 27328
rect 1577 27298 1643 27301
rect 200 27296 1643 27298
rect 200 27240 1582 27296
rect 1638 27240 1643 27296
rect 200 27238 1643 27240
rect 200 27208 800 27238
rect 1577 27235 1643 27238
rect 38285 27298 38351 27301
rect 39200 27298 39800 27328
rect 38285 27296 39800 27298
rect 38285 27240 38290 27296
rect 38346 27240 39800 27296
rect 38285 27238 39800 27240
rect 38285 27235 38351 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 39200 27208 39800 27238
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 200 25938 800 25968
rect 1669 25938 1735 25941
rect 200 25936 1735 25938
rect 200 25880 1674 25936
rect 1730 25880 1735 25936
rect 200 25878 1735 25880
rect 200 25848 800 25878
rect 1669 25875 1735 25878
rect 38285 25938 38351 25941
rect 39200 25938 39800 25968
rect 38285 25936 39800 25938
rect 38285 25880 38290 25936
rect 38346 25880 39800 25936
rect 38285 25878 39800 25880
rect 38285 25875 38351 25878
rect 39200 25848 39800 25878
rect 10501 25804 10567 25805
rect 10501 25802 10548 25804
rect 10456 25800 10548 25802
rect 10456 25744 10506 25800
rect 10456 25742 10548 25744
rect 10501 25740 10548 25742
rect 10612 25740 10618 25804
rect 10501 25739 10567 25740
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 38193 25258 38259 25261
rect 39200 25258 39800 25288
rect 38193 25256 39800 25258
rect 38193 25200 38198 25256
rect 38254 25200 39800 25256
rect 38193 25198 39800 25200
rect 38193 25195 38259 25198
rect 39200 25168 39800 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 200 24578 800 24608
rect 1761 24578 1827 24581
rect 200 24576 1827 24578
rect 200 24520 1766 24576
rect 1822 24520 1827 24576
rect 200 24518 1827 24520
rect 200 24488 800 24518
rect 1761 24515 1827 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 3182 24244 3188 24308
rect 3252 24306 3258 24308
rect 11053 24306 11119 24309
rect 3252 24304 11119 24306
rect 3252 24248 11058 24304
rect 11114 24248 11119 24304
rect 3252 24246 11119 24248
rect 3252 24244 3258 24246
rect 11053 24243 11119 24246
rect 18321 24034 18387 24037
rect 18454 24034 18460 24036
rect 18321 24032 18460 24034
rect 18321 23976 18326 24032
rect 18382 23976 18460 24032
rect 18321 23974 18460 23976
rect 18321 23971 18387 23974
rect 18454 23972 18460 23974
rect 18524 23972 18530 24036
rect 19570 23968 19886 23969
rect 200 23898 800 23928
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 1577 23898 1643 23901
rect 200 23896 1643 23898
rect 200 23840 1582 23896
rect 1638 23840 1643 23896
rect 200 23838 1643 23840
rect 200 23808 800 23838
rect 1577 23835 1643 23838
rect 37457 23898 37523 23901
rect 39200 23898 39800 23928
rect 37457 23896 39800 23898
rect 37457 23840 37462 23896
rect 37518 23840 39800 23896
rect 37457 23838 39800 23840
rect 37457 23835 37523 23838
rect 39200 23808 39800 23838
rect 1710 23428 1716 23492
rect 1780 23490 1786 23492
rect 1945 23490 2011 23493
rect 1780 23488 2011 23490
rect 1780 23432 1950 23488
rect 2006 23432 2011 23488
rect 1780 23430 2011 23432
rect 1780 23428 1786 23430
rect 1945 23427 2011 23430
rect 15653 23492 15719 23493
rect 15653 23488 15700 23492
rect 15764 23490 15770 23492
rect 15653 23432 15658 23488
rect 15653 23428 15700 23432
rect 15764 23430 15810 23490
rect 15764 23428 15770 23430
rect 15653 23427 15719 23428
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 200 22538 800 22568
rect 1761 22538 1827 22541
rect 200 22536 1827 22538
rect 200 22480 1766 22536
rect 1822 22480 1827 22536
rect 200 22478 1827 22480
rect 200 22448 800 22478
rect 1761 22475 1827 22478
rect 38193 22538 38259 22541
rect 39200 22538 39800 22568
rect 38193 22536 39800 22538
rect 38193 22480 38198 22536
rect 38254 22480 39800 22536
rect 38193 22478 39800 22480
rect 38193 22475 38259 22478
rect 39200 22448 39800 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 15377 21994 15443 21997
rect 15745 21994 15811 21997
rect 15377 21992 15811 21994
rect 15377 21936 15382 21992
rect 15438 21936 15750 21992
rect 15806 21936 15811 21992
rect 15377 21934 15811 21936
rect 15377 21931 15443 21934
rect 15745 21931 15811 21934
rect 15837 21858 15903 21861
rect 18597 21858 18663 21861
rect 15837 21856 18663 21858
rect 15837 21800 15842 21856
rect 15898 21800 18602 21856
rect 18658 21800 18663 21856
rect 15837 21798 18663 21800
rect 15837 21795 15903 21798
rect 18597 21795 18663 21798
rect 38193 21858 38259 21861
rect 39200 21858 39800 21888
rect 38193 21856 39800 21858
rect 38193 21800 38198 21856
rect 38254 21800 39800 21856
rect 38193 21798 39800 21800
rect 38193 21795 38259 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 39200 21768 39800 21798
rect 19570 21727 19886 21728
rect 13169 21314 13235 21317
rect 17953 21314 18019 21317
rect 13169 21312 18019 21314
rect 13169 21256 13174 21312
rect 13230 21256 17958 21312
rect 18014 21256 18019 21312
rect 13169 21254 18019 21256
rect 13169 21251 13235 21254
rect 17953 21251 18019 21254
rect 4210 21248 4526 21249
rect 200 21178 800 21208
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 1669 21178 1735 21181
rect 200 21176 1735 21178
rect 200 21120 1674 21176
rect 1730 21120 1735 21176
rect 200 21118 1735 21120
rect 200 21088 800 21118
rect 1669 21115 1735 21118
rect 14365 21178 14431 21181
rect 22001 21178 22067 21181
rect 14365 21176 22067 21178
rect 14365 21120 14370 21176
rect 14426 21120 22006 21176
rect 22062 21120 22067 21176
rect 14365 21118 22067 21120
rect 14365 21115 14431 21118
rect 22001 21115 22067 21118
rect 12985 21042 13051 21045
rect 16941 21042 17007 21045
rect 12985 21040 17007 21042
rect 12985 20984 12990 21040
rect 13046 20984 16946 21040
rect 17002 20984 17007 21040
rect 12985 20982 17007 20984
rect 12985 20979 13051 20982
rect 16941 20979 17007 20982
rect 17401 21042 17467 21045
rect 18597 21042 18663 21045
rect 17401 21040 18663 21042
rect 17401 20984 17406 21040
rect 17462 20984 18602 21040
rect 18658 20984 18663 21040
rect 17401 20982 18663 20984
rect 17401 20979 17467 20982
rect 18597 20979 18663 20982
rect 22737 21042 22803 21045
rect 23749 21042 23815 21045
rect 22737 21040 23815 21042
rect 22737 20984 22742 21040
rect 22798 20984 23754 21040
rect 23810 20984 23815 21040
rect 22737 20982 23815 20984
rect 22737 20979 22803 20982
rect 23749 20979 23815 20982
rect 4521 20770 4587 20773
rect 4838 20770 4844 20772
rect 4521 20768 4844 20770
rect 4521 20712 4526 20768
rect 4582 20712 4844 20768
rect 4521 20710 4844 20712
rect 4521 20707 4587 20710
rect 4838 20708 4844 20710
rect 4908 20708 4914 20772
rect 9581 20770 9647 20773
rect 13261 20770 13327 20773
rect 9581 20768 13327 20770
rect 9581 20712 9586 20768
rect 9642 20712 13266 20768
rect 13322 20712 13327 20768
rect 9581 20710 13327 20712
rect 9581 20707 9647 20710
rect 13261 20707 13327 20710
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 200 20498 800 20528
rect 1577 20498 1643 20501
rect 200 20496 1643 20498
rect 200 20440 1582 20496
rect 1638 20440 1643 20496
rect 200 20438 1643 20440
rect 200 20408 800 20438
rect 1577 20435 1643 20438
rect 38285 20498 38351 20501
rect 39200 20498 39800 20528
rect 38285 20496 39800 20498
rect 38285 20440 38290 20496
rect 38346 20440 39800 20496
rect 38285 20438 39800 20440
rect 38285 20435 38351 20438
rect 39200 20408 39800 20438
rect 14273 20362 14339 20365
rect 14406 20362 14412 20364
rect 14273 20360 14412 20362
rect 14273 20304 14278 20360
rect 14334 20304 14412 20360
rect 14273 20302 14412 20304
rect 14273 20299 14339 20302
rect 14406 20300 14412 20302
rect 14476 20300 14482 20364
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 10869 19412 10935 19413
rect 10869 19408 10916 19412
rect 10980 19410 10986 19412
rect 12617 19410 12683 19413
rect 15929 19410 15995 19413
rect 37273 19410 37339 19413
rect 10869 19352 10874 19408
rect 10869 19348 10916 19352
rect 10980 19350 11026 19410
rect 12617 19408 12818 19410
rect 12617 19352 12622 19408
rect 12678 19352 12818 19408
rect 12617 19350 12818 19352
rect 10980 19348 10986 19350
rect 10869 19347 10935 19348
rect 12617 19347 12683 19350
rect 12065 19274 12131 19277
rect 12617 19274 12683 19277
rect 12065 19272 12683 19274
rect 12065 19216 12070 19272
rect 12126 19216 12622 19272
rect 12678 19216 12683 19272
rect 12065 19214 12683 19216
rect 12065 19211 12131 19214
rect 12617 19211 12683 19214
rect 200 19138 800 19168
rect 1761 19138 1827 19141
rect 200 19136 1827 19138
rect 200 19080 1766 19136
rect 1822 19080 1827 19136
rect 200 19078 1827 19080
rect 12758 19138 12818 19350
rect 15929 19408 37339 19410
rect 15929 19352 15934 19408
rect 15990 19352 37278 19408
rect 37334 19352 37339 19408
rect 15929 19350 37339 19352
rect 15929 19347 15995 19350
rect 37273 19347 37339 19350
rect 12985 19138 13051 19141
rect 12758 19136 13051 19138
rect 12758 19080 12990 19136
rect 13046 19080 13051 19136
rect 12758 19078 13051 19080
rect 200 19048 800 19078
rect 1761 19075 1827 19078
rect 12985 19075 13051 19078
rect 38193 19138 38259 19141
rect 39200 19138 39800 19168
rect 38193 19136 39800 19138
rect 38193 19080 38198 19136
rect 38254 19080 39800 19136
rect 38193 19078 39800 19080
rect 38193 19075 38259 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 39200 19048 39800 19078
rect 34930 19007 35246 19008
rect 11237 19002 11303 19005
rect 16665 19002 16731 19005
rect 11237 19000 16731 19002
rect 11237 18944 11242 19000
rect 11298 18944 16670 19000
rect 16726 18944 16731 19000
rect 11237 18942 16731 18944
rect 11237 18939 11303 18942
rect 16665 18939 16731 18942
rect 11697 18730 11763 18733
rect 11830 18730 11836 18732
rect 11697 18728 11836 18730
rect 11697 18672 11702 18728
rect 11758 18672 11836 18728
rect 11697 18670 11836 18672
rect 11697 18667 11763 18670
rect 11830 18668 11836 18670
rect 11900 18668 11906 18732
rect 20110 18668 20116 18732
rect 20180 18730 20186 18732
rect 20253 18730 20319 18733
rect 20180 18728 20319 18730
rect 20180 18672 20258 18728
rect 20314 18672 20319 18728
rect 20180 18670 20319 18672
rect 20180 18668 20186 18670
rect 20253 18667 20319 18670
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 11329 18458 11395 18461
rect 11789 18458 11855 18461
rect 11329 18456 11530 18458
rect 11329 18400 11334 18456
rect 11390 18400 11530 18456
rect 11329 18398 11530 18400
rect 11329 18395 11395 18398
rect 11470 18186 11530 18398
rect 11789 18456 12450 18458
rect 11789 18400 11794 18456
rect 11850 18400 12450 18456
rect 11789 18398 12450 18400
rect 11789 18395 11855 18398
rect 12390 18322 12450 18398
rect 39200 18368 39800 18488
rect 15837 18322 15903 18325
rect 12390 18320 15903 18322
rect 12390 18264 15842 18320
rect 15898 18264 15903 18320
rect 12390 18262 15903 18264
rect 15837 18259 15903 18262
rect 11697 18186 11763 18189
rect 11470 18184 11763 18186
rect 11470 18128 11702 18184
rect 11758 18128 11763 18184
rect 11470 18126 11763 18128
rect 11697 18123 11763 18126
rect 21582 18124 21588 18188
rect 21652 18186 21658 18188
rect 28901 18186 28967 18189
rect 21652 18184 28967 18186
rect 21652 18128 28906 18184
rect 28962 18128 28967 18184
rect 21652 18126 28967 18128
rect 21652 18124 21658 18126
rect 28901 18123 28967 18126
rect 17350 17988 17356 18052
rect 17420 18050 17426 18052
rect 20529 18050 20595 18053
rect 17420 18048 20595 18050
rect 17420 17992 20534 18048
rect 20590 17992 20595 18048
rect 17420 17990 20595 17992
rect 17420 17988 17426 17990
rect 20529 17987 20595 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 200 17778 800 17808
rect 1577 17778 1643 17781
rect 200 17776 1643 17778
rect 200 17720 1582 17776
rect 1638 17720 1643 17776
rect 200 17718 1643 17720
rect 200 17688 800 17718
rect 1577 17715 1643 17718
rect 4245 17642 4311 17645
rect 8886 17642 8892 17644
rect 4245 17640 8892 17642
rect 4245 17584 4250 17640
rect 4306 17584 8892 17640
rect 4245 17582 8892 17584
rect 4245 17579 4311 17582
rect 8886 17580 8892 17582
rect 8956 17580 8962 17644
rect 11329 17642 11395 17645
rect 13670 17642 13676 17644
rect 11329 17640 13676 17642
rect 11329 17584 11334 17640
rect 11390 17584 13676 17640
rect 11329 17582 13676 17584
rect 11329 17579 11395 17582
rect 13670 17580 13676 17582
rect 13740 17642 13746 17644
rect 16113 17642 16179 17645
rect 13740 17640 16179 17642
rect 13740 17584 16118 17640
rect 16174 17584 16179 17640
rect 13740 17582 16179 17584
rect 13740 17580 13746 17582
rect 16113 17579 16179 17582
rect 19977 17642 20043 17645
rect 20294 17642 20300 17644
rect 19977 17640 20300 17642
rect 19977 17584 19982 17640
rect 20038 17584 20300 17640
rect 19977 17582 20300 17584
rect 19977 17579 20043 17582
rect 20294 17580 20300 17582
rect 20364 17580 20370 17644
rect 8477 17506 8543 17509
rect 14273 17506 14339 17509
rect 8477 17504 14339 17506
rect 8477 17448 8482 17504
rect 8538 17448 14278 17504
rect 14334 17448 14339 17504
rect 8477 17446 14339 17448
rect 8477 17443 8543 17446
rect 14273 17443 14339 17446
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 12341 17370 12407 17373
rect 13721 17370 13787 17373
rect 12341 17368 13787 17370
rect 12341 17312 12346 17368
rect 12402 17312 13726 17368
rect 13782 17312 13787 17368
rect 12341 17310 13787 17312
rect 12341 17307 12407 17310
rect 13721 17307 13787 17310
rect 9765 17234 9831 17237
rect 18413 17234 18479 17237
rect 9765 17232 18479 17234
rect 9765 17176 9770 17232
rect 9826 17176 18418 17232
rect 18474 17176 18479 17232
rect 9765 17174 18479 17176
rect 9765 17171 9831 17174
rect 200 17098 800 17128
rect 12252 17101 12312 17174
rect 18413 17171 18479 17174
rect 1761 17098 1827 17101
rect 200 17096 1827 17098
rect 200 17040 1766 17096
rect 1822 17040 1827 17096
rect 200 17038 1827 17040
rect 200 17008 800 17038
rect 1761 17035 1827 17038
rect 10225 17098 10291 17101
rect 10869 17098 10935 17101
rect 10225 17096 10935 17098
rect 10225 17040 10230 17096
rect 10286 17040 10874 17096
rect 10930 17040 10935 17096
rect 10225 17038 10935 17040
rect 10225 17035 10291 17038
rect 10869 17035 10935 17038
rect 12249 17096 12315 17101
rect 12249 17040 12254 17096
rect 12310 17040 12315 17096
rect 12249 17035 12315 17040
rect 17953 17098 18019 17101
rect 19374 17098 19380 17100
rect 17953 17096 19380 17098
rect 17953 17040 17958 17096
rect 18014 17040 19380 17096
rect 17953 17038 19380 17040
rect 17953 17035 18019 17038
rect 19374 17036 19380 17038
rect 19444 17036 19450 17100
rect 19609 17098 19675 17101
rect 20713 17098 20779 17101
rect 19609 17096 20779 17098
rect 19609 17040 19614 17096
rect 19670 17040 20718 17096
rect 20774 17040 20779 17096
rect 19609 17038 20779 17040
rect 19609 17035 19675 17038
rect 20713 17035 20779 17038
rect 38193 17098 38259 17101
rect 39200 17098 39800 17128
rect 38193 17096 39800 17098
rect 38193 17040 38198 17096
rect 38254 17040 39800 17096
rect 38193 17038 39800 17040
rect 38193 17035 38259 17038
rect 39200 17008 39800 17038
rect 9673 16962 9739 16965
rect 11605 16962 11671 16965
rect 9673 16960 11671 16962
rect 9673 16904 9678 16960
rect 9734 16904 11610 16960
rect 11666 16904 11671 16960
rect 9673 16902 11671 16904
rect 9673 16899 9739 16902
rect 11605 16899 11671 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 10593 16826 10659 16829
rect 11094 16826 11100 16828
rect 10593 16824 11100 16826
rect 10593 16768 10598 16824
rect 10654 16768 11100 16824
rect 10593 16766 11100 16768
rect 10593 16763 10659 16766
rect 11094 16764 11100 16766
rect 11164 16764 11170 16828
rect 7833 16690 7899 16693
rect 7966 16690 7972 16692
rect 7833 16688 7972 16690
rect 7833 16632 7838 16688
rect 7894 16632 7972 16688
rect 7833 16630 7972 16632
rect 7833 16627 7899 16630
rect 7966 16628 7972 16630
rect 8036 16628 8042 16692
rect 10869 16690 10935 16693
rect 13486 16690 13492 16692
rect 10869 16688 13492 16690
rect 10869 16632 10874 16688
rect 10930 16632 13492 16688
rect 10869 16630 13492 16632
rect 10869 16627 10935 16630
rect 13486 16628 13492 16630
rect 13556 16628 13562 16692
rect 19517 16690 19583 16693
rect 25814 16690 25820 16692
rect 19517 16688 25820 16690
rect 19517 16632 19522 16688
rect 19578 16632 25820 16688
rect 19517 16630 25820 16632
rect 19517 16627 19583 16630
rect 25814 16628 25820 16630
rect 25884 16628 25890 16692
rect 20805 16554 20871 16557
rect 23381 16554 23447 16557
rect 20805 16552 23447 16554
rect 20805 16496 20810 16552
rect 20866 16496 23386 16552
rect 23442 16496 23447 16552
rect 20805 16494 23447 16496
rect 20805 16491 20871 16494
rect 23381 16491 23447 16494
rect 8017 16418 8083 16421
rect 12566 16418 12572 16420
rect 8017 16416 12572 16418
rect 8017 16360 8022 16416
rect 8078 16360 12572 16416
rect 8017 16358 12572 16360
rect 8017 16355 8083 16358
rect 12566 16356 12572 16358
rect 12636 16356 12642 16420
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 14089 16146 14155 16149
rect 16573 16146 16639 16149
rect 22461 16146 22527 16149
rect 14089 16144 22527 16146
rect 14089 16088 14094 16144
rect 14150 16088 16578 16144
rect 16634 16088 22466 16144
rect 22522 16088 22527 16144
rect 14089 16086 22527 16088
rect 14089 16083 14155 16086
rect 16573 16083 16639 16086
rect 22461 16083 22527 16086
rect 13445 16012 13511 16013
rect 13445 16010 13492 16012
rect 13400 16008 13492 16010
rect 13400 15952 13450 16008
rect 13400 15950 13492 15952
rect 13445 15948 13492 15950
rect 13556 15948 13562 16012
rect 13445 15947 13511 15948
rect 4210 15808 4526 15809
rect 200 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 1761 15738 1827 15741
rect 200 15736 1827 15738
rect 200 15680 1766 15736
rect 1822 15680 1827 15736
rect 200 15678 1827 15680
rect 200 15648 800 15678
rect 1761 15675 1827 15678
rect 9765 15738 9831 15741
rect 18689 15738 18755 15741
rect 9765 15736 18755 15738
rect 9765 15680 9770 15736
rect 9826 15680 18694 15736
rect 18750 15680 18755 15736
rect 9765 15678 18755 15680
rect 9765 15675 9831 15678
rect 18689 15675 18755 15678
rect 38193 15738 38259 15741
rect 39200 15738 39800 15768
rect 38193 15736 39800 15738
rect 38193 15680 38198 15736
rect 38254 15680 39800 15736
rect 38193 15678 39800 15680
rect 38193 15675 38259 15678
rect 39200 15648 39800 15678
rect 8017 15602 8083 15605
rect 8293 15602 8359 15605
rect 8017 15600 8359 15602
rect 8017 15544 8022 15600
rect 8078 15544 8298 15600
rect 8354 15544 8359 15600
rect 8017 15542 8359 15544
rect 8017 15539 8083 15542
rect 8293 15539 8359 15542
rect 8477 15602 8543 15605
rect 9581 15602 9647 15605
rect 8477 15600 9647 15602
rect 8477 15544 8482 15600
rect 8538 15544 9586 15600
rect 9642 15544 9647 15600
rect 8477 15542 9647 15544
rect 8477 15539 8543 15542
rect 9581 15539 9647 15542
rect 11973 15602 12039 15605
rect 14089 15602 14155 15605
rect 11973 15600 14155 15602
rect 11973 15544 11978 15600
rect 12034 15544 14094 15600
rect 14150 15544 14155 15600
rect 11973 15542 14155 15544
rect 11973 15539 12039 15542
rect 14089 15539 14155 15542
rect 17125 15604 17191 15605
rect 17125 15600 17172 15604
rect 17236 15602 17242 15604
rect 19333 15602 19399 15605
rect 20478 15602 20484 15604
rect 17125 15544 17130 15600
rect 17125 15540 17172 15544
rect 17236 15542 17282 15602
rect 19333 15600 20484 15602
rect 19333 15544 19338 15600
rect 19394 15544 20484 15600
rect 19333 15542 20484 15544
rect 17236 15540 17242 15542
rect 17125 15539 17191 15540
rect 19333 15539 19399 15542
rect 20478 15540 20484 15542
rect 20548 15540 20554 15604
rect 7557 15466 7623 15469
rect 9765 15466 9831 15469
rect 7557 15464 9831 15466
rect 7557 15408 7562 15464
rect 7618 15408 9770 15464
rect 9826 15408 9831 15464
rect 7557 15406 9831 15408
rect 7557 15403 7623 15406
rect 9765 15403 9831 15406
rect 12341 15466 12407 15469
rect 12985 15466 13051 15469
rect 12341 15464 13051 15466
rect 12341 15408 12346 15464
rect 12402 15408 12990 15464
rect 13046 15408 13051 15464
rect 12341 15406 13051 15408
rect 12341 15403 12407 15406
rect 12985 15403 13051 15406
rect 13813 15466 13879 15469
rect 15377 15466 15443 15469
rect 17953 15466 18019 15469
rect 13813 15464 18019 15466
rect 13813 15408 13818 15464
rect 13874 15408 15382 15464
rect 15438 15408 17958 15464
rect 18014 15408 18019 15464
rect 13813 15406 18019 15408
rect 13813 15403 13879 15406
rect 15377 15403 15443 15406
rect 17953 15403 18019 15406
rect 19517 15466 19583 15469
rect 20529 15466 20595 15469
rect 19517 15464 20595 15466
rect 19517 15408 19522 15464
rect 19578 15408 20534 15464
rect 20590 15408 20595 15464
rect 19517 15406 20595 15408
rect 19517 15403 19583 15406
rect 20529 15403 20595 15406
rect 12801 15330 12867 15333
rect 13302 15330 13308 15332
rect 12801 15328 13308 15330
rect 12801 15272 12806 15328
rect 12862 15272 13308 15328
rect 12801 15270 13308 15272
rect 12801 15267 12867 15270
rect 13302 15268 13308 15270
rect 13372 15268 13378 15332
rect 14590 15268 14596 15332
rect 14660 15330 14666 15332
rect 14825 15330 14891 15333
rect 14660 15328 14891 15330
rect 14660 15272 14830 15328
rect 14886 15272 14891 15328
rect 14660 15270 14891 15272
rect 14660 15268 14666 15270
rect 14825 15267 14891 15270
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 13077 15194 13143 15197
rect 13537 15194 13603 15197
rect 13077 15192 13603 15194
rect 13077 15136 13082 15192
rect 13138 15136 13542 15192
rect 13598 15136 13603 15192
rect 13077 15134 13603 15136
rect 13077 15131 13143 15134
rect 13537 15131 13603 15134
rect 20621 15196 20687 15197
rect 20621 15192 20668 15196
rect 20732 15194 20738 15196
rect 20621 15136 20626 15192
rect 20621 15132 20668 15136
rect 20732 15134 20778 15194
rect 20732 15132 20738 15134
rect 20621 15131 20687 15132
rect 10961 15058 11027 15061
rect 12525 15058 12591 15061
rect 10961 15056 12591 15058
rect 10961 15000 10966 15056
rect 11022 15000 12530 15056
rect 12586 15000 12591 15056
rect 10961 14998 12591 15000
rect 10961 14995 11027 14998
rect 12525 14995 12591 14998
rect 19374 14996 19380 15060
rect 19444 15058 19450 15060
rect 20069 15058 20135 15061
rect 19444 15056 20135 15058
rect 19444 15000 20074 15056
rect 20130 15000 20135 15056
rect 19444 14998 20135 15000
rect 19444 14996 19450 14998
rect 20069 14995 20135 14998
rect 38101 15058 38167 15061
rect 39200 15058 39800 15088
rect 38101 15056 39800 15058
rect 38101 15000 38106 15056
rect 38162 15000 39800 15056
rect 38101 14998 39800 15000
rect 38101 14995 38167 14998
rect 39200 14968 39800 14998
rect 11881 14922 11947 14925
rect 13813 14922 13879 14925
rect 11881 14920 13879 14922
rect 11881 14864 11886 14920
rect 11942 14864 13818 14920
rect 13874 14864 13879 14920
rect 11881 14862 13879 14864
rect 11881 14859 11947 14862
rect 13813 14859 13879 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 19517 14650 19583 14653
rect 23197 14650 23263 14653
rect 19517 14648 23263 14650
rect 19517 14592 19522 14648
rect 19578 14592 23202 14648
rect 23258 14592 23263 14648
rect 19517 14590 23263 14592
rect 19517 14587 19583 14590
rect 23197 14587 23263 14590
rect 6085 14514 6151 14517
rect 8477 14514 8543 14517
rect 6085 14512 8543 14514
rect 6085 14456 6090 14512
rect 6146 14456 8482 14512
rect 8538 14456 8543 14512
rect 6085 14454 8543 14456
rect 6085 14451 6151 14454
rect 8477 14451 8543 14454
rect 9765 14514 9831 14517
rect 10961 14514 11027 14517
rect 20437 14514 20503 14517
rect 9765 14512 20503 14514
rect 9765 14456 9770 14512
rect 9826 14456 10966 14512
rect 11022 14456 20442 14512
rect 20498 14456 20503 14512
rect 9765 14454 20503 14456
rect 9765 14451 9831 14454
rect 10961 14451 11027 14454
rect 20437 14451 20503 14454
rect 200 14378 800 14408
rect 1761 14378 1827 14381
rect 200 14376 1827 14378
rect 200 14320 1766 14376
rect 1822 14320 1827 14376
rect 200 14318 1827 14320
rect 200 14288 800 14318
rect 1761 14315 1827 14318
rect 4705 14378 4771 14381
rect 7833 14378 7899 14381
rect 9121 14378 9187 14381
rect 16113 14380 16179 14381
rect 4705 14376 9187 14378
rect 4705 14320 4710 14376
rect 4766 14320 7838 14376
rect 7894 14320 9126 14376
rect 9182 14320 9187 14376
rect 4705 14318 9187 14320
rect 4705 14315 4771 14318
rect 7833 14315 7899 14318
rect 9121 14315 9187 14318
rect 16062 14316 16068 14380
rect 16132 14378 16179 14380
rect 16297 14378 16363 14381
rect 16132 14376 16363 14378
rect 16174 14320 16302 14376
rect 16358 14320 16363 14376
rect 16132 14318 16363 14320
rect 16132 14316 16179 14318
rect 16113 14315 16179 14316
rect 16297 14315 16363 14318
rect 18137 14242 18203 14245
rect 18638 14242 18644 14244
rect 18137 14240 18644 14242
rect 18137 14184 18142 14240
rect 18198 14184 18644 14240
rect 18137 14182 18644 14184
rect 18137 14179 18203 14182
rect 18638 14180 18644 14182
rect 18708 14180 18714 14244
rect 20294 14180 20300 14244
rect 20364 14242 20370 14244
rect 20437 14242 20503 14245
rect 20364 14240 20503 14242
rect 20364 14184 20442 14240
rect 20498 14184 20503 14240
rect 20364 14182 20503 14184
rect 20364 14180 20370 14182
rect 20437 14179 20503 14182
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 5073 13970 5139 13973
rect 6913 13970 6979 13973
rect 11513 13970 11579 13973
rect 11789 13970 11855 13973
rect 5073 13968 11855 13970
rect 5073 13912 5078 13968
rect 5134 13912 6918 13968
rect 6974 13912 11518 13968
rect 11574 13912 11794 13968
rect 11850 13912 11855 13968
rect 5073 13910 11855 13912
rect 5073 13907 5139 13910
rect 6913 13907 6979 13910
rect 11513 13907 11579 13910
rect 11789 13907 11855 13910
rect 12341 13970 12407 13973
rect 15009 13970 15075 13973
rect 12341 13968 15075 13970
rect 12341 13912 12346 13968
rect 12402 13912 15014 13968
rect 15070 13912 15075 13968
rect 12341 13910 15075 13912
rect 12341 13907 12407 13910
rect 15009 13907 15075 13910
rect 1894 13772 1900 13836
rect 1964 13834 1970 13836
rect 3693 13834 3759 13837
rect 1964 13832 3759 13834
rect 1964 13776 3698 13832
rect 3754 13776 3759 13832
rect 1964 13774 3759 13776
rect 1964 13772 1970 13774
rect 3693 13771 3759 13774
rect 11881 13834 11947 13837
rect 18229 13834 18295 13837
rect 11881 13832 18295 13834
rect 11881 13776 11886 13832
rect 11942 13776 18234 13832
rect 18290 13776 18295 13832
rect 11881 13774 18295 13776
rect 11881 13771 11947 13774
rect 18229 13771 18295 13774
rect 200 13698 800 13728
rect 1761 13698 1827 13701
rect 200 13696 1827 13698
rect 200 13640 1766 13696
rect 1822 13640 1827 13696
rect 200 13638 1827 13640
rect 200 13608 800 13638
rect 1761 13635 1827 13638
rect 12985 13698 13051 13701
rect 13629 13700 13695 13701
rect 13629 13698 13676 13700
rect 12985 13696 13676 13698
rect 12985 13640 12990 13696
rect 13046 13640 13634 13696
rect 12985 13638 13676 13640
rect 12985 13635 13051 13638
rect 13629 13636 13676 13638
rect 13740 13636 13746 13700
rect 38193 13698 38259 13701
rect 39200 13698 39800 13728
rect 38193 13696 39800 13698
rect 38193 13640 38198 13696
rect 38254 13640 39800 13696
rect 38193 13638 39800 13640
rect 13629 13635 13695 13636
rect 38193 13635 38259 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 39200 13608 39800 13638
rect 34930 13567 35246 13568
rect 6821 13562 6887 13565
rect 9121 13562 9187 13565
rect 6821 13560 9187 13562
rect 6821 13504 6826 13560
rect 6882 13504 9126 13560
rect 9182 13504 9187 13560
rect 6821 13502 9187 13504
rect 6821 13499 6887 13502
rect 9121 13499 9187 13502
rect 10910 13500 10916 13564
rect 10980 13562 10986 13564
rect 15653 13562 15719 13565
rect 10980 13560 15719 13562
rect 10980 13504 15658 13560
rect 15714 13504 15719 13560
rect 10980 13502 15719 13504
rect 10980 13500 10986 13502
rect 15653 13499 15719 13502
rect 6821 13426 6887 13429
rect 12525 13426 12591 13429
rect 6821 13424 12591 13426
rect 6821 13368 6826 13424
rect 6882 13368 12530 13424
rect 12586 13368 12591 13424
rect 6821 13366 12591 13368
rect 6821 13363 6887 13366
rect 12525 13363 12591 13366
rect 13486 13364 13492 13428
rect 13556 13426 13562 13428
rect 24393 13426 24459 13429
rect 13556 13424 24459 13426
rect 13556 13368 24398 13424
rect 24454 13368 24459 13424
rect 13556 13366 24459 13368
rect 13556 13364 13562 13366
rect 24393 13363 24459 13366
rect 19701 13290 19767 13293
rect 25589 13290 25655 13293
rect 19701 13288 25655 13290
rect 19701 13232 19706 13288
rect 19762 13232 25594 13288
rect 25650 13232 25655 13288
rect 19701 13230 25655 13232
rect 19701 13227 19767 13230
rect 25589 13227 25655 13230
rect 9121 13154 9187 13157
rect 9581 13154 9647 13157
rect 9121 13152 9647 13154
rect 9121 13096 9126 13152
rect 9182 13096 9586 13152
rect 9642 13096 9647 13152
rect 9121 13094 9647 13096
rect 9121 13091 9187 13094
rect 9581 13091 9647 13094
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 19977 13018 20043 13021
rect 20478 13018 20484 13020
rect 19977 13016 20484 13018
rect 19977 12960 19982 13016
rect 20038 12960 20484 13016
rect 19977 12958 20484 12960
rect 19977 12955 20043 12958
rect 20478 12956 20484 12958
rect 20548 12956 20554 13020
rect 4889 12882 4955 12885
rect 9673 12882 9739 12885
rect 10542 12882 10548 12884
rect 4889 12880 10548 12882
rect 4889 12824 4894 12880
rect 4950 12824 9678 12880
rect 9734 12824 10548 12880
rect 4889 12822 10548 12824
rect 4889 12819 4955 12822
rect 9673 12819 9739 12822
rect 10542 12820 10548 12822
rect 10612 12820 10618 12884
rect 22645 12882 22711 12885
rect 23105 12882 23171 12885
rect 22645 12880 23171 12882
rect 22645 12824 22650 12880
rect 22706 12824 23110 12880
rect 23166 12824 23171 12880
rect 22645 12822 23171 12824
rect 22645 12819 22711 12822
rect 23105 12819 23171 12822
rect 7373 12746 7439 12749
rect 10225 12746 10291 12749
rect 12801 12746 12867 12749
rect 16941 12746 17007 12749
rect 7373 12744 17007 12746
rect 7373 12688 7378 12744
rect 7434 12688 10230 12744
rect 10286 12688 12806 12744
rect 12862 12688 16946 12744
rect 17002 12688 17007 12744
rect 7373 12686 17007 12688
rect 7373 12683 7439 12686
rect 10225 12683 10291 12686
rect 12801 12683 12867 12686
rect 16941 12683 17007 12686
rect 26877 12746 26943 12749
rect 27245 12746 27311 12749
rect 37365 12746 37431 12749
rect 26877 12744 37431 12746
rect 26877 12688 26882 12744
rect 26938 12688 27250 12744
rect 27306 12688 37370 12744
rect 37426 12688 37431 12744
rect 26877 12686 37431 12688
rect 26877 12683 26943 12686
rect 27245 12683 27311 12686
rect 37365 12683 37431 12686
rect 5533 12610 5599 12613
rect 6177 12610 6243 12613
rect 10685 12610 10751 12613
rect 11421 12610 11487 12613
rect 5533 12608 11487 12610
rect 5533 12552 5538 12608
rect 5594 12552 6182 12608
rect 6238 12552 10690 12608
rect 10746 12552 11426 12608
rect 11482 12552 11487 12608
rect 5533 12550 11487 12552
rect 5533 12547 5599 12550
rect 6177 12547 6243 12550
rect 10685 12547 10751 12550
rect 11421 12547 11487 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 7557 12474 7623 12477
rect 8109 12474 8175 12477
rect 7557 12472 8175 12474
rect 7557 12416 7562 12472
rect 7618 12416 8114 12472
rect 8170 12416 8175 12472
rect 7557 12414 8175 12416
rect 7557 12411 7623 12414
rect 8109 12411 8175 12414
rect 9765 12474 9831 12477
rect 13169 12474 13235 12477
rect 18873 12474 18939 12477
rect 9765 12472 18939 12474
rect 9765 12416 9770 12472
rect 9826 12416 13174 12472
rect 13230 12416 18878 12472
rect 18934 12416 18939 12472
rect 9765 12414 18939 12416
rect 9765 12411 9831 12414
rect 13169 12411 13235 12414
rect 18873 12411 18939 12414
rect 21541 12474 21607 12477
rect 23473 12474 23539 12477
rect 21541 12472 23539 12474
rect 21541 12416 21546 12472
rect 21602 12416 23478 12472
rect 23534 12416 23539 12472
rect 21541 12414 23539 12416
rect 21541 12411 21607 12414
rect 23473 12411 23539 12414
rect 200 12338 800 12368
rect 1761 12338 1827 12341
rect 200 12336 1827 12338
rect 200 12280 1766 12336
rect 1822 12280 1827 12336
rect 200 12278 1827 12280
rect 200 12248 800 12278
rect 1761 12275 1827 12278
rect 10409 12338 10475 12341
rect 11421 12338 11487 12341
rect 10409 12336 11487 12338
rect 10409 12280 10414 12336
rect 10470 12280 11426 12336
rect 11482 12280 11487 12336
rect 10409 12278 11487 12280
rect 10409 12275 10475 12278
rect 11421 12275 11487 12278
rect 20621 12338 20687 12341
rect 28349 12338 28415 12341
rect 20621 12336 28415 12338
rect 20621 12280 20626 12336
rect 20682 12280 28354 12336
rect 28410 12280 28415 12336
rect 20621 12278 28415 12280
rect 20621 12275 20687 12278
rect 28349 12275 28415 12278
rect 38193 12338 38259 12341
rect 39200 12338 39800 12368
rect 38193 12336 39800 12338
rect 38193 12280 38198 12336
rect 38254 12280 39800 12336
rect 38193 12278 39800 12280
rect 38193 12275 38259 12278
rect 39200 12248 39800 12278
rect 9673 12202 9739 12205
rect 12525 12202 12591 12205
rect 9673 12200 12591 12202
rect 9673 12144 9678 12200
rect 9734 12144 12530 12200
rect 12586 12144 12591 12200
rect 9673 12142 12591 12144
rect 9673 12139 9739 12142
rect 12525 12139 12591 12142
rect 18638 12140 18644 12204
rect 18708 12202 18714 12204
rect 22093 12202 22159 12205
rect 18708 12200 22159 12202
rect 18708 12144 22098 12200
rect 22154 12144 22159 12200
rect 18708 12142 22159 12144
rect 18708 12140 18714 12142
rect 22093 12139 22159 12142
rect 23013 12202 23079 12205
rect 23289 12202 23355 12205
rect 23013 12200 23355 12202
rect 23013 12144 23018 12200
rect 23074 12144 23294 12200
rect 23350 12144 23355 12200
rect 23013 12142 23355 12144
rect 23013 12139 23079 12142
rect 23289 12139 23355 12142
rect 15561 12066 15627 12069
rect 18597 12066 18663 12069
rect 15561 12064 18663 12066
rect 15561 12008 15566 12064
rect 15622 12008 18602 12064
rect 18658 12008 18663 12064
rect 15561 12006 18663 12008
rect 15561 12003 15627 12006
rect 18597 12003 18663 12006
rect 23381 12066 23447 12069
rect 23974 12066 23980 12068
rect 23381 12064 23980 12066
rect 23381 12008 23386 12064
rect 23442 12008 23980 12064
rect 23381 12006 23980 12008
rect 23381 12003 23447 12006
rect 23974 12004 23980 12006
rect 24044 12066 24050 12068
rect 24485 12066 24551 12069
rect 24044 12064 24551 12066
rect 24044 12008 24490 12064
rect 24546 12008 24551 12064
rect 24044 12006 24551 12008
rect 24044 12004 24050 12006
rect 24485 12003 24551 12006
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 11513 11930 11579 11933
rect 11513 11928 12450 11930
rect 11513 11872 11518 11928
rect 11574 11872 12450 11928
rect 11513 11870 12450 11872
rect 11513 11867 11579 11870
rect 9489 11794 9555 11797
rect 11789 11794 11855 11797
rect 9489 11792 11855 11794
rect 9489 11736 9494 11792
rect 9550 11736 11794 11792
rect 11850 11736 11855 11792
rect 9489 11734 11855 11736
rect 12390 11794 12450 11870
rect 13445 11794 13511 11797
rect 12390 11792 13511 11794
rect 12390 11736 13450 11792
rect 13506 11736 13511 11792
rect 12390 11734 13511 11736
rect 9489 11731 9555 11734
rect 11789 11731 11855 11734
rect 13445 11731 13511 11734
rect 9857 11658 9923 11661
rect 12433 11658 12499 11661
rect 24209 11660 24275 11661
rect 9857 11656 12499 11658
rect 9857 11600 9862 11656
rect 9918 11600 12438 11656
rect 12494 11600 12499 11656
rect 9857 11598 12499 11600
rect 9857 11595 9923 11598
rect 12433 11595 12499 11598
rect 24158 11596 24164 11660
rect 24228 11658 24275 11660
rect 24228 11656 24320 11658
rect 24270 11600 24320 11656
rect 24228 11598 24320 11600
rect 24228 11596 24275 11598
rect 24209 11595 24275 11596
rect 12893 11522 12959 11525
rect 12574 11520 12959 11522
rect 12574 11464 12898 11520
rect 12954 11464 12959 11520
rect 12574 11462 12959 11464
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 6453 11250 6519 11253
rect 8569 11250 8635 11253
rect 6453 11248 8635 11250
rect 6453 11192 6458 11248
rect 6514 11192 8574 11248
rect 8630 11192 8635 11248
rect 6453 11190 8635 11192
rect 6453 11187 6519 11190
rect 8569 11187 8635 11190
rect 200 10978 800 11008
rect 1761 10978 1827 10981
rect 200 10976 1827 10978
rect 200 10920 1766 10976
rect 1822 10920 1827 10976
rect 200 10918 1827 10920
rect 200 10888 800 10918
rect 1761 10915 1827 10918
rect 12433 10978 12499 10981
rect 12574 10978 12634 11462
rect 12893 11459 12959 11462
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 14089 11250 14155 11253
rect 15285 11250 15351 11253
rect 14089 11248 15351 11250
rect 14089 11192 14094 11248
rect 14150 11192 15290 11248
rect 15346 11192 15351 11248
rect 14089 11190 15351 11192
rect 14089 11187 14155 11190
rect 15285 11187 15351 11190
rect 12433 10976 12634 10978
rect 12433 10920 12438 10976
rect 12494 10920 12634 10976
rect 12433 10918 12634 10920
rect 38193 10978 38259 10981
rect 39200 10978 39800 11008
rect 38193 10976 39800 10978
rect 38193 10920 38198 10976
rect 38254 10920 39800 10976
rect 38193 10918 39800 10920
rect 12433 10915 12499 10918
rect 38193 10915 38259 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 39200 10888 39800 10918
rect 19570 10847 19886 10848
rect 10777 10842 10843 10845
rect 16297 10842 16363 10845
rect 10777 10840 16363 10842
rect 10777 10784 10782 10840
rect 10838 10784 16302 10840
rect 16358 10784 16363 10840
rect 10777 10782 16363 10784
rect 10777 10779 10843 10782
rect 16297 10779 16363 10782
rect 4210 10368 4526 10369
rect 200 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 1761 10298 1827 10301
rect 200 10296 1827 10298
rect 200 10240 1766 10296
rect 1822 10240 1827 10296
rect 200 10238 1827 10240
rect 200 10208 800 10238
rect 1761 10235 1827 10238
rect 12566 10236 12572 10300
rect 12636 10298 12642 10300
rect 26969 10298 27035 10301
rect 12636 10296 27035 10298
rect 12636 10240 26974 10296
rect 27030 10240 27035 10296
rect 12636 10238 27035 10240
rect 12636 10236 12642 10238
rect 26969 10235 27035 10238
rect 38193 10298 38259 10301
rect 39200 10298 39800 10328
rect 38193 10296 39800 10298
rect 38193 10240 38198 10296
rect 38254 10240 39800 10296
rect 38193 10238 39800 10240
rect 38193 10235 38259 10238
rect 39200 10208 39800 10238
rect 17861 10162 17927 10165
rect 18454 10162 18460 10164
rect 17861 10160 18460 10162
rect 17861 10104 17866 10160
rect 17922 10104 18460 10160
rect 17861 10102 18460 10104
rect 17861 10099 17927 10102
rect 18454 10100 18460 10102
rect 18524 10100 18530 10164
rect 20662 10100 20668 10164
rect 20732 10162 20738 10164
rect 24669 10162 24735 10165
rect 20732 10160 24735 10162
rect 20732 10104 24674 10160
rect 24730 10104 24735 10160
rect 20732 10102 24735 10104
rect 20732 10100 20738 10102
rect 24669 10099 24735 10102
rect 9949 10026 10015 10029
rect 10593 10026 10659 10029
rect 9949 10024 10659 10026
rect 9949 9968 9954 10024
rect 10010 9968 10598 10024
rect 10654 9968 10659 10024
rect 9949 9966 10659 9968
rect 9949 9963 10015 9966
rect 10593 9963 10659 9966
rect 9765 9890 9831 9893
rect 10225 9890 10291 9893
rect 9765 9888 10291 9890
rect 9765 9832 9770 9888
rect 9826 9832 10230 9888
rect 10286 9832 10291 9888
rect 9765 9830 10291 9832
rect 9765 9827 9831 9830
rect 10225 9827 10291 9830
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 3785 9754 3851 9757
rect 4797 9754 4863 9757
rect 3785 9752 4863 9754
rect 3785 9696 3790 9752
rect 3846 9696 4802 9752
rect 4858 9696 4863 9752
rect 3785 9694 4863 9696
rect 3785 9691 3851 9694
rect 4797 9691 4863 9694
rect 6545 9754 6611 9757
rect 9581 9754 9647 9757
rect 6545 9752 9647 9754
rect 6545 9696 6550 9752
rect 6606 9696 9586 9752
rect 9642 9696 9647 9752
rect 6545 9694 9647 9696
rect 6545 9691 6611 9694
rect 9581 9691 9647 9694
rect 4521 9618 4587 9621
rect 9765 9618 9831 9621
rect 4521 9616 9831 9618
rect 4521 9560 4526 9616
rect 4582 9560 9770 9616
rect 9826 9560 9831 9616
rect 4521 9558 9831 9560
rect 4521 9555 4587 9558
rect 9765 9555 9831 9558
rect 10409 9618 10475 9621
rect 13077 9618 13143 9621
rect 10409 9616 13143 9618
rect 10409 9560 10414 9616
rect 10470 9560 13082 9616
rect 13138 9560 13143 9616
rect 10409 9558 13143 9560
rect 10409 9555 10475 9558
rect 13077 9555 13143 9558
rect 14590 9556 14596 9620
rect 14660 9618 14666 9620
rect 18781 9618 18847 9621
rect 14660 9616 18847 9618
rect 14660 9560 18786 9616
rect 18842 9560 18847 9616
rect 14660 9558 18847 9560
rect 14660 9556 14666 9558
rect 18781 9555 18847 9558
rect 3325 9482 3391 9485
rect 13537 9482 13603 9485
rect 24025 9484 24091 9485
rect 3325 9480 13603 9482
rect 3325 9424 3330 9480
rect 3386 9424 13542 9480
rect 13598 9424 13603 9480
rect 3325 9422 13603 9424
rect 3325 9419 3391 9422
rect 13537 9419 13603 9422
rect 23974 9420 23980 9484
rect 24044 9482 24091 9484
rect 24044 9480 24136 9482
rect 24086 9424 24136 9480
rect 24044 9422 24136 9424
rect 24044 9420 24091 9422
rect 24025 9419 24091 9420
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 7925 9210 7991 9213
rect 8385 9210 8451 9213
rect 7925 9208 8451 9210
rect 7925 9152 7930 9208
rect 7986 9152 8390 9208
rect 8446 9152 8451 9208
rect 7925 9150 8451 9152
rect 7925 9147 7991 9150
rect 8385 9147 8451 9150
rect 4061 9074 4127 9077
rect 9489 9074 9555 9077
rect 4061 9072 9555 9074
rect 4061 9016 4066 9072
rect 4122 9016 9494 9072
rect 9550 9016 9555 9072
rect 4061 9014 9555 9016
rect 4061 9011 4127 9014
rect 9489 9011 9555 9014
rect 12249 9074 12315 9077
rect 16297 9074 16363 9077
rect 16573 9074 16639 9077
rect 12249 9072 19350 9074
rect 12249 9016 12254 9072
rect 12310 9016 16302 9072
rect 16358 9016 16578 9072
rect 16634 9016 19350 9072
rect 12249 9014 19350 9016
rect 12249 9011 12315 9014
rect 16297 9011 16363 9014
rect 16573 9011 16639 9014
rect 200 8938 800 8968
rect 1761 8938 1827 8941
rect 200 8936 1827 8938
rect 200 8880 1766 8936
rect 1822 8880 1827 8936
rect 200 8878 1827 8880
rect 200 8848 800 8878
rect 1761 8875 1827 8878
rect 9581 8938 9647 8941
rect 14590 8938 14596 8940
rect 9581 8936 14596 8938
rect 9581 8880 9586 8936
rect 9642 8880 14596 8936
rect 9581 8878 14596 8880
rect 9581 8875 9647 8878
rect 14590 8876 14596 8878
rect 14660 8876 14666 8940
rect 19290 8938 19350 9014
rect 20713 8938 20779 8941
rect 19290 8936 20779 8938
rect 19290 8880 20718 8936
rect 20774 8880 20779 8936
rect 19290 8878 20779 8880
rect 20713 8875 20779 8878
rect 38285 8938 38351 8941
rect 39200 8938 39800 8968
rect 38285 8936 39800 8938
rect 38285 8880 38290 8936
rect 38346 8880 39800 8936
rect 38285 8878 39800 8880
rect 38285 8875 38351 8878
rect 39200 8848 39800 8878
rect 12433 8802 12499 8805
rect 15745 8802 15811 8805
rect 12433 8800 15811 8802
rect 12433 8744 12438 8800
rect 12494 8744 15750 8800
rect 15806 8744 15811 8800
rect 12433 8742 15811 8744
rect 12433 8739 12499 8742
rect 15745 8739 15811 8742
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 8845 8668 8911 8669
rect 8845 8666 8892 8668
rect 8800 8664 8892 8666
rect 8956 8666 8962 8668
rect 15101 8666 15167 8669
rect 17350 8666 17356 8668
rect 8956 8664 17356 8666
rect 8800 8608 8850 8664
rect 8956 8608 15106 8664
rect 15162 8608 17356 8664
rect 8800 8606 8892 8608
rect 8845 8604 8892 8606
rect 8956 8606 17356 8608
rect 8956 8604 8962 8606
rect 8845 8603 8911 8604
rect 15101 8603 15167 8606
rect 17350 8604 17356 8606
rect 17420 8604 17426 8668
rect 12341 8530 12407 8533
rect 13629 8530 13695 8533
rect 12341 8528 13695 8530
rect 12341 8472 12346 8528
rect 12402 8472 13634 8528
rect 13690 8472 13695 8528
rect 12341 8470 13695 8472
rect 12341 8467 12407 8470
rect 13629 8467 13695 8470
rect 1577 8394 1643 8397
rect 28625 8394 28691 8397
rect 1577 8392 28691 8394
rect 1577 8336 1582 8392
rect 1638 8336 28630 8392
rect 28686 8336 28691 8392
rect 1577 8334 28691 8336
rect 1577 8331 1643 8334
rect 28625 8331 28691 8334
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 4061 7986 4127 7989
rect 4838 7986 4844 7988
rect 4061 7984 4844 7986
rect 4061 7928 4066 7984
rect 4122 7928 4844 7984
rect 4061 7926 4844 7928
rect 4061 7923 4127 7926
rect 4838 7924 4844 7926
rect 4908 7924 4914 7988
rect 22369 7986 22435 7989
rect 23749 7986 23815 7989
rect 22369 7984 23815 7986
rect 22369 7928 22374 7984
rect 22430 7928 23754 7984
rect 23810 7928 23815 7984
rect 22369 7926 23815 7928
rect 22369 7923 22435 7926
rect 23749 7923 23815 7926
rect 4521 7714 4587 7717
rect 8293 7714 8359 7717
rect 4521 7712 8359 7714
rect 4521 7656 4526 7712
rect 4582 7656 8298 7712
rect 8354 7656 8359 7712
rect 4521 7654 8359 7656
rect 4521 7651 4587 7654
rect 8293 7651 8359 7654
rect 19570 7648 19886 7649
rect 200 7578 800 7608
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 1761 7578 1827 7581
rect 200 7576 1827 7578
rect 200 7520 1766 7576
rect 1822 7520 1827 7576
rect 200 7518 1827 7520
rect 200 7488 800 7518
rect 1761 7515 1827 7518
rect 5349 7578 5415 7581
rect 10225 7578 10291 7581
rect 5349 7576 10291 7578
rect 5349 7520 5354 7576
rect 5410 7520 10230 7576
rect 10286 7520 10291 7576
rect 5349 7518 10291 7520
rect 5349 7515 5415 7518
rect 10225 7515 10291 7518
rect 37457 7578 37523 7581
rect 39200 7578 39800 7608
rect 37457 7576 39800 7578
rect 37457 7520 37462 7576
rect 37518 7520 39800 7576
rect 37457 7518 39800 7520
rect 37457 7515 37523 7518
rect 39200 7488 39800 7518
rect 3693 7442 3759 7445
rect 7833 7442 7899 7445
rect 3693 7440 7899 7442
rect 3693 7384 3698 7440
rect 3754 7384 7838 7440
rect 7894 7384 7899 7440
rect 3693 7382 7899 7384
rect 3693 7379 3759 7382
rect 7833 7379 7899 7382
rect 15653 7442 15719 7445
rect 19977 7442 20043 7445
rect 15653 7440 20043 7442
rect 15653 7384 15658 7440
rect 15714 7384 19982 7440
rect 20038 7384 20043 7440
rect 15653 7382 20043 7384
rect 15653 7379 15719 7382
rect 19977 7379 20043 7382
rect 5073 7306 5139 7309
rect 9397 7306 9463 7309
rect 5073 7304 9463 7306
rect 5073 7248 5078 7304
rect 5134 7248 9402 7304
rect 9458 7248 9463 7304
rect 5073 7246 9463 7248
rect 5073 7243 5139 7246
rect 9397 7243 9463 7246
rect 13302 7244 13308 7308
rect 13372 7306 13378 7308
rect 19609 7306 19675 7309
rect 21081 7306 21147 7309
rect 13372 7246 16682 7306
rect 13372 7244 13378 7246
rect 12157 7170 12223 7173
rect 16389 7170 16455 7173
rect 12157 7168 16455 7170
rect 12157 7112 12162 7168
rect 12218 7112 16394 7168
rect 16450 7112 16455 7168
rect 12157 7110 16455 7112
rect 16622 7170 16682 7246
rect 19609 7304 21147 7306
rect 19609 7248 19614 7304
rect 19670 7248 21086 7304
rect 21142 7248 21147 7304
rect 19609 7246 21147 7248
rect 19609 7243 19675 7246
rect 21081 7243 21147 7246
rect 24209 7170 24275 7173
rect 24853 7170 24919 7173
rect 16622 7168 24919 7170
rect 16622 7112 24214 7168
rect 24270 7112 24858 7168
rect 24914 7112 24919 7168
rect 16622 7110 24919 7112
rect 12157 7107 12223 7110
rect 16389 7107 16455 7110
rect 24209 7107 24275 7110
rect 24853 7107 24919 7110
rect 26233 7170 26299 7173
rect 27981 7170 28047 7173
rect 26233 7168 28047 7170
rect 26233 7112 26238 7168
rect 26294 7112 27986 7168
rect 28042 7112 28047 7168
rect 26233 7110 28047 7112
rect 26233 7107 26299 7110
rect 27981 7107 28047 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 11881 7034 11947 7037
rect 17401 7034 17467 7037
rect 11881 7032 17467 7034
rect 11881 6976 11886 7032
rect 11942 6976 17406 7032
rect 17462 6976 17467 7032
rect 11881 6974 17467 6976
rect 11881 6971 11947 6974
rect 17401 6971 17467 6974
rect 200 6898 800 6928
rect 1393 6898 1459 6901
rect 200 6896 1459 6898
rect 200 6840 1398 6896
rect 1454 6840 1459 6896
rect 200 6838 1459 6840
rect 200 6808 800 6838
rect 1393 6835 1459 6838
rect 4337 6898 4403 6901
rect 7557 6898 7623 6901
rect 4337 6896 7623 6898
rect 4337 6840 4342 6896
rect 4398 6840 7562 6896
rect 7618 6840 7623 6896
rect 4337 6838 7623 6840
rect 4337 6835 4403 6838
rect 7557 6835 7623 6838
rect 11145 6898 11211 6901
rect 12157 6898 12223 6901
rect 11145 6896 12223 6898
rect 11145 6840 11150 6896
rect 11206 6840 12162 6896
rect 12218 6840 12223 6896
rect 11145 6838 12223 6840
rect 11145 6835 11211 6838
rect 12157 6835 12223 6838
rect 38285 6898 38351 6901
rect 39200 6898 39800 6928
rect 38285 6896 39800 6898
rect 38285 6840 38290 6896
rect 38346 6840 39800 6896
rect 38285 6838 39800 6840
rect 38285 6835 38351 6838
rect 39200 6808 39800 6838
rect 1669 6762 1735 6765
rect 8385 6762 8451 6765
rect 1669 6760 8451 6762
rect 1669 6704 1674 6760
rect 1730 6704 8390 6760
rect 8446 6704 8451 6760
rect 1669 6702 8451 6704
rect 1669 6699 1735 6702
rect 8385 6699 8451 6702
rect 12065 6762 12131 6765
rect 14365 6762 14431 6765
rect 12065 6760 14431 6762
rect 12065 6704 12070 6760
rect 12126 6704 14370 6760
rect 14426 6704 14431 6760
rect 12065 6702 14431 6704
rect 12065 6699 12131 6702
rect 14365 6699 14431 6702
rect 19609 6762 19675 6765
rect 20805 6762 20871 6765
rect 21173 6762 21239 6765
rect 19609 6760 21239 6762
rect 19609 6704 19614 6760
rect 19670 6704 20810 6760
rect 20866 6704 21178 6760
rect 21234 6704 21239 6760
rect 19609 6702 21239 6704
rect 19609 6699 19675 6702
rect 20805 6699 20871 6702
rect 21173 6699 21239 6702
rect 21541 6762 21607 6765
rect 26601 6762 26667 6765
rect 21541 6760 26667 6762
rect 21541 6704 21546 6760
rect 21602 6704 26606 6760
rect 26662 6704 26667 6760
rect 21541 6702 26667 6704
rect 21541 6699 21607 6702
rect 26601 6699 26667 6702
rect 5073 6626 5139 6629
rect 8661 6626 8727 6629
rect 5073 6624 8727 6626
rect 5073 6568 5078 6624
rect 5134 6568 8666 6624
rect 8722 6568 8727 6624
rect 5073 6566 8727 6568
rect 5073 6563 5139 6566
rect 8661 6563 8727 6566
rect 22001 6626 22067 6629
rect 23473 6626 23539 6629
rect 22001 6624 23539 6626
rect 22001 6568 22006 6624
rect 22062 6568 23478 6624
rect 23534 6568 23539 6624
rect 22001 6566 23539 6568
rect 22001 6563 22067 6566
rect 23473 6563 23539 6566
rect 24945 6626 25011 6629
rect 26325 6626 26391 6629
rect 24945 6624 26391 6626
rect 24945 6568 24950 6624
rect 25006 6568 26330 6624
rect 26386 6568 26391 6624
rect 24945 6566 26391 6568
rect 24945 6563 25011 6566
rect 26325 6563 26391 6566
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 8385 6490 8451 6493
rect 10317 6490 10383 6493
rect 8385 6488 10383 6490
rect 8385 6432 8390 6488
rect 8446 6432 10322 6488
rect 10378 6432 10383 6488
rect 8385 6430 10383 6432
rect 8385 6427 8451 6430
rect 10317 6427 10383 6430
rect 21817 6490 21883 6493
rect 23289 6490 23355 6493
rect 26785 6490 26851 6493
rect 21817 6488 26851 6490
rect 21817 6432 21822 6488
rect 21878 6432 23294 6488
rect 23350 6432 26790 6488
rect 26846 6432 26851 6488
rect 21817 6430 26851 6432
rect 21817 6427 21883 6430
rect 23289 6427 23355 6430
rect 26785 6427 26851 6430
rect 4061 6354 4127 6357
rect 18638 6354 18644 6356
rect 4061 6352 18644 6354
rect 4061 6296 4066 6352
rect 4122 6296 18644 6352
rect 4061 6294 18644 6296
rect 4061 6291 4127 6294
rect 18638 6292 18644 6294
rect 18708 6292 18714 6356
rect 19701 6354 19767 6357
rect 21265 6354 21331 6357
rect 19701 6352 21331 6354
rect 19701 6296 19706 6352
rect 19762 6296 21270 6352
rect 21326 6296 21331 6352
rect 19701 6294 21331 6296
rect 19701 6291 19767 6294
rect 21265 6291 21331 6294
rect 27153 6354 27219 6357
rect 27613 6354 27679 6357
rect 27153 6352 27679 6354
rect 27153 6296 27158 6352
rect 27214 6296 27618 6352
rect 27674 6296 27679 6352
rect 27153 6294 27679 6296
rect 27153 6291 27219 6294
rect 27613 6291 27679 6294
rect 7966 6156 7972 6220
rect 8036 6218 8042 6220
rect 8661 6218 8727 6221
rect 9581 6218 9647 6221
rect 8036 6216 9647 6218
rect 8036 6160 8666 6216
rect 8722 6160 9586 6216
rect 9642 6160 9647 6216
rect 8036 6158 9647 6160
rect 8036 6156 8042 6158
rect 8661 6155 8727 6158
rect 9581 6155 9647 6158
rect 10225 6218 10291 6221
rect 29729 6218 29795 6221
rect 10225 6216 29795 6218
rect 10225 6160 10230 6216
rect 10286 6160 29734 6216
rect 29790 6160 29795 6216
rect 10225 6158 29795 6160
rect 10225 6155 10291 6158
rect 29729 6155 29795 6158
rect 6637 6082 6703 6085
rect 9949 6082 10015 6085
rect 6637 6080 10015 6082
rect 6637 6024 6642 6080
rect 6698 6024 9954 6080
rect 10010 6024 10015 6080
rect 6637 6022 10015 6024
rect 6637 6019 6703 6022
rect 9949 6019 10015 6022
rect 11329 6082 11395 6085
rect 18413 6082 18479 6085
rect 11329 6080 18479 6082
rect 11329 6024 11334 6080
rect 11390 6024 18418 6080
rect 18474 6024 18479 6080
rect 11329 6022 18479 6024
rect 11329 6019 11395 6022
rect 18413 6019 18479 6022
rect 21173 6082 21239 6085
rect 29637 6082 29703 6085
rect 21173 6080 29703 6082
rect 21173 6024 21178 6080
rect 21234 6024 29642 6080
rect 29698 6024 29703 6080
rect 21173 6022 29703 6024
rect 21173 6019 21239 6022
rect 29637 6019 29703 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 6269 5946 6335 5949
rect 12249 5946 12315 5949
rect 28533 5946 28599 5949
rect 6269 5944 12315 5946
rect 6269 5888 6274 5944
rect 6330 5888 12254 5944
rect 12310 5888 12315 5944
rect 6269 5886 12315 5888
rect 6269 5883 6335 5886
rect 12249 5883 12315 5886
rect 22050 5944 28599 5946
rect 22050 5888 28538 5944
rect 28594 5888 28599 5944
rect 22050 5886 28599 5888
rect 22050 5813 22110 5886
rect 28533 5883 28599 5886
rect 6913 5810 6979 5813
rect 7925 5810 7991 5813
rect 6913 5808 7991 5810
rect 6913 5752 6918 5808
rect 6974 5752 7930 5808
rect 7986 5752 7991 5808
rect 6913 5750 7991 5752
rect 6913 5747 6979 5750
rect 7925 5747 7991 5750
rect 8477 5810 8543 5813
rect 14406 5810 14412 5812
rect 8477 5808 14412 5810
rect 8477 5752 8482 5808
rect 8538 5752 14412 5808
rect 8477 5750 14412 5752
rect 8477 5747 8543 5750
rect 14406 5748 14412 5750
rect 14476 5810 14482 5812
rect 14641 5810 14707 5813
rect 14476 5808 14707 5810
rect 14476 5752 14646 5808
rect 14702 5752 14707 5808
rect 14476 5750 14707 5752
rect 14476 5748 14482 5750
rect 14641 5747 14707 5750
rect 22001 5808 22110 5813
rect 22001 5752 22006 5808
rect 22062 5752 22110 5808
rect 22001 5750 22110 5752
rect 22737 5810 22803 5813
rect 29913 5810 29979 5813
rect 22737 5808 29979 5810
rect 22737 5752 22742 5808
rect 22798 5752 29918 5808
rect 29974 5752 29979 5808
rect 22737 5750 29979 5752
rect 22001 5747 22067 5750
rect 22737 5747 22803 5750
rect 29913 5747 29979 5750
rect 6545 5674 6611 5677
rect 11145 5674 11211 5677
rect 6545 5672 11211 5674
rect 6545 5616 6550 5672
rect 6606 5616 11150 5672
rect 11206 5616 11211 5672
rect 6545 5614 11211 5616
rect 6545 5611 6611 5614
rect 11145 5611 11211 5614
rect 12341 5674 12407 5677
rect 18229 5674 18295 5677
rect 21541 5676 21607 5677
rect 21541 5674 21588 5676
rect 12341 5672 18295 5674
rect 12341 5616 12346 5672
rect 12402 5616 18234 5672
rect 18290 5616 18295 5672
rect 12341 5614 18295 5616
rect 21460 5672 21588 5674
rect 21652 5674 21658 5676
rect 25681 5674 25747 5677
rect 25814 5674 25820 5676
rect 21460 5616 21546 5672
rect 21460 5614 21588 5616
rect 12341 5611 12407 5614
rect 18229 5611 18295 5614
rect 21541 5612 21588 5614
rect 21652 5614 25514 5674
rect 21652 5612 21658 5614
rect 21541 5611 21607 5612
rect 200 5538 800 5568
rect 1577 5538 1643 5541
rect 200 5536 1643 5538
rect 200 5480 1582 5536
rect 1638 5480 1643 5536
rect 200 5478 1643 5480
rect 200 5448 800 5478
rect 1577 5475 1643 5478
rect 3325 5538 3391 5541
rect 9213 5538 9279 5541
rect 3325 5536 9279 5538
rect 3325 5480 3330 5536
rect 3386 5480 9218 5536
rect 9274 5480 9279 5536
rect 3325 5478 9279 5480
rect 3325 5475 3391 5478
rect 9213 5475 9279 5478
rect 10593 5538 10659 5541
rect 15101 5538 15167 5541
rect 10593 5536 15167 5538
rect 10593 5480 10598 5536
rect 10654 5480 15106 5536
rect 15162 5480 15167 5536
rect 10593 5478 15167 5480
rect 10593 5475 10659 5478
rect 15101 5475 15167 5478
rect 20069 5538 20135 5541
rect 21725 5538 21791 5541
rect 20069 5536 21791 5538
rect 20069 5480 20074 5536
rect 20130 5480 21730 5536
rect 21786 5480 21791 5536
rect 20069 5478 21791 5480
rect 20069 5475 20135 5478
rect 21725 5475 21791 5478
rect 21909 5538 21975 5541
rect 22461 5538 22527 5541
rect 24025 5540 24091 5541
rect 23974 5538 23980 5540
rect 21909 5536 22527 5538
rect 21909 5480 21914 5536
rect 21970 5480 22466 5536
rect 22522 5480 22527 5536
rect 21909 5478 22527 5480
rect 23934 5478 23980 5538
rect 24044 5536 24091 5540
rect 24086 5480 24091 5536
rect 21909 5475 21975 5478
rect 22461 5475 22527 5478
rect 23974 5476 23980 5478
rect 24044 5476 24091 5480
rect 25454 5538 25514 5614
rect 25681 5672 25820 5674
rect 25681 5616 25686 5672
rect 25742 5616 25820 5672
rect 25681 5614 25820 5616
rect 25681 5611 25747 5614
rect 25814 5612 25820 5614
rect 25884 5612 25890 5676
rect 29361 5674 29427 5677
rect 26006 5672 29427 5674
rect 26006 5616 29366 5672
rect 29422 5616 29427 5672
rect 26006 5614 29427 5616
rect 26006 5538 26066 5614
rect 29361 5611 29427 5614
rect 25454 5478 26066 5538
rect 26325 5538 26391 5541
rect 28625 5538 28691 5541
rect 26325 5536 28691 5538
rect 26325 5480 26330 5536
rect 26386 5480 28630 5536
rect 28686 5480 28691 5536
rect 26325 5478 28691 5480
rect 24025 5475 24091 5476
rect 26325 5475 26391 5478
rect 28625 5475 28691 5478
rect 38193 5538 38259 5541
rect 39200 5538 39800 5568
rect 38193 5536 39800 5538
rect 38193 5480 38198 5536
rect 38254 5480 39800 5536
rect 38193 5478 39800 5480
rect 38193 5475 38259 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 39200 5448 39800 5478
rect 19570 5407 19886 5408
rect 1577 5402 1643 5405
rect 1894 5402 1900 5404
rect 1577 5400 1900 5402
rect 1577 5344 1582 5400
rect 1638 5344 1900 5400
rect 1577 5342 1900 5344
rect 1577 5339 1643 5342
rect 1894 5340 1900 5342
rect 1964 5340 1970 5404
rect 6821 5402 6887 5405
rect 7189 5402 7255 5405
rect 6821 5400 7255 5402
rect 6821 5344 6826 5400
rect 6882 5344 7194 5400
rect 7250 5344 7255 5400
rect 6821 5342 7255 5344
rect 6821 5339 6887 5342
rect 7189 5339 7255 5342
rect 7465 5402 7531 5405
rect 12801 5402 12867 5405
rect 7465 5400 12867 5402
rect 7465 5344 7470 5400
rect 7526 5344 12806 5400
rect 12862 5344 12867 5400
rect 7465 5342 12867 5344
rect 7465 5339 7531 5342
rect 12801 5339 12867 5342
rect 20529 5402 20595 5405
rect 26417 5402 26483 5405
rect 20529 5400 26483 5402
rect 20529 5344 20534 5400
rect 20590 5344 26422 5400
rect 26478 5344 26483 5400
rect 20529 5342 26483 5344
rect 20529 5339 20595 5342
rect 26417 5339 26483 5342
rect 3785 5266 3851 5269
rect 6913 5266 6979 5269
rect 3785 5264 6979 5266
rect 3785 5208 3790 5264
rect 3846 5208 6918 5264
rect 6974 5208 6979 5264
rect 3785 5206 6979 5208
rect 3785 5203 3851 5206
rect 6913 5203 6979 5206
rect 7189 5266 7255 5269
rect 10501 5266 10567 5269
rect 7189 5264 10567 5266
rect 7189 5208 7194 5264
rect 7250 5208 10506 5264
rect 10562 5208 10567 5264
rect 7189 5206 10567 5208
rect 7189 5203 7255 5206
rect 10501 5203 10567 5206
rect 16021 5266 16087 5269
rect 30373 5266 30439 5269
rect 16021 5264 30439 5266
rect 16021 5208 16026 5264
rect 16082 5208 30378 5264
rect 30434 5208 30439 5264
rect 16021 5206 30439 5208
rect 16021 5203 16087 5206
rect 30373 5203 30439 5206
rect 4521 5130 4587 5133
rect 9121 5130 9187 5133
rect 4521 5128 9187 5130
rect 4521 5072 4526 5128
rect 4582 5072 9126 5128
rect 9182 5072 9187 5128
rect 4521 5070 9187 5072
rect 4521 5067 4587 5070
rect 9121 5067 9187 5070
rect 14641 5130 14707 5133
rect 28349 5130 28415 5133
rect 14641 5128 28415 5130
rect 14641 5072 14646 5128
rect 14702 5072 28354 5128
rect 28410 5072 28415 5128
rect 14641 5070 28415 5072
rect 14641 5067 14707 5070
rect 28349 5067 28415 5070
rect 12065 4994 12131 4997
rect 13261 4994 13327 4997
rect 12065 4992 13327 4994
rect 12065 4936 12070 4992
rect 12126 4936 13266 4992
rect 13322 4936 13327 4992
rect 12065 4934 13327 4936
rect 12065 4931 12131 4934
rect 13261 4931 13327 4934
rect 21909 4994 21975 4997
rect 24577 4994 24643 4997
rect 28165 4994 28231 4997
rect 21909 4992 28231 4994
rect 21909 4936 21914 4992
rect 21970 4936 24582 4992
rect 24638 4936 28170 4992
rect 28226 4936 28231 4992
rect 21909 4934 28231 4936
rect 21909 4931 21975 4934
rect 24577 4931 24643 4934
rect 28165 4931 28231 4934
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 5073 4858 5139 4861
rect 12985 4858 13051 4861
rect 5073 4856 13051 4858
rect 5073 4800 5078 4856
rect 5134 4800 12990 4856
rect 13046 4800 13051 4856
rect 5073 4798 13051 4800
rect 5073 4795 5139 4798
rect 12985 4795 13051 4798
rect 19517 4858 19583 4861
rect 21909 4858 21975 4861
rect 19517 4856 21975 4858
rect 19517 4800 19522 4856
rect 19578 4800 21914 4856
rect 21970 4800 21975 4856
rect 19517 4798 21975 4800
rect 19517 4795 19583 4798
rect 21909 4795 21975 4798
rect 25037 4858 25103 4861
rect 28809 4858 28875 4861
rect 25037 4856 28875 4858
rect 25037 4800 25042 4856
rect 25098 4800 28814 4856
rect 28870 4800 28875 4856
rect 25037 4798 28875 4800
rect 25037 4795 25103 4798
rect 28809 4795 28875 4798
rect 3233 4722 3299 4725
rect 5993 4722 6059 4725
rect 3233 4720 6059 4722
rect 3233 4664 3238 4720
rect 3294 4664 5998 4720
rect 6054 4664 6059 4720
rect 3233 4662 6059 4664
rect 3233 4659 3299 4662
rect 5993 4659 6059 4662
rect 9121 4722 9187 4725
rect 27889 4722 27955 4725
rect 28349 4722 28415 4725
rect 9121 4720 28415 4722
rect 9121 4664 9126 4720
rect 9182 4664 27894 4720
rect 27950 4664 28354 4720
rect 28410 4664 28415 4720
rect 9121 4662 28415 4664
rect 9121 4659 9187 4662
rect 27889 4659 27955 4662
rect 28349 4659 28415 4662
rect 5717 4586 5783 4589
rect 14641 4586 14707 4589
rect 5717 4584 14707 4586
rect 5717 4528 5722 4584
rect 5778 4528 14646 4584
rect 14702 4528 14707 4584
rect 5717 4526 14707 4528
rect 5717 4523 5783 4526
rect 14641 4523 14707 4526
rect 14825 4586 14891 4589
rect 16021 4586 16087 4589
rect 14825 4584 16087 4586
rect 14825 4528 14830 4584
rect 14886 4528 16026 4584
rect 16082 4528 16087 4584
rect 14825 4526 16087 4528
rect 14825 4523 14891 4526
rect 16021 4523 16087 4526
rect 24761 4586 24827 4589
rect 26233 4586 26299 4589
rect 24761 4584 26299 4586
rect 24761 4528 24766 4584
rect 24822 4528 26238 4584
rect 26294 4528 26299 4584
rect 24761 4526 26299 4528
rect 24761 4523 24827 4526
rect 26233 4523 26299 4526
rect 26417 4586 26483 4589
rect 28717 4586 28783 4589
rect 26417 4584 28783 4586
rect 26417 4528 26422 4584
rect 26478 4528 28722 4584
rect 28778 4528 28783 4584
rect 26417 4526 28783 4528
rect 26417 4523 26483 4526
rect 28717 4523 28783 4526
rect 4797 4450 4863 4453
rect 9949 4450 10015 4453
rect 4797 4448 10015 4450
rect 4797 4392 4802 4448
rect 4858 4392 9954 4448
rect 10010 4392 10015 4448
rect 4797 4390 10015 4392
rect 4797 4387 4863 4390
rect 9949 4387 10015 4390
rect 21449 4450 21515 4453
rect 23841 4450 23907 4453
rect 21449 4448 23907 4450
rect 21449 4392 21454 4448
rect 21510 4392 23846 4448
rect 23902 4392 23907 4448
rect 21449 4390 23907 4392
rect 21449 4387 21515 4390
rect 23841 4387 23907 4390
rect 25497 4450 25563 4453
rect 30465 4450 30531 4453
rect 25497 4448 30531 4450
rect 25497 4392 25502 4448
rect 25558 4392 30470 4448
rect 30526 4392 30531 4448
rect 25497 4390 30531 4392
rect 25497 4387 25563 4390
rect 30465 4387 30531 4390
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 6177 4314 6243 4317
rect 4110 4312 6243 4314
rect 4110 4256 6182 4312
rect 6238 4256 6243 4312
rect 4110 4254 6243 4256
rect 200 4178 800 4208
rect 1761 4178 1827 4181
rect 200 4176 1827 4178
rect 200 4120 1766 4176
rect 1822 4120 1827 4176
rect 200 4118 1827 4120
rect 200 4088 800 4118
rect 1761 4115 1827 4118
rect 3785 4178 3851 4181
rect 3969 4178 4035 4181
rect 4110 4178 4170 4254
rect 6177 4251 6243 4254
rect 9489 4314 9555 4317
rect 12525 4314 12591 4317
rect 9489 4312 12591 4314
rect 9489 4256 9494 4312
rect 9550 4256 12530 4312
rect 12586 4256 12591 4312
rect 9489 4254 12591 4256
rect 9489 4251 9555 4254
rect 12525 4251 12591 4254
rect 20253 4314 20319 4317
rect 30373 4314 30439 4317
rect 20253 4312 30439 4314
rect 20253 4256 20258 4312
rect 20314 4256 30378 4312
rect 30434 4256 30439 4312
rect 20253 4254 30439 4256
rect 20253 4251 20319 4254
rect 30373 4251 30439 4254
rect 3785 4176 4170 4178
rect 3785 4120 3790 4176
rect 3846 4120 3974 4176
rect 4030 4120 4170 4176
rect 3785 4118 4170 4120
rect 7005 4178 7071 4181
rect 8293 4178 8359 4181
rect 7005 4176 8359 4178
rect 7005 4120 7010 4176
rect 7066 4120 8298 4176
rect 8354 4120 8359 4176
rect 7005 4118 8359 4120
rect 3785 4115 3851 4118
rect 3969 4115 4035 4118
rect 7005 4115 7071 4118
rect 8293 4115 8359 4118
rect 16205 4178 16271 4181
rect 17166 4178 17172 4180
rect 16205 4176 17172 4178
rect 16205 4120 16210 4176
rect 16266 4120 17172 4176
rect 16205 4118 17172 4120
rect 16205 4115 16271 4118
rect 17166 4116 17172 4118
rect 17236 4116 17242 4180
rect 18873 4178 18939 4181
rect 20989 4178 21055 4181
rect 21449 4178 21515 4181
rect 18873 4176 21515 4178
rect 18873 4120 18878 4176
rect 18934 4120 20994 4176
rect 21050 4120 21454 4176
rect 21510 4120 21515 4176
rect 18873 4118 21515 4120
rect 18873 4115 18939 4118
rect 20989 4115 21055 4118
rect 21449 4115 21515 4118
rect 21633 4178 21699 4181
rect 27613 4178 27679 4181
rect 21633 4176 27679 4178
rect 21633 4120 21638 4176
rect 21694 4120 27618 4176
rect 27674 4120 27679 4176
rect 21633 4118 27679 4120
rect 21633 4115 21699 4118
rect 27613 4115 27679 4118
rect 38101 4178 38167 4181
rect 39200 4178 39800 4208
rect 38101 4176 39800 4178
rect 38101 4120 38106 4176
rect 38162 4120 39800 4176
rect 38101 4118 39800 4120
rect 38101 4115 38167 4118
rect 39200 4088 39800 4118
rect 4153 4042 4219 4045
rect 14549 4042 14615 4045
rect 4153 4040 14615 4042
rect 4153 3984 4158 4040
rect 4214 3984 14554 4040
rect 14610 3984 14615 4040
rect 4153 3982 14615 3984
rect 4153 3979 4219 3982
rect 14549 3979 14615 3982
rect 18229 4042 18295 4045
rect 21817 4042 21883 4045
rect 18229 4040 21883 4042
rect 18229 3984 18234 4040
rect 18290 3984 21822 4040
rect 21878 3984 21883 4040
rect 18229 3982 21883 3984
rect 18229 3979 18295 3982
rect 21817 3979 21883 3982
rect 24117 4044 24183 4045
rect 24117 4040 24164 4044
rect 24228 4042 24234 4044
rect 24761 4042 24827 4045
rect 27981 4042 28047 4045
rect 24117 3984 24122 4040
rect 24117 3980 24164 3984
rect 24228 3982 24274 4042
rect 24761 4040 28047 4042
rect 24761 3984 24766 4040
rect 24822 3984 27986 4040
rect 28042 3984 28047 4040
rect 24761 3982 28047 3984
rect 24228 3980 24234 3982
rect 24117 3979 24183 3980
rect 24761 3979 24827 3982
rect 27981 3979 28047 3982
rect 29269 4042 29335 4045
rect 32489 4042 32555 4045
rect 29269 4040 32555 4042
rect 29269 3984 29274 4040
rect 29330 3984 32494 4040
rect 32550 3984 32555 4040
rect 29269 3982 32555 3984
rect 29269 3979 29335 3982
rect 32489 3979 32555 3982
rect 7925 3906 7991 3909
rect 8845 3906 8911 3909
rect 7925 3904 8911 3906
rect 7925 3848 7930 3904
rect 7986 3848 8850 3904
rect 8906 3848 8911 3904
rect 7925 3846 8911 3848
rect 7925 3843 7991 3846
rect 8845 3843 8911 3846
rect 11830 3844 11836 3908
rect 11900 3906 11906 3908
rect 16297 3906 16363 3909
rect 11900 3904 16363 3906
rect 11900 3848 16302 3904
rect 16358 3848 16363 3904
rect 11900 3846 16363 3848
rect 11900 3844 11906 3846
rect 16297 3843 16363 3846
rect 19374 3844 19380 3908
rect 19444 3844 19450 3908
rect 20069 3906 20135 3909
rect 29729 3906 29795 3909
rect 20069 3904 29795 3906
rect 20069 3848 20074 3904
rect 20130 3848 29734 3904
rect 29790 3848 29795 3904
rect 20069 3846 29795 3848
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 19382 3773 19442 3844
rect 20069 3843 20135 3846
rect 29729 3843 29795 3846
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 9489 3770 9555 3773
rect 10685 3770 10751 3773
rect 15694 3770 15700 3772
rect 9489 3768 10751 3770
rect 9489 3712 9494 3768
rect 9550 3712 10690 3768
rect 10746 3712 10751 3768
rect 9489 3710 10751 3712
rect 9489 3707 9555 3710
rect 10685 3707 10751 3710
rect 12390 3710 15700 3770
rect 2221 3634 2287 3637
rect 12390 3634 12450 3710
rect 15694 3708 15700 3710
rect 15764 3708 15770 3772
rect 19333 3768 19442 3773
rect 19333 3712 19338 3768
rect 19394 3712 19442 3768
rect 19333 3710 19442 3712
rect 19977 3770 20043 3773
rect 20110 3770 20116 3772
rect 19977 3768 20116 3770
rect 19977 3712 19982 3768
rect 20038 3712 20116 3768
rect 19977 3710 20116 3712
rect 19333 3707 19399 3710
rect 19977 3707 20043 3710
rect 20110 3708 20116 3710
rect 20180 3708 20186 3772
rect 22461 3770 22527 3773
rect 20302 3768 22527 3770
rect 20302 3712 22466 3768
rect 22522 3712 22527 3768
rect 20302 3710 22527 3712
rect 2221 3632 12450 3634
rect 2221 3576 2226 3632
rect 2282 3576 12450 3632
rect 2221 3574 12450 3576
rect 18413 3634 18479 3637
rect 19333 3634 19399 3637
rect 18413 3632 19399 3634
rect 18413 3576 18418 3632
rect 18474 3576 19338 3632
rect 19394 3576 19399 3632
rect 18413 3574 19399 3576
rect 2221 3571 2287 3574
rect 18413 3571 18479 3574
rect 19333 3571 19399 3574
rect 19517 3634 19583 3637
rect 20302 3634 20362 3710
rect 22461 3707 22527 3710
rect 23381 3770 23447 3773
rect 30281 3770 30347 3773
rect 23381 3768 30347 3770
rect 23381 3712 23386 3768
rect 23442 3712 30286 3768
rect 30342 3712 30347 3768
rect 23381 3710 30347 3712
rect 23381 3707 23447 3710
rect 30281 3707 30347 3710
rect 19517 3632 20362 3634
rect 19517 3576 19522 3632
rect 19578 3576 20362 3632
rect 19517 3574 20362 3576
rect 20529 3634 20595 3637
rect 30649 3634 30715 3637
rect 20529 3632 30715 3634
rect 20529 3576 20534 3632
rect 20590 3576 30654 3632
rect 30710 3576 30715 3632
rect 20529 3574 30715 3576
rect 19517 3571 19583 3574
rect 20529 3571 20595 3574
rect 30649 3571 30715 3574
rect 200 3498 800 3528
rect 1761 3498 1827 3501
rect 200 3496 1827 3498
rect 200 3440 1766 3496
rect 1822 3440 1827 3496
rect 200 3438 1827 3440
rect 200 3408 800 3438
rect 1761 3435 1827 3438
rect 4521 3498 4587 3501
rect 8385 3498 8451 3501
rect 4521 3496 8451 3498
rect 4521 3440 4526 3496
rect 4582 3440 8390 3496
rect 8446 3440 8451 3496
rect 4521 3438 8451 3440
rect 4521 3435 4587 3438
rect 8385 3435 8451 3438
rect 9397 3498 9463 3501
rect 19287 3498 19353 3501
rect 9397 3496 19353 3498
rect 9397 3440 9402 3496
rect 9458 3440 19292 3496
rect 19348 3440 19353 3496
rect 9397 3438 19353 3440
rect 9397 3435 9463 3438
rect 19287 3435 19353 3438
rect 19609 3498 19675 3501
rect 24669 3498 24735 3501
rect 26877 3498 26943 3501
rect 19609 3496 23122 3498
rect 19609 3440 19614 3496
rect 19670 3440 23122 3496
rect 19609 3438 23122 3440
rect 19609 3435 19675 3438
rect 3141 3362 3207 3365
rect 8569 3362 8635 3365
rect 3141 3360 8635 3362
rect 3141 3304 3146 3360
rect 3202 3304 8574 3360
rect 8630 3304 8635 3360
rect 3141 3302 8635 3304
rect 3141 3299 3207 3302
rect 8569 3299 8635 3302
rect 12617 3362 12683 3365
rect 16062 3362 16068 3364
rect 12617 3360 16068 3362
rect 12617 3304 12622 3360
rect 12678 3304 16068 3360
rect 12617 3302 16068 3304
rect 12617 3299 12683 3302
rect 16062 3300 16068 3302
rect 16132 3300 16138 3364
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 3141 3226 3207 3229
rect 15101 3226 15167 3229
rect 3141 3224 15167 3226
rect 3141 3168 3146 3224
rect 3202 3168 15106 3224
rect 15162 3168 15167 3224
rect 3141 3166 15167 3168
rect 3141 3163 3207 3166
rect 15101 3163 15167 3166
rect 2405 3090 2471 3093
rect 11881 3090 11947 3093
rect 13629 3090 13695 3093
rect 2405 3088 7620 3090
rect 2405 3032 2410 3088
rect 2466 3032 7620 3088
rect 2405 3030 7620 3032
rect 2405 3027 2471 3030
rect 7560 2818 7620 3030
rect 11881 3088 13695 3090
rect 11881 3032 11886 3088
rect 11942 3032 13634 3088
rect 13690 3032 13695 3088
rect 11881 3030 13695 3032
rect 11881 3027 11947 3030
rect 13629 3027 13695 3030
rect 14825 3090 14891 3093
rect 19609 3090 19675 3093
rect 14825 3088 19675 3090
rect 14825 3032 14830 3088
rect 14886 3032 19614 3088
rect 19670 3032 19675 3088
rect 14825 3030 19675 3032
rect 23062 3090 23122 3438
rect 24669 3496 26943 3498
rect 24669 3440 24674 3496
rect 24730 3440 26882 3496
rect 26938 3440 26943 3496
rect 24669 3438 26943 3440
rect 24669 3435 24735 3438
rect 26877 3435 26943 3438
rect 27061 3498 27127 3501
rect 28257 3498 28323 3501
rect 27061 3496 28323 3498
rect 27061 3440 27066 3496
rect 27122 3440 28262 3496
rect 28318 3440 28323 3496
rect 27061 3438 28323 3440
rect 27061 3435 27127 3438
rect 28257 3435 28323 3438
rect 38193 3498 38259 3501
rect 39200 3498 39800 3528
rect 38193 3496 39800 3498
rect 38193 3440 38198 3496
rect 38254 3440 39800 3496
rect 38193 3438 39800 3440
rect 38193 3435 38259 3438
rect 39200 3408 39800 3438
rect 23289 3362 23355 3365
rect 26233 3362 26299 3365
rect 23289 3360 26299 3362
rect 23289 3304 23294 3360
rect 23350 3304 26238 3360
rect 26294 3304 26299 3360
rect 23289 3302 26299 3304
rect 23289 3299 23355 3302
rect 26233 3299 26299 3302
rect 27245 3362 27311 3365
rect 31661 3362 31727 3365
rect 27245 3360 31727 3362
rect 27245 3304 27250 3360
rect 27306 3304 31666 3360
rect 31722 3304 31727 3360
rect 27245 3302 31727 3304
rect 27245 3299 27311 3302
rect 31661 3299 31727 3302
rect 26233 3226 26299 3229
rect 30465 3226 30531 3229
rect 26233 3224 30531 3226
rect 26233 3168 26238 3224
rect 26294 3168 30470 3224
rect 30526 3168 30531 3224
rect 26233 3166 30531 3168
rect 26233 3163 26299 3166
rect 30465 3163 30531 3166
rect 27337 3090 27403 3093
rect 30373 3090 30439 3093
rect 23062 3030 26802 3090
rect 14825 3027 14891 3030
rect 19609 3027 19675 3030
rect 11973 2954 12039 2957
rect 26509 2954 26575 2957
rect 11973 2952 26575 2954
rect 11973 2896 11978 2952
rect 12034 2896 26514 2952
rect 26570 2896 26575 2952
rect 11973 2894 26575 2896
rect 26742 2954 26802 3030
rect 27337 3088 30439 3090
rect 27337 3032 27342 3088
rect 27398 3032 30378 3088
rect 30434 3032 30439 3088
rect 27337 3030 30439 3032
rect 27337 3027 27403 3030
rect 30373 3027 30439 3030
rect 30833 2954 30899 2957
rect 26742 2952 30899 2954
rect 26742 2896 30838 2952
rect 30894 2896 30899 2952
rect 26742 2894 30899 2896
rect 11973 2891 12039 2894
rect 26509 2891 26575 2894
rect 30833 2891 30899 2894
rect 12617 2818 12683 2821
rect 7560 2816 12683 2818
rect 7560 2760 12622 2816
rect 12678 2760 12683 2816
rect 7560 2758 12683 2760
rect 12617 2755 12683 2758
rect 13353 2818 13419 2821
rect 20253 2818 20319 2821
rect 13353 2816 20319 2818
rect 13353 2760 13358 2816
rect 13414 2760 20258 2816
rect 20314 2760 20319 2816
rect 13353 2758 20319 2760
rect 13353 2755 13419 2758
rect 20253 2755 20319 2758
rect 26417 2818 26483 2821
rect 32397 2818 32463 2821
rect 26417 2816 32463 2818
rect 26417 2760 26422 2816
rect 26478 2760 32402 2816
rect 32458 2760 32463 2816
rect 26417 2758 32463 2760
rect 26417 2755 26483 2758
rect 32397 2755 32463 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 1669 2684 1735 2685
rect 3141 2684 3207 2685
rect 1669 2680 1716 2684
rect 1780 2682 1786 2684
rect 1669 2624 1674 2680
rect 1669 2620 1716 2624
rect 1780 2622 1826 2682
rect 3141 2680 3188 2684
rect 3252 2682 3258 2684
rect 14457 2682 14523 2685
rect 29177 2682 29243 2685
rect 3141 2624 3146 2680
rect 1780 2620 1786 2622
rect 3141 2620 3188 2624
rect 3252 2622 3298 2682
rect 14457 2680 29243 2682
rect 14457 2624 14462 2680
rect 14518 2624 29182 2680
rect 29238 2624 29243 2680
rect 14457 2622 29243 2624
rect 3252 2620 3258 2622
rect 1669 2619 1735 2620
rect 3141 2619 3207 2620
rect 14457 2619 14523 2622
rect 29177 2619 29243 2622
rect 19333 2546 19399 2549
rect 19609 2546 19675 2549
rect 19333 2544 19675 2546
rect 19333 2488 19338 2544
rect 19394 2488 19614 2544
rect 19670 2488 19675 2544
rect 19333 2486 19675 2488
rect 19333 2483 19399 2486
rect 19609 2483 19675 2486
rect 22737 2546 22803 2549
rect 29729 2546 29795 2549
rect 22737 2544 29795 2546
rect 22737 2488 22742 2544
rect 22798 2488 29734 2544
rect 29790 2488 29795 2544
rect 22737 2486 29795 2488
rect 22737 2483 22803 2486
rect 29729 2483 29795 2486
rect 19374 2348 19380 2412
rect 19444 2410 19450 2412
rect 19517 2410 19583 2413
rect 19444 2408 19583 2410
rect 19444 2352 19522 2408
rect 19578 2352 19583 2408
rect 19444 2350 19583 2352
rect 19444 2348 19450 2350
rect 19517 2347 19583 2350
rect 19701 2410 19767 2413
rect 21909 2410 21975 2413
rect 19701 2408 21975 2410
rect 19701 2352 19706 2408
rect 19762 2352 21914 2408
rect 21970 2352 21975 2408
rect 19701 2350 21975 2352
rect 19701 2347 19767 2350
rect 21909 2347 21975 2350
rect 11053 2276 11119 2277
rect 11053 2272 11100 2276
rect 11164 2274 11170 2276
rect 11053 2216 11058 2272
rect 11053 2212 11100 2216
rect 11164 2214 11210 2274
rect 11164 2212 11170 2214
rect 11053 2211 11119 2212
rect 19570 2208 19886 2209
rect 200 2138 800 2168
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 1853 2138 1919 2141
rect 200 2136 1919 2138
rect 200 2080 1858 2136
rect 1914 2080 1919 2136
rect 200 2078 1919 2080
rect 200 2048 800 2078
rect 1853 2075 1919 2078
rect 37181 2138 37247 2141
rect 39200 2138 39800 2168
rect 37181 2136 39800 2138
rect 37181 2080 37186 2136
rect 37242 2080 39800 2136
rect 37181 2078 39800 2080
rect 37181 2075 37247 2078
rect 39200 2048 39800 2078
rect 3049 914 3115 917
rect 1718 912 3115 914
rect 1718 856 3054 912
rect 3110 856 3115 912
rect 1718 854 3115 856
rect 200 778 800 808
rect 1718 778 1778 854
rect 3049 851 3115 854
rect 200 718 1778 778
rect 37825 778 37891 781
rect 39200 778 39800 808
rect 37825 776 39800 778
rect 37825 720 37830 776
rect 37886 720 39800 776
rect 37825 718 39800 720
rect 200 688 800 718
rect 37825 715 37891 718
rect 39200 688 39800 718
rect 37089 98 37155 101
rect 39200 98 39800 128
rect 37089 96 39800 98
rect 37089 40 37094 96
rect 37150 40 39800 96
rect 37089 38 39800 40
rect 37089 35 37155 38
rect 39200 8 39800 38
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 10548 25800 10612 25804
rect 10548 25744 10562 25800
rect 10562 25744 10612 25800
rect 10548 25740 10612 25744
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 3188 24244 3252 24308
rect 18460 23972 18524 24036
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 1716 23428 1780 23492
rect 15700 23488 15764 23492
rect 15700 23432 15714 23488
rect 15714 23432 15764 23488
rect 15700 23428 15764 23432
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 4844 20708 4908 20772
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 14412 20300 14476 20364
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 10916 19408 10980 19412
rect 10916 19352 10930 19408
rect 10930 19352 10980 19408
rect 10916 19348 10980 19352
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 11836 18668 11900 18732
rect 20116 18668 20180 18732
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 21588 18124 21652 18188
rect 17356 17988 17420 18052
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 8892 17580 8956 17644
rect 13676 17580 13740 17644
rect 20300 17580 20364 17644
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 19380 17036 19444 17100
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 11100 16764 11164 16828
rect 7972 16628 8036 16692
rect 13492 16628 13556 16692
rect 25820 16628 25884 16692
rect 12572 16356 12636 16420
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 13492 16008 13556 16012
rect 13492 15952 13506 16008
rect 13506 15952 13556 16008
rect 13492 15948 13556 15952
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 17172 15600 17236 15604
rect 17172 15544 17186 15600
rect 17186 15544 17236 15600
rect 17172 15540 17236 15544
rect 20484 15540 20548 15604
rect 13308 15268 13372 15332
rect 14596 15268 14660 15332
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 20668 15192 20732 15196
rect 20668 15136 20682 15192
rect 20682 15136 20732 15192
rect 20668 15132 20732 15136
rect 19380 14996 19444 15060
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 16068 14376 16132 14380
rect 16068 14320 16118 14376
rect 16118 14320 16132 14376
rect 16068 14316 16132 14320
rect 18644 14180 18708 14244
rect 20300 14180 20364 14244
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 1900 13772 1964 13836
rect 13676 13696 13740 13700
rect 13676 13640 13690 13696
rect 13690 13640 13740 13696
rect 13676 13636 13740 13640
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 10916 13500 10980 13564
rect 13492 13364 13556 13428
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 20484 12956 20548 13020
rect 10548 12820 10612 12884
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 18644 12140 18708 12204
rect 23980 12004 24044 12068
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 24164 11656 24228 11660
rect 24164 11600 24214 11656
rect 24214 11600 24228 11656
rect 24164 11596 24228 11600
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 12572 10236 12636 10300
rect 18460 10100 18524 10164
rect 20668 10100 20732 10164
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 14596 9556 14660 9620
rect 23980 9480 24044 9484
rect 23980 9424 24030 9480
rect 24030 9424 24044 9480
rect 23980 9420 24044 9424
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 14596 8876 14660 8940
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 8892 8664 8956 8668
rect 8892 8608 8906 8664
rect 8906 8608 8956 8664
rect 8892 8604 8956 8608
rect 17356 8604 17420 8668
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 4844 7924 4908 7988
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 13308 7244 13372 7308
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 18644 6292 18708 6356
rect 7972 6156 8036 6220
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 14412 5748 14476 5812
rect 21588 5672 21652 5676
rect 21588 5616 21602 5672
rect 21602 5616 21652 5672
rect 21588 5612 21652 5616
rect 23980 5536 24044 5540
rect 23980 5480 24030 5536
rect 24030 5480 24044 5536
rect 23980 5476 24044 5480
rect 25820 5612 25884 5676
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 1900 5340 1964 5404
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 17172 4116 17236 4180
rect 24164 4040 24228 4044
rect 24164 3984 24178 4040
rect 24178 3984 24228 4040
rect 24164 3980 24228 3984
rect 11836 3844 11900 3908
rect 19380 3844 19444 3908
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 15700 3708 15764 3772
rect 20116 3708 20180 3772
rect 16068 3300 16132 3364
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 1716 2680 1780 2684
rect 1716 2624 1730 2680
rect 1730 2624 1780 2680
rect 1716 2620 1780 2624
rect 3188 2680 3252 2684
rect 3188 2624 3202 2680
rect 3202 2624 3252 2680
rect 3188 2620 3252 2624
rect 19380 2348 19444 2412
rect 11100 2272 11164 2276
rect 11100 2216 11114 2272
rect 11114 2216 11164 2272
rect 11100 2212 11164 2216
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 10547 25804 10613 25805
rect 10547 25740 10548 25804
rect 10612 25740 10613 25804
rect 10547 25739 10613 25740
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 3187 24308 3253 24309
rect 3187 24244 3188 24308
rect 3252 24244 3253 24308
rect 3187 24243 3253 24244
rect 1715 23492 1781 23493
rect 1715 23428 1716 23492
rect 1780 23428 1781 23492
rect 1715 23427 1781 23428
rect 1718 2685 1778 23427
rect 1899 13836 1965 13837
rect 1899 13772 1900 13836
rect 1964 13772 1965 13836
rect 1899 13771 1965 13772
rect 1902 5405 1962 13771
rect 1899 5404 1965 5405
rect 1899 5340 1900 5404
rect 1964 5340 1965 5404
rect 1899 5339 1965 5340
rect 3190 2685 3250 24243
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4843 20772 4909 20773
rect 4843 20708 4844 20772
rect 4908 20708 4909 20772
rect 4843 20707 4909 20708
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4846 7989 4906 20707
rect 8891 17644 8957 17645
rect 8891 17580 8892 17644
rect 8956 17580 8957 17644
rect 8891 17579 8957 17580
rect 7971 16692 8037 16693
rect 7971 16628 7972 16692
rect 8036 16628 8037 16692
rect 7971 16627 8037 16628
rect 4843 7988 4909 7989
rect 4843 7924 4844 7988
rect 4908 7924 4909 7988
rect 4843 7923 4909 7924
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 7974 6221 8034 16627
rect 8894 8669 8954 17579
rect 10550 12885 10610 25739
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 18459 24036 18525 24037
rect 18459 23972 18460 24036
rect 18524 23972 18525 24036
rect 18459 23971 18525 23972
rect 15699 23492 15765 23493
rect 15699 23428 15700 23492
rect 15764 23428 15765 23492
rect 15699 23427 15765 23428
rect 14411 20364 14477 20365
rect 14411 20300 14412 20364
rect 14476 20300 14477 20364
rect 14411 20299 14477 20300
rect 10915 19412 10981 19413
rect 10915 19348 10916 19412
rect 10980 19348 10981 19412
rect 10915 19347 10981 19348
rect 10918 13565 10978 19347
rect 11835 18732 11901 18733
rect 11835 18668 11836 18732
rect 11900 18668 11901 18732
rect 11835 18667 11901 18668
rect 11099 16828 11165 16829
rect 11099 16764 11100 16828
rect 11164 16764 11165 16828
rect 11099 16763 11165 16764
rect 10915 13564 10981 13565
rect 10915 13500 10916 13564
rect 10980 13500 10981 13564
rect 10915 13499 10981 13500
rect 10547 12884 10613 12885
rect 10547 12820 10548 12884
rect 10612 12820 10613 12884
rect 10547 12819 10613 12820
rect 8891 8668 8957 8669
rect 8891 8604 8892 8668
rect 8956 8604 8957 8668
rect 8891 8603 8957 8604
rect 7971 6220 8037 6221
rect 7971 6156 7972 6220
rect 8036 6156 8037 6220
rect 7971 6155 8037 6156
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 1715 2684 1781 2685
rect 1715 2620 1716 2684
rect 1780 2620 1781 2684
rect 1715 2619 1781 2620
rect 3187 2684 3253 2685
rect 3187 2620 3188 2684
rect 3252 2620 3253 2684
rect 3187 2619 3253 2620
rect 4208 2128 4528 2688
rect 11102 2277 11162 16763
rect 11838 3909 11898 18667
rect 13675 17644 13741 17645
rect 13675 17580 13676 17644
rect 13740 17580 13741 17644
rect 13675 17579 13741 17580
rect 13491 16692 13557 16693
rect 13491 16628 13492 16692
rect 13556 16628 13557 16692
rect 13491 16627 13557 16628
rect 12571 16420 12637 16421
rect 12571 16356 12572 16420
rect 12636 16356 12637 16420
rect 12571 16355 12637 16356
rect 12574 10301 12634 16355
rect 13494 16013 13554 16627
rect 13491 16012 13557 16013
rect 13491 15948 13492 16012
rect 13556 15948 13557 16012
rect 13491 15947 13557 15948
rect 13307 15332 13373 15333
rect 13307 15268 13308 15332
rect 13372 15268 13373 15332
rect 13307 15267 13373 15268
rect 12571 10300 12637 10301
rect 12571 10236 12572 10300
rect 12636 10236 12637 10300
rect 12571 10235 12637 10236
rect 13310 7309 13370 15267
rect 13494 13429 13554 15947
rect 13678 13701 13738 17579
rect 13675 13700 13741 13701
rect 13675 13636 13676 13700
rect 13740 13636 13741 13700
rect 13675 13635 13741 13636
rect 13491 13428 13557 13429
rect 13491 13364 13492 13428
rect 13556 13364 13557 13428
rect 13491 13363 13557 13364
rect 13307 7308 13373 7309
rect 13307 7244 13308 7308
rect 13372 7244 13373 7308
rect 13307 7243 13373 7244
rect 14414 5813 14474 20299
rect 14595 15332 14661 15333
rect 14595 15268 14596 15332
rect 14660 15268 14661 15332
rect 14595 15267 14661 15268
rect 14598 9621 14658 15267
rect 14595 9620 14661 9621
rect 14595 9556 14596 9620
rect 14660 9556 14661 9620
rect 14595 9555 14661 9556
rect 14598 8941 14658 9555
rect 14595 8940 14661 8941
rect 14595 8876 14596 8940
rect 14660 8876 14661 8940
rect 14595 8875 14661 8876
rect 14411 5812 14477 5813
rect 14411 5748 14412 5812
rect 14476 5748 14477 5812
rect 14411 5747 14477 5748
rect 11835 3908 11901 3909
rect 11835 3844 11836 3908
rect 11900 3844 11901 3908
rect 11835 3843 11901 3844
rect 15702 3773 15762 23427
rect 17355 18052 17421 18053
rect 17355 17988 17356 18052
rect 17420 17988 17421 18052
rect 17355 17987 17421 17988
rect 17171 15604 17237 15605
rect 17171 15540 17172 15604
rect 17236 15540 17237 15604
rect 17171 15539 17237 15540
rect 16067 14380 16133 14381
rect 16067 14316 16068 14380
rect 16132 14316 16133 14380
rect 16067 14315 16133 14316
rect 15699 3772 15765 3773
rect 15699 3708 15700 3772
rect 15764 3708 15765 3772
rect 15699 3707 15765 3708
rect 16070 3365 16130 14315
rect 17174 4181 17234 15539
rect 17358 8669 17418 17987
rect 18462 10165 18522 23971
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 20115 18732 20181 18733
rect 20115 18668 20116 18732
rect 20180 18668 20181 18732
rect 20115 18667 20181 18668
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19379 17100 19445 17101
rect 19379 17036 19380 17100
rect 19444 17036 19445 17100
rect 19379 17035 19445 17036
rect 19382 15061 19442 17035
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19379 15060 19445 15061
rect 19379 14996 19380 15060
rect 19444 14996 19445 15060
rect 19379 14995 19445 14996
rect 18643 14244 18709 14245
rect 18643 14180 18644 14244
rect 18708 14180 18709 14244
rect 18643 14179 18709 14180
rect 18646 12205 18706 14179
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 18643 12204 18709 12205
rect 18643 12140 18644 12204
rect 18708 12140 18709 12204
rect 18643 12139 18709 12140
rect 18459 10164 18525 10165
rect 18459 10100 18460 10164
rect 18524 10100 18525 10164
rect 18459 10099 18525 10100
rect 17355 8668 17421 8669
rect 17355 8604 17356 8668
rect 17420 8604 17421 8668
rect 17355 8603 17421 8604
rect 18646 6357 18706 12139
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 18643 6356 18709 6357
rect 18643 6292 18644 6356
rect 18708 6292 18709 6356
rect 18643 6291 18709 6292
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 17171 4180 17237 4181
rect 17171 4116 17172 4180
rect 17236 4116 17237 4180
rect 17171 4115 17237 4116
rect 19379 3908 19445 3909
rect 19379 3844 19380 3908
rect 19444 3844 19445 3908
rect 19379 3843 19445 3844
rect 16067 3364 16133 3365
rect 16067 3300 16068 3364
rect 16132 3300 16133 3364
rect 16067 3299 16133 3300
rect 19382 2413 19442 3843
rect 19568 3296 19888 4320
rect 20118 3773 20178 18667
rect 21587 18188 21653 18189
rect 21587 18124 21588 18188
rect 21652 18124 21653 18188
rect 21587 18123 21653 18124
rect 20299 17644 20365 17645
rect 20299 17580 20300 17644
rect 20364 17580 20365 17644
rect 20299 17579 20365 17580
rect 20302 14245 20362 17579
rect 20483 15604 20549 15605
rect 20483 15540 20484 15604
rect 20548 15540 20549 15604
rect 20483 15539 20549 15540
rect 20299 14244 20365 14245
rect 20299 14180 20300 14244
rect 20364 14180 20365 14244
rect 20299 14179 20365 14180
rect 20486 13021 20546 15539
rect 20667 15196 20733 15197
rect 20667 15132 20668 15196
rect 20732 15132 20733 15196
rect 20667 15131 20733 15132
rect 20483 13020 20549 13021
rect 20483 12956 20484 13020
rect 20548 12956 20549 13020
rect 20483 12955 20549 12956
rect 20670 10165 20730 15131
rect 20667 10164 20733 10165
rect 20667 10100 20668 10164
rect 20732 10100 20733 10164
rect 20667 10099 20733 10100
rect 21590 5677 21650 18123
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 25819 16692 25885 16693
rect 25819 16628 25820 16692
rect 25884 16628 25885 16692
rect 25819 16627 25885 16628
rect 23979 12068 24045 12069
rect 23979 12004 23980 12068
rect 24044 12004 24045 12068
rect 23979 12003 24045 12004
rect 23982 9485 24042 12003
rect 24163 11660 24229 11661
rect 24163 11596 24164 11660
rect 24228 11596 24229 11660
rect 24163 11595 24229 11596
rect 23979 9484 24045 9485
rect 23979 9420 23980 9484
rect 24044 9420 24045 9484
rect 23979 9419 24045 9420
rect 21587 5676 21653 5677
rect 21587 5612 21588 5676
rect 21652 5612 21653 5676
rect 21587 5611 21653 5612
rect 23982 5541 24042 9419
rect 23979 5540 24045 5541
rect 23979 5476 23980 5540
rect 24044 5476 24045 5540
rect 23979 5475 24045 5476
rect 24166 4045 24226 11595
rect 25822 5677 25882 16627
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 25819 5676 25885 5677
rect 25819 5612 25820 5676
rect 25884 5612 25885 5676
rect 25819 5611 25885 5612
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 24163 4044 24229 4045
rect 24163 3980 24164 4044
rect 24228 3980 24229 4044
rect 24163 3979 24229 3980
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 20115 3772 20181 3773
rect 20115 3708 20116 3772
rect 20180 3708 20181 3772
rect 20115 3707 20181 3708
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19379 2412 19445 2413
rect 19379 2348 19380 2412
rect 19444 2348 19445 2412
rect 19379 2347 19445 2348
rect 11099 2276 11165 2277
rect 11099 2212 11100 2276
rect 11164 2212 11165 2276
rect 11099 2211 11165 2212
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 30360 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1667941163
transform 1 0 37996 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1667941163
transform 1 0 2116 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18
timestamp 1667941163
transform 1 0 2760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4140 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1667941163
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1667941163
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89
timestamp 1667941163
transform 1 0 9292 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1667941163
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117
timestamp 1667941163
transform 1 0 11868 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1667941163
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_145
timestamp 1667941163
transform 1 0 14444 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1667941163
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_173
timestamp 1667941163
transform 1 0 17020 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1667941163
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_219
timestamp 1667941163
transform 1 0 21252 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1667941163
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_230 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 22264 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_236
timestamp 1667941163
transform 1 0 22816 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1667941163
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_265
timestamp 1667941163
transform 1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1667941163
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_286
timestamp 1667941163
transform 1 0 27416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_294
timestamp 1667941163
transform 1 0 28152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1667941163
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1667941163
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_315
timestamp 1667941163
transform 1 0 30084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_323
timestamp 1667941163
transform 1 0 30820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_330
timestamp 1667941163
transform 1 0 31464 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_349
timestamp 1667941163
transform 1 0 33212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_357
timestamp 1667941163
transform 1 0 33948 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1667941163
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_371
timestamp 1667941163
transform 1 0 35236 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_377
timestamp 1667941163
transform 1 0 35788 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_382
timestamp 1667941163
transform 1 0 36248 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1667941163
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_405
timestamp 1667941163
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1667941163
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_16
timestamp 1667941163
transform 1 0 2576 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_23
timestamp 1667941163
transform 1 0 3220 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_30
timestamp 1667941163
transform 1 0 3864 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1667941163
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_63 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6900 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_71
timestamp 1667941163
transform 1 0 7636 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_96
timestamp 1667941163
transform 1 0 9936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_103
timestamp 1667941163
transform 1 0 10580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1667941163
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_117
timestamp 1667941163
transform 1 0 11868 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_121
timestamp 1667941163
transform 1 0 12236 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_129
timestamp 1667941163
transform 1 0 12972 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_154
timestamp 1667941163
transform 1 0 15272 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1667941163
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_193
timestamp 1667941163
transform 1 0 18860 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_218
timestamp 1667941163
transform 1 0 21160 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_247
timestamp 1667941163
transform 1 0 23828 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_264
timestamp 1667941163
transform 1 0 25392 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_277
timestamp 1667941163
transform 1 0 26588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_292
timestamp 1667941163
transform 1 0 27968 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_299
timestamp 1667941163
transform 1 0 28612 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_306
timestamp 1667941163
transform 1 0 29256 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_313
timestamp 1667941163
transform 1 0 29900 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_320
timestamp 1667941163
transform 1 0 30544 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_327
timestamp 1667941163
transform 1 0 31188 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_334
timestamp 1667941163
transform 1 0 31832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_342
timestamp 1667941163
transform 1 0 32568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_349
timestamp 1667941163
transform 1 0 33212 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_356 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 33856 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_368
timestamp 1667941163
transform 1 0 34960 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_377
timestamp 1667941163
transform 1 0 35788 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_385
timestamp 1667941163
transform 1 0 36524 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1667941163
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_9
timestamp 1667941163
transform 1 0 1932 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_13
timestamp 1667941163
transform 1 0 2300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_19
timestamp 1667941163
transform 1 0 2852 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1667941163
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_34
timestamp 1667941163
transform 1 0 4232 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_58
timestamp 1667941163
transform 1 0 6440 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1667941163
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_91
timestamp 1667941163
transform 1 0 9476 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_118
timestamp 1667941163
transform 1 0 11960 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_126
timestamp 1667941163
transform 1 0 12696 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1667941163
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_163
timestamp 1667941163
transform 1 0 16100 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_170
timestamp 1667941163
transform 1 0 16744 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1667941163
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_222
timestamp 1667941163
transform 1 0 21528 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_229
timestamp 1667941163
transform 1 0 22172 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_242
timestamp 1667941163
transform 1 0 23368 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_249
timestamp 1667941163
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_264
timestamp 1667941163
transform 1 0 25392 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_277
timestamp 1667941163
transform 1 0 26588 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_294
timestamp 1667941163
transform 1 0 28152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1667941163
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1667941163
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_314
timestamp 1667941163
transform 1 0 29992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_321
timestamp 1667941163
transform 1 0 30636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_328
timestamp 1667941163
transform 1 0 31280 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_335
timestamp 1667941163
transform 1 0 31924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_342
timestamp 1667941163
transform 1 0 32568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_349
timestamp 1667941163
transform 1 0 33212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_356
timestamp 1667941163
transform 1 0 33856 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1667941163
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1667941163
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_405
timestamp 1667941163
transform 1 0 38364 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_9
timestamp 1667941163
transform 1 0 1932 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_13
timestamp 1667941163
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_20
timestamp 1667941163
transform 1 0 2944 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 1667941163
transform 1 0 3588 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_34
timestamp 1667941163
transform 1 0 4232 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_41
timestamp 1667941163
transform 1 0 4876 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_49
timestamp 1667941163
transform 1 0 5612 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1667941163
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_88
timestamp 1667941163
transform 1 0 9200 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_94
timestamp 1667941163
transform 1 0 9752 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_106
timestamp 1667941163
transform 1 0 10856 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_117
timestamp 1667941163
transform 1 0 11868 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_138
timestamp 1667941163
transform 1 0 13800 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1667941163
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_183
timestamp 1667941163
transform 1 0 17940 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_208
timestamp 1667941163
transform 1 0 20240 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_215
timestamp 1667941163
transform 1 0 20884 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1667941163
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_231
timestamp 1667941163
transform 1 0 22356 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_235
timestamp 1667941163
transform 1 0 22724 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_252
timestamp 1667941163
transform 1 0 24288 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_265
timestamp 1667941163
transform 1 0 25484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1667941163
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_286
timestamp 1667941163
transform 1 0 27416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_293
timestamp 1667941163
transform 1 0 28060 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_300
timestamp 1667941163
transform 1 0 28704 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_307
timestamp 1667941163
transform 1 0 29348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_314
timestamp 1667941163
transform 1 0 29992 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_321
timestamp 1667941163
transform 1 0 30636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_328
timestamp 1667941163
transform 1 0 31280 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_342
timestamp 1667941163
transform 1 0 32568 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_357
timestamp 1667941163
transform 1 0 33948 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_369
timestamp 1667941163
transform 1 0 35052 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_381
timestamp 1667941163
transform 1 0 36156 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_389
timestamp 1667941163
transform 1 0 36892 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_401
timestamp 1667941163
transform 1 0 37996 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_9
timestamp 1667941163
transform 1 0 1932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_15
timestamp 1667941163
transform 1 0 2484 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_19
timestamp 1667941163
transform 1 0 2852 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1667941163
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_57
timestamp 1667941163
transform 1 0 6348 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1667941163
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1667941163
transform 1 0 9476 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_112
timestamp 1667941163
transform 1 0 11408 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_137
timestamp 1667941163
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_145
timestamp 1667941163
transform 1 0 14444 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_166
timestamp 1667941163
transform 1 0 16376 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_172
timestamp 1667941163
transform 1 0 16928 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp 1667941163
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_220
timestamp 1667941163
transform 1 0 21344 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_244
timestamp 1667941163
transform 1 0 23552 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_257
timestamp 1667941163
transform 1 0 24748 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_271
timestamp 1667941163
transform 1 0 26036 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_275
timestamp 1667941163
transform 1 0 26404 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_289
timestamp 1667941163
transform 1 0 27692 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_296
timestamp 1667941163
transform 1 0 28336 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_303
timestamp 1667941163
transform 1 0 28980 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1667941163
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_314
timestamp 1667941163
transform 1 0 29992 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_328
timestamp 1667941163
transform 1 0 31280 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_335
timestamp 1667941163
transform 1 0 31924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_342
timestamp 1667941163
transform 1 0 32568 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_350
timestamp 1667941163
transform 1 0 33304 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_355
timestamp 1667941163
transform 1 0 33764 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1667941163
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1667941163
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_405
timestamp 1667941163
transform 1 0 38364 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_8
timestamp 1667941163
transform 1 0 1840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_12
timestamp 1667941163
transform 1 0 2208 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_16
timestamp 1667941163
transform 1 0 2576 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_23
timestamp 1667941163
transform 1 0 3220 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_30
timestamp 1667941163
transform 1 0 3864 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1667941163
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_62
timestamp 1667941163
transform 1 0 6808 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_86
timestamp 1667941163
transform 1 0 9016 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1667941163
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_138
timestamp 1667941163
transform 1 0 13800 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_162
timestamp 1667941163
transform 1 0 16008 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_192
timestamp 1667941163
transform 1 0 18768 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_220
timestamp 1667941163
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_231
timestamp 1667941163
transform 1 0 22356 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_235
timestamp 1667941163
transform 1 0 22724 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_252
timestamp 1667941163
transform 1 0 24288 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_259
timestamp 1667941163
transform 1 0 24932 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_278
timestamp 1667941163
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_286
timestamp 1667941163
transform 1 0 27416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_293
timestamp 1667941163
transform 1 0 28060 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_300
timestamp 1667941163
transform 1 0 28704 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_307
timestamp 1667941163
transform 1 0 29348 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_314
timestamp 1667941163
transform 1 0 29992 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_321
timestamp 1667941163
transform 1 0 30636 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_333
timestamp 1667941163
transform 1 0 31740 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1667941163
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1667941163
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1667941163
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1667941163
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1667941163
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1667941163
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_12
timestamp 1667941163
transform 1 0 2208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_19
timestamp 1667941163
transform 1 0 2852 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1667941163
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_57
timestamp 1667941163
transform 1 0 6348 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1667941163
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_109
timestamp 1667941163
transform 1 0 11132 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_117
timestamp 1667941163
transform 1 0 11868 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1667941163
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_164
timestamp 1667941163
transform 1 0 16192 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_172
timestamp 1667941163
transform 1 0 16928 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1667941163
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_224
timestamp 1667941163
transform 1 0 21712 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_233
timestamp 1667941163
transform 1 0 22540 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_246
timestamp 1667941163
transform 1 0 23736 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_268
timestamp 1667941163
transform 1 0 25760 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_275
timestamp 1667941163
transform 1 0 26404 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_282
timestamp 1667941163
transform 1 0 27048 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_289
timestamp 1667941163
transform 1 0 27692 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_296
timestamp 1667941163
transform 1 0 28336 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_303
timestamp 1667941163
transform 1 0 28980 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1667941163
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_314
timestamp 1667941163
transform 1 0 29992 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_326
timestamp 1667941163
transform 1 0 31096 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_338
timestamp 1667941163
transform 1 0 32200 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_350
timestamp 1667941163
transform 1 0 33304 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_362
timestamp 1667941163
transform 1 0 34408 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1667941163
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1667941163
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_405
timestamp 1667941163
transform 1 0 38364 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_14
timestamp 1667941163
transform 1 0 2392 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_31
timestamp 1667941163
transform 1 0 3956 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_40
timestamp 1667941163
transform 1 0 4784 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_47
timestamp 1667941163
transform 1 0 5428 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1667941163
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_70
timestamp 1667941163
transform 1 0 7544 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_74
timestamp 1667941163
transform 1 0 7912 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_78
timestamp 1667941163
transform 1 0 8280 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_103
timestamp 1667941163
transform 1 0 10580 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1667941163
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_136
timestamp 1667941163
transform 1 0 13616 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_160
timestamp 1667941163
transform 1 0 15824 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_195
timestamp 1667941163
transform 1 0 19044 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_201
timestamp 1667941163
transform 1 0 19596 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1667941163
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_235
timestamp 1667941163
transform 1 0 22724 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_243
timestamp 1667941163
transform 1 0 23460 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_257
timestamp 1667941163
transform 1 0 24748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_261
timestamp 1667941163
transform 1 0 25116 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_275
timestamp 1667941163
transform 1 0 26404 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1667941163
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_287
timestamp 1667941163
transform 1 0 27508 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_294
timestamp 1667941163
transform 1 0 28152 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_301
timestamp 1667941163
transform 1 0 28796 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_313
timestamp 1667941163
transform 1 0 29900 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1667941163
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1667941163
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1667941163
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1667941163
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1667941163
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1667941163
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_385
timestamp 1667941163
transform 1 0 36524 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_389
timestamp 1667941163
transform 1 0 36892 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_8
timestamp 1667941163
transform 1 0 1840 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_20
timestamp 1667941163
transform 1 0 2944 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_33
timestamp 1667941163
transform 1 0 4140 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_37
timestamp 1667941163
transform 1 0 4508 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_44
timestamp 1667941163
transform 1 0 5152 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_51
timestamp 1667941163
transform 1 0 5796 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_58
timestamp 1667941163
transform 1 0 6440 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1667941163
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_96
timestamp 1667941163
transform 1 0 9936 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_111
timestamp 1667941163
transform 1 0 11316 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_135
timestamp 1667941163
transform 1 0 13524 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1667941163
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_165
timestamp 1667941163
transform 1 0 16284 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1667941163
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_201
timestamp 1667941163
transform 1 0 19596 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_222
timestamp 1667941163
transform 1 0 21528 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_229
timestamp 1667941163
transform 1 0 22172 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_236
timestamp 1667941163
transform 1 0 22816 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_243
timestamp 1667941163
transform 1 0 23460 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1667941163
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_257
timestamp 1667941163
transform 1 0 24748 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_271
timestamp 1667941163
transform 1 0 26036 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_288
timestamp 1667941163
transform 1 0 27600 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_295
timestamp 1667941163
transform 1 0 28244 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_302
timestamp 1667941163
transform 1 0 28888 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1667941163
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1667941163
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1667941163
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1667941163
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1667941163
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1667941163
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_401
timestamp 1667941163
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_17
timestamp 1667941163
transform 1 0 2668 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_26
timestamp 1667941163
transform 1 0 3496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_33
timestamp 1667941163
transform 1 0 4140 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_40
timestamp 1667941163
transform 1 0 4784 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_47
timestamp 1667941163
transform 1 0 5428 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1667941163
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_85
timestamp 1667941163
transform 1 0 8924 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1667941163
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_138
timestamp 1667941163
transform 1 0 13800 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_162
timestamp 1667941163
transform 1 0 16008 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_174
timestamp 1667941163
transform 1 0 17112 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_198
timestamp 1667941163
transform 1 0 19320 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1667941163
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_238
timestamp 1667941163
transform 1 0 23000 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_246
timestamp 1667941163
transform 1 0 23736 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_256
timestamp 1667941163
transform 1 0 24656 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_263
timestamp 1667941163
transform 1 0 25300 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_270
timestamp 1667941163
transform 1 0 25944 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp 1667941163
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_286
timestamp 1667941163
transform 1 0 27416 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1667941163
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1667941163
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1667941163
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1667941163
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1667941163
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_357
timestamp 1667941163
transform 1 0 33948 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_363
timestamp 1667941163
transform 1 0 34500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_375
timestamp 1667941163
transform 1 0 35604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_387
timestamp 1667941163
transform 1 0 36708 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1667941163
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_401
timestamp 1667941163
transform 1 0 37996 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_12
timestamp 1667941163
transform 1 0 2208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_19
timestamp 1667941163
transform 1 0 2852 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1667941163
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_34
timestamp 1667941163
transform 1 0 4232 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_38
timestamp 1667941163
transform 1 0 4600 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_42
timestamp 1667941163
transform 1 0 4968 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_49
timestamp 1667941163
transform 1 0 5612 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_56
timestamp 1667941163
transform 1 0 6256 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_60
timestamp 1667941163
transform 1 0 6624 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1667941163
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_108
timestamp 1667941163
transform 1 0 11040 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_116
timestamp 1667941163
transform 1 0 11776 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1667941163
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_167
timestamp 1667941163
transform 1 0 16468 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_173
timestamp 1667941163
transform 1 0 17020 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1667941163
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_225
timestamp 1667941163
transform 1 0 21804 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_237
timestamp 1667941163
transform 1 0 22908 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_243
timestamp 1667941163
transform 1 0 23460 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1667941163
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_258
timestamp 1667941163
transform 1 0 24840 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_265
timestamp 1667941163
transform 1 0 25484 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_271
timestamp 1667941163
transform 1 0 26036 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_285
timestamp 1667941163
transform 1 0 27324 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_292
timestamp 1667941163
transform 1 0 27968 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_304
timestamp 1667941163
transform 1 0 29072 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1667941163
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1667941163
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1667941163
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1667941163
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1667941163
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_389
timestamp 1667941163
transform 1 0 36892 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_405
timestamp 1667941163
transform 1 0 38364 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_8
timestamp 1667941163
transform 1 0 1840 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_15
timestamp 1667941163
transform 1 0 2484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_22
timestamp 1667941163
transform 1 0 3128 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_26
timestamp 1667941163
transform 1 0 3496 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_30
timestamp 1667941163
transform 1 0 3864 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1667941163
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_62
timestamp 1667941163
transform 1 0 6808 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_77
timestamp 1667941163
transform 1 0 8188 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_102
timestamp 1667941163
transform 1 0 10488 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_106
timestamp 1667941163
transform 1 0 10856 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1667941163
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_124
timestamp 1667941163
transform 1 0 12512 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_151
timestamp 1667941163
transform 1 0 14996 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1667941163
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_191
timestamp 1667941163
transform 1 0 18676 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_218
timestamp 1667941163
transform 1 0 21160 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_233
timestamp 1667941163
transform 1 0 22540 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_239
timestamp 1667941163
transform 1 0 23092 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_248
timestamp 1667941163
transform 1 0 23920 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_255
timestamp 1667941163
transform 1 0 24564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_262
timestamp 1667941163
transform 1 0 25208 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_268
timestamp 1667941163
transform 1 0 25760 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_272
timestamp 1667941163
transform 1 0 26128 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_286
timestamp 1667941163
transform 1 0 27416 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_294
timestamp 1667941163
transform 1 0 28152 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_300
timestamp 1667941163
transform 1 0 28704 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_314
timestamp 1667941163
transform 1 0 29992 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_321
timestamp 1667941163
transform 1 0 30636 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_333
timestamp 1667941163
transform 1 0 31740 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1667941163
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1667941163
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1667941163
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1667941163
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_9
timestamp 1667941163
transform 1 0 1932 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_16
timestamp 1667941163
transform 1 0 2576 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_20
timestamp 1667941163
transform 1 0 2944 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1667941163
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_36
timestamp 1667941163
transform 1 0 4416 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_43
timestamp 1667941163
transform 1 0 5060 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_58
timestamp 1667941163
transform 1 0 6440 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1667941163
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_107
timestamp 1667941163
transform 1 0 10948 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_132
timestamp 1667941163
transform 1 0 13248 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_164
timestamp 1667941163
transform 1 0 16192 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_171
timestamp 1667941163
transform 1 0 16836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1667941163
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_224
timestamp 1667941163
transform 1 0 21712 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_236
timestamp 1667941163
transform 1 0 22816 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_240
timestamp 1667941163
transform 1 0 23184 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_247
timestamp 1667941163
transform 1 0 23828 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1667941163
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_257
timestamp 1667941163
transform 1 0 24748 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_271
timestamp 1667941163
transform 1 0 26036 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_283
timestamp 1667941163
transform 1 0 27140 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_295
timestamp 1667941163
transform 1 0 28244 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_302
timestamp 1667941163
transform 1 0 28888 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_319
timestamp 1667941163
transform 1 0 30452 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_326
timestamp 1667941163
transform 1 0 31096 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_338
timestamp 1667941163
transform 1 0 32200 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_350
timestamp 1667941163
transform 1 0 33304 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_362
timestamp 1667941163
transform 1 0 34408 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1667941163
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_401
timestamp 1667941163
transform 1 0 37996 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_405
timestamp 1667941163
transform 1 0 38364 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_9
timestamp 1667941163
transform 1 0 1932 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_16
timestamp 1667941163
transform 1 0 2576 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_22
timestamp 1667941163
transform 1 0 3128 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_26
timestamp 1667941163
transform 1 0 3496 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_33
timestamp 1667941163
transform 1 0 4140 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_40
timestamp 1667941163
transform 1 0 4784 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_49
timestamp 1667941163
transform 1 0 5612 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1667941163
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_69
timestamp 1667941163
transform 1 0 7452 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_92
timestamp 1667941163
transform 1 0 9568 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_98
timestamp 1667941163
transform 1 0 10120 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1667941163
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_118
timestamp 1667941163
transform 1 0 11960 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_143
timestamp 1667941163
transform 1 0 14260 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_158
timestamp 1667941163
transform 1 0 15640 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_165
timestamp 1667941163
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_195
timestamp 1667941163
transform 1 0 19044 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_219
timestamp 1667941163
transform 1 0 21252 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1667941163
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_237
timestamp 1667941163
transform 1 0 22908 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_243
timestamp 1667941163
transform 1 0 23460 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_257
timestamp 1667941163
transform 1 0 24748 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_269
timestamp 1667941163
transform 1 0 25852 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_277
timestamp 1667941163
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1667941163
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_305
timestamp 1667941163
transform 1 0 29164 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_310
timestamp 1667941163
transform 1 0 29624 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_314
timestamp 1667941163
transform 1 0 29992 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_318
timestamp 1667941163
transform 1 0 30360 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_325
timestamp 1667941163
transform 1 0 31004 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_332
timestamp 1667941163
transform 1 0 31648 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1667941163
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1667941163
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1667941163
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1667941163
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_12
timestamp 1667941163
transform 1 0 2208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_19
timestamp 1667941163
transform 1 0 2852 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1667941163
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_34
timestamp 1667941163
transform 1 0 4232 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_46
timestamp 1667941163
transform 1 0 5336 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_58
timestamp 1667941163
transform 1 0 6440 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1667941163
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_113
timestamp 1667941163
transform 1 0 11500 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1667941163
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_149
timestamp 1667941163
transform 1 0 14812 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_153
timestamp 1667941163
transform 1 0 15180 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_161
timestamp 1667941163
transform 1 0 15916 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_185
timestamp 1667941163
transform 1 0 18124 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_192
timestamp 1667941163
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_223
timestamp 1667941163
transform 1 0 21620 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_235
timestamp 1667941163
transform 1 0 22724 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_241
timestamp 1667941163
transform 1 0 23276 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_249
timestamp 1667941163
transform 1 0 24012 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_268
timestamp 1667941163
transform 1 0 25760 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_280
timestamp 1667941163
transform 1 0 26864 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_292
timestamp 1667941163
transform 1 0 27968 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_304
timestamp 1667941163
transform 1 0 29072 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1667941163
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1667941163
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1667941163
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1667941163
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1667941163
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_389
timestamp 1667941163
transform 1 0 36892 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_397
timestamp 1667941163
transform 1 0 37628 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_402
timestamp 1667941163
transform 1 0 38088 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_406
timestamp 1667941163
transform 1 0 38456 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_8
timestamp 1667941163
transform 1 0 1840 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_19
timestamp 1667941163
transform 1 0 2852 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_27
timestamp 1667941163
transform 1 0 3588 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_31
timestamp 1667941163
transform 1 0 3956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_43
timestamp 1667941163
transform 1 0 5060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1667941163
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_65
timestamp 1667941163
transform 1 0 7084 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_88
timestamp 1667941163
transform 1 0 9200 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_96
timestamp 1667941163
transform 1 0 9936 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_101
timestamp 1667941163
transform 1 0 10396 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 1667941163
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_122
timestamp 1667941163
transform 1 0 12328 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_129
timestamp 1667941163
transform 1 0 12972 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_154
timestamp 1667941163
transform 1 0 15272 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1667941163
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_193
timestamp 1667941163
transform 1 0 18860 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1667941163
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1667941163
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_236
timestamp 1667941163
transform 1 0 22816 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_257
timestamp 1667941163
transform 1 0 24748 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_268
timestamp 1667941163
transform 1 0 25760 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1667941163
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_305
timestamp 1667941163
transform 1 0 29164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_309
timestamp 1667941163
transform 1 0 29532 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_321
timestamp 1667941163
transform 1 0 30636 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_333
timestamp 1667941163
transform 1 0 31740 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_364
timestamp 1667941163
transform 1 0 34592 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1667941163
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1667941163
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1667941163
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_8
timestamp 1667941163
transform 1 0 1840 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_12
timestamp 1667941163
transform 1 0 2208 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_16
timestamp 1667941163
transform 1 0 2576 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1667941163
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_53
timestamp 1667941163
transform 1 0 5980 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_61
timestamp 1667941163
transform 1 0 6716 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1667941163
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_111
timestamp 1667941163
transform 1 0 11316 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1667941163
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_166
timestamp 1667941163
transform 1 0 16376 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_190
timestamp 1667941163
transform 1 0 18584 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_210
timestamp 1667941163
transform 1 0 20424 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_222
timestamp 1667941163
transform 1 0 21528 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_234
timestamp 1667941163
transform 1 0 22632 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_238
timestamp 1667941163
transform 1 0 23000 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_242
timestamp 1667941163
transform 1 0 23368 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_249
timestamp 1667941163
transform 1 0 24012 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_259
timestamp 1667941163
transform 1 0 24932 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_269
timestamp 1667941163
transform 1 0 25852 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_276
timestamp 1667941163
transform 1 0 26496 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_288
timestamp 1667941163
transform 1 0 27600 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_293
timestamp 1667941163
transform 1 0 28060 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_305
timestamp 1667941163
transform 1 0 29164 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_314
timestamp 1667941163
transform 1 0 29992 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_326
timestamp 1667941163
transform 1 0 31096 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_338
timestamp 1667941163
transform 1 0 32200 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_350
timestamp 1667941163
transform 1 0 33304 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_362
timestamp 1667941163
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_389
timestamp 1667941163
transform 1 0 36892 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_393
timestamp 1667941163
transform 1 0 37260 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_397
timestamp 1667941163
transform 1 0 37628 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_405
timestamp 1667941163
transform 1 0 38364 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1667941163
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1667941163
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1667941163
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1667941163
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1667941163
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_69
timestamp 1667941163
transform 1 0 7452 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_73
timestamp 1667941163
transform 1 0 7820 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_97
timestamp 1667941163
transform 1 0 10028 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_105
timestamp 1667941163
transform 1 0 10764 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1667941163
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_136
timestamp 1667941163
transform 1 0 13616 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_160
timestamp 1667941163
transform 1 0 15824 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_173
timestamp 1667941163
transform 1 0 17020 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_195
timestamp 1667941163
transform 1 0 19044 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1667941163
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_229
timestamp 1667941163
transform 1 0 22172 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_233
timestamp 1667941163
transform 1 0 22540 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_252
timestamp 1667941163
transform 1 0 24288 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_259
timestamp 1667941163
transform 1 0 24932 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_276
timestamp 1667941163
transform 1 0 26496 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_292
timestamp 1667941163
transform 1 0 27968 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_304
timestamp 1667941163
transform 1 0 29072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_315
timestamp 1667941163
transform 1 0 30084 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_322
timestamp 1667941163
transform 1 0 30728 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_334
timestamp 1667941163
transform 1 0 31832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_342
timestamp 1667941163
transform 1 0 32568 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_354
timestamp 1667941163
transform 1 0 33672 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_366
timestamp 1667941163
transform 1 0 34776 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_378
timestamp 1667941163
transform 1 0 35880 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_390
timestamp 1667941163
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1667941163
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1667941163
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1667941163
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_53
timestamp 1667941163
transform 1 0 5980 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1667941163
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_90
timestamp 1667941163
transform 1 0 9384 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_97
timestamp 1667941163
transform 1 0 10028 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_124
timestamp 1667941163
transform 1 0 12512 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_131
timestamp 1667941163
transform 1 0 13156 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1667941163
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_147
timestamp 1667941163
transform 1 0 14628 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_154
timestamp 1667941163
transform 1 0 15272 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_160
timestamp 1667941163
transform 1 0 15824 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_184
timestamp 1667941163
transform 1 0 18032 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_191
timestamp 1667941163
transform 1 0 18676 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1667941163
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_228
timestamp 1667941163
transform 1 0 22080 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_249
timestamp 1667941163
transform 1 0 24012 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_263
timestamp 1667941163
transform 1 0 25300 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_270
timestamp 1667941163
transform 1 0 25944 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1667941163
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_289
timestamp 1667941163
transform 1 0 27692 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_295
timestamp 1667941163
transform 1 0 28244 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_299
timestamp 1667941163
transform 1 0 28612 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1667941163
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_316
timestamp 1667941163
transform 1 0 30176 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_328
timestamp 1667941163
transform 1 0 31280 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_340
timestamp 1667941163
transform 1 0 32384 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_352
timestamp 1667941163
transform 1 0 33488 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1667941163
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_401
timestamp 1667941163
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_9
timestamp 1667941163
transform 1 0 1932 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_21
timestamp 1667941163
transform 1 0 3036 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_29
timestamp 1667941163
transform 1 0 3772 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_34
timestamp 1667941163
transform 1 0 4232 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_42
timestamp 1667941163
transform 1 0 4968 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_47
timestamp 1667941163
transform 1 0 5428 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1667941163
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_68
timestamp 1667941163
transform 1 0 7360 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_93
timestamp 1667941163
transform 1 0 9660 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_97
timestamp 1667941163
transform 1 0 10028 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_104
timestamp 1667941163
transform 1 0 10672 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_140
timestamp 1667941163
transform 1 0 13984 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_144
timestamp 1667941163
transform 1 0 14352 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1667941163
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_191
timestamp 1667941163
transform 1 0 18676 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1667941163
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_234
timestamp 1667941163
transform 1 0 22632 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_241
timestamp 1667941163
transform 1 0 23276 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_249
timestamp 1667941163
transform 1 0 24012 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_259
timestamp 1667941163
transform 1 0 24932 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_275
timestamp 1667941163
transform 1 0 26404 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1667941163
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_289
timestamp 1667941163
transform 1 0 27692 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_300
timestamp 1667941163
transform 1 0 28704 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_307
timestamp 1667941163
transform 1 0 29348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_319
timestamp 1667941163
transform 1 0 30452 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1667941163
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1667941163
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1667941163
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1667941163
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1667941163
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1667941163
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1667941163
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1667941163
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1667941163
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_40
timestamp 1667941163
transform 1 0 4784 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_47
timestamp 1667941163
transform 1 0 5428 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_54
timestamp 1667941163
transform 1 0 6072 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1667941163
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_107
timestamp 1667941163
transform 1 0 10948 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_115
timestamp 1667941163
transform 1 0 11684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1667941163
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_164
timestamp 1667941163
transform 1 0 16192 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_188
timestamp 1667941163
transform 1 0 18400 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_220
timestamp 1667941163
transform 1 0 21344 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_227
timestamp 1667941163
transform 1 0 21988 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_234
timestamp 1667941163
transform 1 0 22632 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_238
timestamp 1667941163
transform 1 0 23000 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_248
timestamp 1667941163
transform 1 0 23920 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_264
timestamp 1667941163
transform 1 0 25392 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_276
timestamp 1667941163
transform 1 0 26496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_286
timestamp 1667941163
transform 1 0 27416 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_293
timestamp 1667941163
transform 1 0 28060 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_297
timestamp 1667941163
transform 1 0 28428 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_306
timestamp 1667941163
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_314
timestamp 1667941163
transform 1 0 29992 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_325
timestamp 1667941163
transform 1 0 31004 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_337
timestamp 1667941163
transform 1 0 32108 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_349
timestamp 1667941163
transform 1 0 33212 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_361
timestamp 1667941163
transform 1 0 34316 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_401
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_9
timestamp 1667941163
transform 1 0 1932 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_17
timestamp 1667941163
transform 1 0 2668 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_23
timestamp 1667941163
transform 1 0 3220 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_30
timestamp 1667941163
transform 1 0 3864 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_37
timestamp 1667941163
transform 1 0 4508 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_44
timestamp 1667941163
transform 1 0 5152 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_50
timestamp 1667941163
transform 1 0 5704 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1667941163
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_61
timestamp 1667941163
transform 1 0 6716 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_65
timestamp 1667941163
transform 1 0 7084 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_89
timestamp 1667941163
transform 1 0 9292 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_97
timestamp 1667941163
transform 1 0 10028 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1667941163
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_120
timestamp 1667941163
transform 1 0 12144 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_144
timestamp 1667941163
transform 1 0 14352 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1667941163
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1667941163
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_177
timestamp 1667941163
transform 1 0 17388 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_188
timestamp 1667941163
transform 1 0 18400 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_212
timestamp 1667941163
transform 1 0 20608 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_216
timestamp 1667941163
transform 1 0 20976 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_220
timestamp 1667941163
transform 1 0 21344 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_229
timestamp 1667941163
transform 1 0 22172 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_243
timestamp 1667941163
transform 1 0 23460 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_260
timestamp 1667941163
transform 1 0 25024 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_269
timestamp 1667941163
transform 1 0 25852 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_276
timestamp 1667941163
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_286
timestamp 1667941163
transform 1 0 27416 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_293
timestamp 1667941163
transform 1 0 28060 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_299
timestamp 1667941163
transform 1 0 28612 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_308
timestamp 1667941163
transform 1 0 29440 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_315
timestamp 1667941163
transform 1 0 30084 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_327
timestamp 1667941163
transform 1 0 31188 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_331
timestamp 1667941163
transform 1 0 31556 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1667941163
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1667941163
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1667941163
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1667941163
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_8
timestamp 1667941163
transform 1 0 1840 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_14
timestamp 1667941163
transform 1 0 2392 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_23
timestamp 1667941163
transform 1 0 3220 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1667941163
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_34
timestamp 1667941163
transform 1 0 4232 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_40
timestamp 1667941163
transform 1 0 4784 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_44
timestamp 1667941163
transform 1 0 5152 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_51
timestamp 1667941163
transform 1 0 5796 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_58
timestamp 1667941163
transform 1 0 6440 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_65
timestamp 1667941163
transform 1 0 7084 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1667941163
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_98
timestamp 1667941163
transform 1 0 10120 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_106
timestamp 1667941163
transform 1 0 10856 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_128
timestamp 1667941163
transform 1 0 12880 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1667941163
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_149
timestamp 1667941163
transform 1 0 14812 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_153
timestamp 1667941163
transform 1 0 15180 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_157
timestamp 1667941163
transform 1 0 15548 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_174
timestamp 1667941163
transform 1 0 17112 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_182
timestamp 1667941163
transform 1 0 17848 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_187
timestamp 1667941163
transform 1 0 18308 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1667941163
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_206
timestamp 1667941163
transform 1 0 20056 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_213
timestamp 1667941163
transform 1 0 20700 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_219
timestamp 1667941163
transform 1 0 21252 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_229
timestamp 1667941163
transform 1 0 22172 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_242
timestamp 1667941163
transform 1 0 23368 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_249
timestamp 1667941163
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_258
timestamp 1667941163
transform 1 0 24840 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_279
timestamp 1667941163
transform 1 0 26772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_296
timestamp 1667941163
transform 1 0 28336 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_303
timestamp 1667941163
transform 1 0 28980 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1667941163
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_314
timestamp 1667941163
transform 1 0 29992 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_326
timestamp 1667941163
transform 1 0 31096 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_338
timestamp 1667941163
transform 1 0 32200 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_350
timestamp 1667941163
transform 1 0 33304 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_362
timestamp 1667941163
transform 1 0 34408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_370
timestamp 1667941163
transform 1 0 35144 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_382
timestamp 1667941163
transform 1 0 36248 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_394
timestamp 1667941163
transform 1 0 37352 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_406
timestamp 1667941163
transform 1 0 38456 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_10
timestamp 1667941163
transform 1 0 2024 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_22
timestamp 1667941163
transform 1 0 3128 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_33
timestamp 1667941163
transform 1 0 4140 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_40
timestamp 1667941163
transform 1 0 4784 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_47
timestamp 1667941163
transform 1 0 5428 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1667941163
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_65
timestamp 1667941163
transform 1 0 7084 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_73
timestamp 1667941163
transform 1 0 7820 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_78
timestamp 1667941163
transform 1 0 8280 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_95
timestamp 1667941163
transform 1 0 9844 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1667941163
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_128
timestamp 1667941163
transform 1 0 12880 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_145
timestamp 1667941163
transform 1 0 14444 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_158
timestamp 1667941163
transform 1 0 15640 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_162
timestamp 1667941163
transform 1 0 16008 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1667941163
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_190
timestamp 1667941163
transform 1 0 18584 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_197
timestamp 1667941163
transform 1 0 19228 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_214
timestamp 1667941163
transform 1 0 20792 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1667941163
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_240
timestamp 1667941163
transform 1 0 23184 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_252
timestamp 1667941163
transform 1 0 24288 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_267
timestamp 1667941163
transform 1 0 25668 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_274
timestamp 1667941163
transform 1 0 26312 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_291
timestamp 1667941163
transform 1 0 27876 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_305
timestamp 1667941163
transform 1 0 29164 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_312
timestamp 1667941163
transform 1 0 29808 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_324
timestamp 1667941163
transform 1 0 30912 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_328
timestamp 1667941163
transform 1 0 31280 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_345
timestamp 1667941163
transform 1 0 32844 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1667941163
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1667941163
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1667941163
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1667941163
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1667941163
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_10
timestamp 1667941163
transform 1 0 2024 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_17
timestamp 1667941163
transform 1 0 2668 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_25
timestamp 1667941163
transform 1 0 3404 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_40
timestamp 1667941163
transform 1 0 4784 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_47
timestamp 1667941163
transform 1 0 5428 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_54
timestamp 1667941163
transform 1 0 6072 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_61
timestamp 1667941163
transform 1 0 6716 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_68
timestamp 1667941163
transform 1 0 7360 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_75
timestamp 1667941163
transform 1 0 8004 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1667941163
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_100
timestamp 1667941163
transform 1 0 10304 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_104
timestamp 1667941163
transform 1 0 10672 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_118
timestamp 1667941163
transform 1 0 11960 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_124
timestamp 1667941163
transform 1 0 12512 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1667941163
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_158
timestamp 1667941163
transform 1 0 15640 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_162
timestamp 1667941163
transform 1 0 16008 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_174
timestamp 1667941163
transform 1 0 17112 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_186
timestamp 1667941163
transform 1 0 18216 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_190
timestamp 1667941163
transform 1 0 18584 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1667941163
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_201
timestamp 1667941163
transform 1 0 19596 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_205
timestamp 1667941163
transform 1 0 19964 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_222
timestamp 1667941163
transform 1 0 21528 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_229
timestamp 1667941163
transform 1 0 22172 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_236
timestamp 1667941163
transform 1 0 22816 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_244
timestamp 1667941163
transform 1 0 23552 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1667941163
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_263
timestamp 1667941163
transform 1 0 25300 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_270
timestamp 1667941163
transform 1 0 25944 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_277
timestamp 1667941163
transform 1 0 26588 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_293
timestamp 1667941163
transform 1 0 28060 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_300
timestamp 1667941163
transform 1 0 28704 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_314
timestamp 1667941163
transform 1 0 29992 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_326
timestamp 1667941163
transform 1 0 31096 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_338
timestamp 1667941163
transform 1 0 32200 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_350
timestamp 1667941163
transform 1 0 33304 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_362
timestamp 1667941163
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1667941163
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_405
timestamp 1667941163
transform 1 0 38364 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_9
timestamp 1667941163
transform 1 0 1932 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_16
timestamp 1667941163
transform 1 0 2576 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_28
timestamp 1667941163
transform 1 0 3680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_33
timestamp 1667941163
transform 1 0 4140 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_41
timestamp 1667941163
transform 1 0 4876 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_46
timestamp 1667941163
transform 1 0 5336 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_50
timestamp 1667941163
transform 1 0 5704 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1667941163
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_68
timestamp 1667941163
transform 1 0 7360 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_75
timestamp 1667941163
transform 1 0 8004 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_88
timestamp 1667941163
transform 1 0 9200 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1667941163
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1667941163
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_128
timestamp 1667941163
transform 1 0 12880 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_145
timestamp 1667941163
transform 1 0 14444 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_152
timestamp 1667941163
transform 1 0 15088 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_165
timestamp 1667941163
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_176
timestamp 1667941163
transform 1 0 17296 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_183
timestamp 1667941163
transform 1 0 17940 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_200
timestamp 1667941163
transform 1 0 19504 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_213
timestamp 1667941163
transform 1 0 20700 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_220
timestamp 1667941163
transform 1 0 21344 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_230
timestamp 1667941163
transform 1 0 22264 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_243
timestamp 1667941163
transform 1 0 23460 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_255
timestamp 1667941163
transform 1 0 24564 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_259
timestamp 1667941163
transform 1 0 24932 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_268
timestamp 1667941163
transform 1 0 25760 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_295
timestamp 1667941163
transform 1 0 28244 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_302
timestamp 1667941163
transform 1 0 28888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_309
timestamp 1667941163
transform 1 0 29532 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_318
timestamp 1667941163
transform 1 0 30360 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_325
timestamp 1667941163
transform 1 0 31004 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_333
timestamp 1667941163
transform 1 0 31740 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1667941163
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1667941163
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1667941163
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1667941163
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1667941163
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1667941163
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1667941163
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1667941163
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_53
timestamp 1667941163
transform 1 0 5980 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_59
timestamp 1667941163
transform 1 0 6532 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_76
timestamp 1667941163
transform 1 0 8096 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_94
timestamp 1667941163
transform 1 0 9752 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_107
timestamp 1667941163
transform 1 0 10948 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_120
timestamp 1667941163
transform 1 0 12144 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_137
timestamp 1667941163
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_152
timestamp 1667941163
transform 1 0 15088 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_162
timestamp 1667941163
transform 1 0 16008 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_170
timestamp 1667941163
transform 1 0 16744 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_175
timestamp 1667941163
transform 1 0 17204 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_182
timestamp 1667941163
transform 1 0 17848 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_188
timestamp 1667941163
transform 1 0 18400 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1667941163
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_208
timestamp 1667941163
transform 1 0 20240 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_220
timestamp 1667941163
transform 1 0 21344 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_227
timestamp 1667941163
transform 1 0 21988 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_231
timestamp 1667941163
transform 1 0 22356 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_235
timestamp 1667941163
transform 1 0 22724 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_241
timestamp 1667941163
transform 1 0 23276 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1667941163
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1667941163
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_258
timestamp 1667941163
transform 1 0 24840 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_270
timestamp 1667941163
transform 1 0 25944 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_282
timestamp 1667941163
transform 1 0 27048 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_288
timestamp 1667941163
transform 1 0 27600 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_305
timestamp 1667941163
transform 1 0 29164 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_320
timestamp 1667941163
transform 1 0 30544 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_332
timestamp 1667941163
transform 1 0 31648 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_344
timestamp 1667941163
transform 1 0 32752 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_356
timestamp 1667941163
transform 1 0 33856 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1667941163
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_401
timestamp 1667941163
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_8
timestamp 1667941163
transform 1 0 1840 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_20
timestamp 1667941163
transform 1 0 2944 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_45
timestamp 1667941163
transform 1 0 5244 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_53
timestamp 1667941163
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_62
timestamp 1667941163
transform 1 0 6808 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_69
timestamp 1667941163
transform 1 0 7452 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_76
timestamp 1667941163
transform 1 0 8096 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_83
timestamp 1667941163
transform 1 0 8740 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_90
timestamp 1667941163
transform 1 0 9384 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_97
timestamp 1667941163
transform 1 0 10028 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1667941163
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_123
timestamp 1667941163
transform 1 0 12420 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_142
timestamp 1667941163
transform 1 0 14168 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_150
timestamp 1667941163
transform 1 0 14904 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_155
timestamp 1667941163
transform 1 0 15364 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1667941163
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_185
timestamp 1667941163
transform 1 0 18124 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_191
timestamp 1667941163
transform 1 0 18676 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_201
timestamp 1667941163
transform 1 0 19596 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_208
timestamp 1667941163
transform 1 0 20240 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_212
timestamp 1667941163
transform 1 0 20608 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1667941163
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_241
timestamp 1667941163
transform 1 0 23276 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_258
timestamp 1667941163
transform 1 0 24840 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_270
timestamp 1667941163
transform 1 0 25944 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1667941163
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_293
timestamp 1667941163
transform 1 0 28060 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_302
timestamp 1667941163
transform 1 0 28888 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_309
timestamp 1667941163
transform 1 0 29532 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_321
timestamp 1667941163
transform 1 0 30636 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_333
timestamp 1667941163
transform 1 0 31740 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_343
timestamp 1667941163
transform 1 0 32660 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_347
timestamp 1667941163
transform 1 0 33028 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_359
timestamp 1667941163
transform 1 0 34132 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_371
timestamp 1667941163
transform 1 0 35236 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_383
timestamp 1667941163
transform 1 0 36340 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1667941163
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1667941163
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1667941163
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1667941163
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_33
timestamp 1667941163
transform 1 0 4140 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_37
timestamp 1667941163
transform 1 0 4508 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_44
timestamp 1667941163
transform 1 0 5152 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_56
timestamp 1667941163
transform 1 0 6256 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_68
timestamp 1667941163
transform 1 0 7360 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_75
timestamp 1667941163
transform 1 0 8004 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1667941163
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_92
timestamp 1667941163
transform 1 0 9568 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_99
timestamp 1667941163
transform 1 0 10212 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_106
timestamp 1667941163
transform 1 0 10856 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_123
timestamp 1667941163
transform 1 0 12420 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1667941163
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1667941163
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_148
timestamp 1667941163
transform 1 0 14720 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_161
timestamp 1667941163
transform 1 0 15916 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_178
timestamp 1667941163
transform 1 0 17480 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_190
timestamp 1667941163
transform 1 0 18584 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_202
timestamp 1667941163
transform 1 0 19688 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_209
timestamp 1667941163
transform 1 0 20332 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_217
timestamp 1667941163
transform 1 0 21068 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_221
timestamp 1667941163
transform 1 0 21436 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_228
timestamp 1667941163
transform 1 0 22080 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_235
timestamp 1667941163
transform 1 0 22724 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_247
timestamp 1667941163
transform 1 0 23828 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1667941163
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_265
timestamp 1667941163
transform 1 0 25484 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_281
timestamp 1667941163
transform 1 0 26956 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_289
timestamp 1667941163
transform 1 0 27692 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_294
timestamp 1667941163
transform 1 0 28152 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1667941163
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1667941163
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1667941163
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1667941163
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1667941163
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1667941163
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1667941163
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1667941163
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1667941163
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1667941163
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_27
timestamp 1667941163
transform 1 0 3588 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_31
timestamp 1667941163
transform 1 0 3956 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_41
timestamp 1667941163
transform 1 0 4876 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1667941163
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_61
timestamp 1667941163
transform 1 0 6716 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_75
timestamp 1667941163
transform 1 0 8004 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_82
timestamp 1667941163
transform 1 0 8648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_89
timestamp 1667941163
transform 1 0 9292 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_96
timestamp 1667941163
transform 1 0 9936 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_103
timestamp 1667941163
transform 1 0 10580 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1667941163
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_128
timestamp 1667941163
transform 1 0 12880 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_137
timestamp 1667941163
transform 1 0 13708 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_144
timestamp 1667941163
transform 1 0 14352 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1667941163
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1667941163
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_180
timestamp 1667941163
transform 1 0 17664 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_187
timestamp 1667941163
transform 1 0 18308 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_194
timestamp 1667941163
transform 1 0 18952 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_202
timestamp 1667941163
transform 1 0 19688 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_210
timestamp 1667941163
transform 1 0 20424 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_214
timestamp 1667941163
transform 1 0 20792 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1667941163
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1667941163
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_249
timestamp 1667941163
transform 1 0 24012 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_259
timestamp 1667941163
transform 1 0 24932 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_271
timestamp 1667941163
transform 1 0 26036 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1667941163
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_298
timestamp 1667941163
transform 1 0 28520 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_305
timestamp 1667941163
transform 1 0 29164 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_312
timestamp 1667941163
transform 1 0 29808 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_319
timestamp 1667941163
transform 1 0 30452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_331
timestamp 1667941163
transform 1 0 31556 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1667941163
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1667941163
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1667941163
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1667941163
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1667941163
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1667941163
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_8
timestamp 1667941163
transform 1 0 1840 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_20
timestamp 1667941163
transform 1 0 2944 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_41
timestamp 1667941163
transform 1 0 4876 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_49
timestamp 1667941163
transform 1 0 5612 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_54
timestamp 1667941163
transform 1 0 6072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_61
timestamp 1667941163
transform 1 0 6716 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_68
timestamp 1667941163
transform 1 0 7360 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_75
timestamp 1667941163
transform 1 0 8004 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1667941163
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_90
timestamp 1667941163
transform 1 0 9384 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_97
timestamp 1667941163
transform 1 0 10028 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_104
timestamp 1667941163
transform 1 0 10672 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_111
timestamp 1667941163
transform 1 0 11316 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_118
timestamp 1667941163
transform 1 0 11960 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_135
timestamp 1667941163
transform 1 0 13524 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1667941163
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_156
timestamp 1667941163
transform 1 0 15456 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_160
timestamp 1667941163
transform 1 0 15824 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_170
timestamp 1667941163
transform 1 0 16744 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_177
timestamp 1667941163
transform 1 0 17388 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_184
timestamp 1667941163
transform 1 0 18032 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_209
timestamp 1667941163
transform 1 0 20332 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_214
timestamp 1667941163
transform 1 0 20792 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_226
timestamp 1667941163
transform 1 0 21896 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_238
timestamp 1667941163
transform 1 0 23000 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_246
timestamp 1667941163
transform 1 0 23736 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1667941163
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_268
timestamp 1667941163
transform 1 0 25760 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_281
timestamp 1667941163
transform 1 0 26956 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_288
timestamp 1667941163
transform 1 0 27600 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_300
timestamp 1667941163
transform 1 0 28704 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1667941163
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_319
timestamp 1667941163
transform 1 0 30452 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_327
timestamp 1667941163
transform 1 0 31188 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1667941163
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_345
timestamp 1667941163
transform 1 0 32844 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_351
timestamp 1667941163
transform 1 0 33396 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_355
timestamp 1667941163
transform 1 0 33764 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1667941163
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_371
timestamp 1667941163
transform 1 0 35236 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_383
timestamp 1667941163
transform 1 0 36340 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_395
timestamp 1667941163
transform 1 0 37444 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_10
timestamp 1667941163
transform 1 0 2024 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_22
timestamp 1667941163
transform 1 0 3128 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_34
timestamp 1667941163
transform 1 0 4232 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_45
timestamp 1667941163
transform 1 0 5244 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1667941163
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_69
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_90
timestamp 1667941163
transform 1 0 9384 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_98
timestamp 1667941163
transform 1 0 10120 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_103
timestamp 1667941163
transform 1 0 10580 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1667941163
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_124
timestamp 1667941163
transform 1 0 12512 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_141
timestamp 1667941163
transform 1 0 14076 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_145
timestamp 1667941163
transform 1 0 14444 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_149
timestamp 1667941163
transform 1 0 14812 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_156
timestamp 1667941163
transform 1 0 15456 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_160
timestamp 1667941163
transform 1 0 15824 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1667941163
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_178
timestamp 1667941163
transform 1 0 17480 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_185
timestamp 1667941163
transform 1 0 18124 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_197
timestamp 1667941163
transform 1 0 19228 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_209
timestamp 1667941163
transform 1 0 20332 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_217
timestamp 1667941163
transform 1 0 21068 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1667941163
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_237
timestamp 1667941163
transform 1 0 22908 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_241
timestamp 1667941163
transform 1 0 23276 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_248
timestamp 1667941163
transform 1 0 23920 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_254
timestamp 1667941163
transform 1 0 24472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_258
timestamp 1667941163
transform 1 0 24840 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_265
timestamp 1667941163
transform 1 0 25484 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_277
timestamp 1667941163
transform 1 0 26588 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_286
timestamp 1667941163
transform 1 0 27416 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_298
timestamp 1667941163
transform 1 0 28520 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_302
timestamp 1667941163
transform 1 0 28888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_309
timestamp 1667941163
transform 1 0 29532 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_316
timestamp 1667941163
transform 1 0 30176 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_328
timestamp 1667941163
transform 1 0 31280 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1667941163
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1667941163
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1667941163
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1667941163
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1667941163
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1667941163
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1667941163
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1667941163
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_46
timestamp 1667941163
transform 1 0 5336 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_54
timestamp 1667941163
transform 1 0 6072 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_65
timestamp 1667941163
transform 1 0 7084 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1667941163
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_90
timestamp 1667941163
transform 1 0 9384 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_97
timestamp 1667941163
transform 1 0 10028 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_103
timestamp 1667941163
transform 1 0 10580 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_107
timestamp 1667941163
transform 1 0 10948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_116
timestamp 1667941163
transform 1 0 11776 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_135
timestamp 1667941163
transform 1 0 13524 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1667941163
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_156
timestamp 1667941163
transform 1 0 15456 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_167
timestamp 1667941163
transform 1 0 16468 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_174
timestamp 1667941163
transform 1 0 17112 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_191
timestamp 1667941163
transform 1 0 18676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1667941163
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_206
timestamp 1667941163
transform 1 0 20056 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_231
timestamp 1667941163
transform 1 0 22356 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_239
timestamp 1667941163
transform 1 0 23092 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1667941163
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1667941163
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_263
timestamp 1667941163
transform 1 0 25300 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_270
timestamp 1667941163
transform 1 0 25944 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_277
timestamp 1667941163
transform 1 0 26588 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_284
timestamp 1667941163
transform 1 0 27232 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_296
timestamp 1667941163
transform 1 0 28336 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_314
timestamp 1667941163
transform 1 0 29992 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_326
timestamp 1667941163
transform 1 0 31096 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_338
timestamp 1667941163
transform 1 0 32200 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_350
timestamp 1667941163
transform 1 0 33304 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_362
timestamp 1667941163
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1667941163
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_401
timestamp 1667941163
transform 1 0 37996 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1667941163
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1667941163
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1667941163
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1667941163
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1667941163
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_69
timestamp 1667941163
transform 1 0 7452 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_74
timestamp 1667941163
transform 1 0 7912 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_91
timestamp 1667941163
transform 1 0 9476 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_108
timestamp 1667941163
transform 1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_124
timestamp 1667941163
transform 1 0 12512 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_139
timestamp 1667941163
transform 1 0 13892 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_146
timestamp 1667941163
transform 1 0 14536 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_152
timestamp 1667941163
transform 1 0 15088 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1667941163
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_173
timestamp 1667941163
transform 1 0 17020 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_183
timestamp 1667941163
transform 1 0 17940 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_190
timestamp 1667941163
transform 1 0 18584 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_196
timestamp 1667941163
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_210
timestamp 1667941163
transform 1 0 20424 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1667941163
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_236
timestamp 1667941163
transform 1 0 22816 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_249
timestamp 1667941163
transform 1 0 24012 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_261
timestamp 1667941163
transform 1 0 25116 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_267
timestamp 1667941163
transform 1 0 25668 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_276
timestamp 1667941163
transform 1 0 26496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_286
timestamp 1667941163
transform 1 0 27416 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_298
timestamp 1667941163
transform 1 0 28520 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_310
timestamp 1667941163
transform 1 0 29624 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_322
timestamp 1667941163
transform 1 0 30728 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_334
timestamp 1667941163
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1667941163
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1667941163
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1667941163
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1667941163
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_401
timestamp 1667941163
transform 1 0 37996 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1667941163
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1667941163
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1667941163
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_35
timestamp 1667941163
transform 1 0 4324 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_45
timestamp 1667941163
transform 1 0 5244 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_52
timestamp 1667941163
transform 1 0 5888 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_59
timestamp 1667941163
transform 1 0 6532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_71
timestamp 1667941163
transform 1 0 7636 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1667941163
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_90
timestamp 1667941163
transform 1 0 9384 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_96
timestamp 1667941163
transform 1 0 9936 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_106
timestamp 1667941163
transform 1 0 10856 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_118
timestamp 1667941163
transform 1 0 11960 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1667941163
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1667941163
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_145
timestamp 1667941163
transform 1 0 14444 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_159
timestamp 1667941163
transform 1 0 15732 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_176
timestamp 1667941163
transform 1 0 17296 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_184
timestamp 1667941163
transform 1 0 18032 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1667941163
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_204
timestamp 1667941163
transform 1 0 19872 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_217
timestamp 1667941163
transform 1 0 21068 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_229
timestamp 1667941163
transform 1 0 22172 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_235
timestamp 1667941163
transform 1 0 22724 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_248
timestamp 1667941163
transform 1 0 23920 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_259
timestamp 1667941163
transform 1 0 24932 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_263
timestamp 1667941163
transform 1 0 25300 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_275
timestamp 1667941163
transform 1 0 26404 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_287
timestamp 1667941163
transform 1 0 27508 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_299
timestamp 1667941163
transform 1 0 28612 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1667941163
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1667941163
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1667941163
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1667941163
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1667941163
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1667941163
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_389
timestamp 1667941163
transform 1 0 36892 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_397
timestamp 1667941163
transform 1 0 37628 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_402
timestamp 1667941163
transform 1 0 38088 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_406
timestamp 1667941163
transform 1 0 38456 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_9
timestamp 1667941163
transform 1 0 1932 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_21
timestamp 1667941163
transform 1 0 3036 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_33
timestamp 1667941163
transform 1 0 4140 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1667941163
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_65
timestamp 1667941163
transform 1 0 7084 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_76
timestamp 1667941163
transform 1 0 8096 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_83
timestamp 1667941163
transform 1 0 8740 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_90
timestamp 1667941163
transform 1 0 9384 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_102
timestamp 1667941163
transform 1 0 10488 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1667941163
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_134
timestamp 1667941163
transform 1 0 13432 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_140
timestamp 1667941163
transform 1 0 13984 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_144
timestamp 1667941163
transform 1 0 14352 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_152
timestamp 1667941163
transform 1 0 15088 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1667941163
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_175
timestamp 1667941163
transform 1 0 17204 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_182
timestamp 1667941163
transform 1 0 17848 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_195
timestamp 1667941163
transform 1 0 19044 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_208
timestamp 1667941163
transform 1 0 20240 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_215
timestamp 1667941163
transform 1 0 20884 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1667941163
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_234
timestamp 1667941163
transform 1 0 22632 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_251
timestamp 1667941163
transform 1 0 24196 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_258
timestamp 1667941163
transform 1 0 24840 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_270
timestamp 1667941163
transform 1 0 25944 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1667941163
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_297
timestamp 1667941163
transform 1 0 28428 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_309
timestamp 1667941163
transform 1 0 29532 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_321
timestamp 1667941163
transform 1 0 30636 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_333
timestamp 1667941163
transform 1 0 31740 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1667941163
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1667941163
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1667941163
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1667941163
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1667941163
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1667941163
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1667941163
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_53
timestamp 1667941163
transform 1 0 5980 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_61
timestamp 1667941163
transform 1 0 6716 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_66
timestamp 1667941163
transform 1 0 7176 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_74
timestamp 1667941163
transform 1 0 7912 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_78
timestamp 1667941163
transform 1 0 8280 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_90
timestamp 1667941163
transform 1 0 9384 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_36_105
timestamp 1667941163
transform 1 0 10764 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_120
timestamp 1667941163
transform 1 0 12144 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_132
timestamp 1667941163
transform 1 0 13248 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_146
timestamp 1667941163
transform 1 0 14536 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_156
timestamp 1667941163
transform 1 0 15456 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_163
timestamp 1667941163
transform 1 0 16100 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_174
timestamp 1667941163
transform 1 0 17112 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_187
timestamp 1667941163
transform 1 0 18308 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1667941163
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_203
timestamp 1667941163
transform 1 0 19780 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_215
timestamp 1667941163
transform 1 0 20884 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_227
timestamp 1667941163
transform 1 0 21988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_239
timestamp 1667941163
transform 1 0 23092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1667941163
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_258
timestamp 1667941163
transform 1 0 24840 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_270
timestamp 1667941163
transform 1 0 25944 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_276
timestamp 1667941163
transform 1 0 26496 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1667941163
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1667941163
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1667941163
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1667941163
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1667941163
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1667941163
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1667941163
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1667941163
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_370
timestamp 1667941163
transform 1 0 35144 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_382
timestamp 1667941163
transform 1 0 36248 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_397
timestamp 1667941163
transform 1 0 37628 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_405
timestamp 1667941163
transform 1 0 38364 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_8
timestamp 1667941163
transform 1 0 1840 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_20
timestamp 1667941163
transform 1 0 2944 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_32
timestamp 1667941163
transform 1 0 4048 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_44
timestamp 1667941163
transform 1 0 5152 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_74
timestamp 1667941163
transform 1 0 7912 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_89
timestamp 1667941163
transform 1 0 9292 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_102
timestamp 1667941163
transform 1 0 10488 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_109
timestamp 1667941163
transform 1 0 11132 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_119
timestamp 1667941163
transform 1 0 12052 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_131
timestamp 1667941163
transform 1 0 13156 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_141
timestamp 1667941163
transform 1 0 14076 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_145
timestamp 1667941163
transform 1 0 14444 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_154
timestamp 1667941163
transform 1 0 15272 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_162
timestamp 1667941163
transform 1 0 16008 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1667941163
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_186
timestamp 1667941163
transform 1 0 18216 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1667941163
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_205
timestamp 1667941163
transform 1 0 19964 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_212
timestamp 1667941163
transform 1 0 20608 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_230
timestamp 1667941163
transform 1 0 22264 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_242
timestamp 1667941163
transform 1 0 23368 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_254
timestamp 1667941163
transform 1 0 24472 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_258
timestamp 1667941163
transform 1 0 24840 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_262
timestamp 1667941163
transform 1 0 25208 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_270
timestamp 1667941163
transform 1 0 25944 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_275
timestamp 1667941163
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1667941163
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_292
timestamp 1667941163
transform 1 0 27968 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_304
timestamp 1667941163
transform 1 0 29072 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_316
timestamp 1667941163
transform 1 0 30176 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_320
timestamp 1667941163
transform 1 0 30544 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_325
timestamp 1667941163
transform 1 0 31004 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_333
timestamp 1667941163
transform 1 0 31740 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1667941163
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1667941163
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1667941163
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1667941163
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1667941163
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1667941163
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1667941163
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1667941163
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1667941163
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1667941163
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1667941163
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_94
timestamp 1667941163
transform 1 0 9752 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_111
timestamp 1667941163
transform 1 0 11316 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_119
timestamp 1667941163
transform 1 0 12052 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_124
timestamp 1667941163
transform 1 0 12512 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1667941163
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_156
timestamp 1667941163
transform 1 0 15456 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_163
timestamp 1667941163
transform 1 0 16100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_169
timestamp 1667941163
transform 1 0 16652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_178
timestamp 1667941163
transform 1 0 17480 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_185
timestamp 1667941163
transform 1 0 18124 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_193
timestamp 1667941163
transform 1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_212
timestamp 1667941163
transform 1 0 20608 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_229
timestamp 1667941163
transform 1 0 22172 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_241
timestamp 1667941163
transform 1 0 23276 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_249
timestamp 1667941163
transform 1 0 24012 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1667941163
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1667941163
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1667941163
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1667941163
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1667941163
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1667941163
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1667941163
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1667941163
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1667941163
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1667941163
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1667941163
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1667941163
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 1667941163
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_12
timestamp 1667941163
transform 1 0 2208 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_24
timestamp 1667941163
transform 1 0 3312 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_36
timestamp 1667941163
transform 1 0 4416 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_40
timestamp 1667941163
transform 1 0 4784 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_52
timestamp 1667941163
transform 1 0 5888 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1667941163
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1667941163
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_93
timestamp 1667941163
transform 1 0 9660 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_97
timestamp 1667941163
transform 1 0 10028 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_101
timestamp 1667941163
transform 1 0 10396 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_109
timestamp 1667941163
transform 1 0 11132 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_120
timestamp 1667941163
transform 1 0 12144 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_126
timestamp 1667941163
transform 1 0 12696 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_136
timestamp 1667941163
transform 1 0 13616 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_144
timestamp 1667941163
transform 1 0 14352 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_149
timestamp 1667941163
transform 1 0 14812 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1667941163
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_174
timestamp 1667941163
transform 1 0 17112 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_180
timestamp 1667941163
transform 1 0 17664 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_184
timestamp 1667941163
transform 1 0 18032 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_198
timestamp 1667941163
transform 1 0 19320 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_214
timestamp 1667941163
transform 1 0 20792 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1667941163
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_236
timestamp 1667941163
transform 1 0 22816 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_253
timestamp 1667941163
transform 1 0 24380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_265
timestamp 1667941163
transform 1 0 25484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_277
timestamp 1667941163
transform 1 0 26588 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1667941163
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_305
timestamp 1667941163
transform 1 0 29164 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_314
timestamp 1667941163
transform 1 0 29992 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_321
timestamp 1667941163
transform 1 0 30636 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_333
timestamp 1667941163
transform 1 0 31740 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1667941163
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1667941163
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1667941163
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1667941163
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1667941163
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1667941163
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1667941163
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1667941163
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1667941163
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1667941163
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1667941163
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1667941163
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1667941163
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1667941163
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_121
timestamp 1667941163
transform 1 0 12236 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_132
timestamp 1667941163
transform 1 0 13248 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_152
timestamp 1667941163
transform 1 0 15088 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_160
timestamp 1667941163
transform 1 0 15824 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_168
timestamp 1667941163
transform 1 0 16560 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_173
timestamp 1667941163
transform 1 0 17020 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_181
timestamp 1667941163
transform 1 0 17756 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_40_190
timestamp 1667941163
transform 1 0 18584 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_205
timestamp 1667941163
transform 1 0 19964 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1667941163
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1667941163
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_233
timestamp 1667941163
transform 1 0 22540 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_247
timestamp 1667941163
transform 1 0 23828 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1667941163
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_263
timestamp 1667941163
transform 1 0 25300 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_275
timestamp 1667941163
transform 1 0 26404 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_287
timestamp 1667941163
transform 1 0 27508 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_299
timestamp 1667941163
transform 1 0 28612 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1667941163
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_314
timestamp 1667941163
transform 1 0 29992 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_326
timestamp 1667941163
transform 1 0 31096 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_338
timestamp 1667941163
transform 1 0 32200 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_350
timestamp 1667941163
transform 1 0 33304 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_362
timestamp 1667941163
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1667941163
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_389
timestamp 1667941163
transform 1 0 36892 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_405
timestamp 1667941163
transform 1 0 38364 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_9
timestamp 1667941163
transform 1 0 1932 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_21
timestamp 1667941163
transform 1 0 3036 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_33
timestamp 1667941163
transform 1 0 4140 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_45
timestamp 1667941163
transform 1 0 5244 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_53
timestamp 1667941163
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1667941163
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1667941163
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_93
timestamp 1667941163
transform 1 0 9660 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_101
timestamp 1667941163
transform 1 0 10396 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_106
timestamp 1667941163
transform 1 0 10856 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_118
timestamp 1667941163
transform 1 0 11960 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_125
timestamp 1667941163
transform 1 0 12604 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_142
timestamp 1667941163
transform 1 0 14168 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_159
timestamp 1667941163
transform 1 0 15732 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1667941163
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_178
timestamp 1667941163
transform 1 0 17480 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_195
timestamp 1667941163
transform 1 0 19044 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_202
timestamp 1667941163
transform 1 0 19688 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_214
timestamp 1667941163
transform 1 0 20792 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1667941163
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_230
timestamp 1667941163
transform 1 0 22264 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_234
timestamp 1667941163
transform 1 0 22632 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_244
timestamp 1667941163
transform 1 0 23552 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_250
timestamp 1667941163
transform 1 0 24104 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_254
timestamp 1667941163
transform 1 0 24472 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_261
timestamp 1667941163
transform 1 0 25116 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_267
timestamp 1667941163
transform 1 0 25668 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_271
timestamp 1667941163
transform 1 0 26036 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1667941163
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1667941163
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1667941163
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_317
timestamp 1667941163
transform 1 0 30268 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_324
timestamp 1667941163
transform 1 0 30912 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1667941163
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1667941163
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1667941163
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1667941163
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1667941163
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1667941163
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1667941163
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_53
timestamp 1667941163
transform 1 0 5980 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_59
timestamp 1667941163
transform 1 0 6532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_71
timestamp 1667941163
transform 1 0 7636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1667941163
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_97
timestamp 1667941163
transform 1 0 10028 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_103
timestamp 1667941163
transform 1 0 10580 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_107
timestamp 1667941163
transform 1 0 10948 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_114
timestamp 1667941163
transform 1 0 11592 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_126
timestamp 1667941163
transform 1 0 12696 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1667941163
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_146
timestamp 1667941163
transform 1 0 14536 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_155
timestamp 1667941163
transform 1 0 15364 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_162
timestamp 1667941163
transform 1 0 16008 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_168
timestamp 1667941163
transform 1 0 16560 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_172
timestamp 1667941163
transform 1 0 16928 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_184
timestamp 1667941163
transform 1 0 18032 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_202
timestamp 1667941163
transform 1 0 19688 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_214
timestamp 1667941163
transform 1 0 20792 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_230
timestamp 1667941163
transform 1 0 22264 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_236
timestamp 1667941163
transform 1 0 22816 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_240
timestamp 1667941163
transform 1 0 23184 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_258
timestamp 1667941163
transform 1 0 24840 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_270
timestamp 1667941163
transform 1 0 25944 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_282
timestamp 1667941163
transform 1 0 27048 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_294
timestamp 1667941163
transform 1 0 28152 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_306
timestamp 1667941163
transform 1 0 29256 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_321
timestamp 1667941163
transform 1 0 30636 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_325
timestamp 1667941163
transform 1 0 31004 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_329
timestamp 1667941163
transform 1 0 31372 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_341
timestamp 1667941163
transform 1 0 32476 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_353
timestamp 1667941163
transform 1 0 33580 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_361
timestamp 1667941163
transform 1 0 34316 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1667941163
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_405
timestamp 1667941163
transform 1 0 38364 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1667941163
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1667941163
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1667941163
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1667941163
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1667941163
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_69
timestamp 1667941163
transform 1 0 7452 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_77
timestamp 1667941163
transform 1 0 8188 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1667941163
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_93
timestamp 1667941163
transform 1 0 9660 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_101
timestamp 1667941163
transform 1 0 10396 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1667941163
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1667941163
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_130
timestamp 1667941163
transform 1 0 13064 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_138
timestamp 1667941163
transform 1 0 13800 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_143
timestamp 1667941163
transform 1 0 14260 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_155
timestamp 1667941163
transform 1 0 15364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1667941163
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_181
timestamp 1667941163
transform 1 0 17756 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_200
timestamp 1667941163
transform 1 0 19504 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_210
timestamp 1667941163
transform 1 0 20424 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1667941163
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1667941163
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_235
timestamp 1667941163
transform 1 0 22724 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_247
timestamp 1667941163
transform 1 0 23828 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_259
timestamp 1667941163
transform 1 0 24932 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_271
timestamp 1667941163
transform 1 0 26036 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1667941163
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1667941163
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1667941163
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_317
timestamp 1667941163
transform 1 0 30268 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_321
timestamp 1667941163
transform 1 0 30636 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_333
timestamp 1667941163
transform 1 0 31740 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1667941163
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1667941163
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1667941163
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1667941163
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1667941163
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_9
timestamp 1667941163
transform 1 0 1932 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_21
timestamp 1667941163
transform 1 0 3036 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1667941163
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1667941163
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1667941163
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1667941163
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1667941163
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_92
timestamp 1667941163
transform 1 0 9568 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_96
timestamp 1667941163
transform 1 0 9936 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_100
timestamp 1667941163
transform 1 0 10304 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_107
timestamp 1667941163
transform 1 0 10948 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_114
timestamp 1667941163
transform 1 0 11592 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_126
timestamp 1667941163
transform 1 0 12696 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1667941163
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_150
timestamp 1667941163
transform 1 0 14904 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_162
timestamp 1667941163
transform 1 0 16008 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_169
timestamp 1667941163
transform 1 0 16652 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_181
timestamp 1667941163
transform 1 0 17756 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_193
timestamp 1667941163
transform 1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_209
timestamp 1667941163
transform 1 0 20332 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_215
timestamp 1667941163
transform 1 0 20884 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_222
timestamp 1667941163
transform 1 0 21528 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_230
timestamp 1667941163
transform 1 0 22264 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_235
timestamp 1667941163
transform 1 0 22724 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_242
timestamp 1667941163
transform 1 0 23368 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 1667941163
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1667941163
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1667941163
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1667941163
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1667941163
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1667941163
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1667941163
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1667941163
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1667941163
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1667941163
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1667941163
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1667941163
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1667941163
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_401
timestamp 1667941163
transform 1 0 37996 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_405
timestamp 1667941163
transform 1 0 38364 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1667941163
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1667941163
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1667941163
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1667941163
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1667941163
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1667941163
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1667941163
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_93
timestamp 1667941163
transform 1 0 9660 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_102
timestamp 1667941163
transform 1 0 10488 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1667941163
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_124
timestamp 1667941163
transform 1 0 12512 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_136
timestamp 1667941163
transform 1 0 13616 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_144
timestamp 1667941163
transform 1 0 14352 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_149
timestamp 1667941163
transform 1 0 14812 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_156
timestamp 1667941163
transform 1 0 15456 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1667941163
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1667941163
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1667941163
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1667941163
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1667941163
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_231
timestamp 1667941163
transform 1 0 22356 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_235
timestamp 1667941163
transform 1 0 22724 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_242
timestamp 1667941163
transform 1 0 23368 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_254
timestamp 1667941163
transform 1 0 24472 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_266
timestamp 1667941163
transform 1 0 25576 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_278
timestamp 1667941163
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1667941163
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1667941163
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1667941163
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1667941163
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1667941163
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1667941163
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1667941163
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1667941163
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1667941163
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1667941163
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1667941163
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1667941163
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1667941163
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1667941163
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1667941163
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1667941163
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1667941163
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_97
timestamp 1667941163
transform 1 0 10028 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_104
timestamp 1667941163
transform 1 0 10672 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_111
timestamp 1667941163
transform 1 0 11316 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_123
timestamp 1667941163
transform 1 0 12420 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_135
timestamp 1667941163
transform 1 0 13524 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1667941163
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_147
timestamp 1667941163
transform 1 0 14628 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_151
timestamp 1667941163
transform 1 0 14996 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_163
timestamp 1667941163
transform 1 0 16100 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_175
timestamp 1667941163
transform 1 0 17204 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_187
timestamp 1667941163
transform 1 0 18308 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1667941163
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1667941163
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1667941163
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1667941163
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1667941163
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1667941163
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1667941163
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1667941163
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1667941163
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1667941163
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1667941163
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1667941163
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1667941163
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1667941163
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1667941163
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1667941163
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1667941163
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_401
timestamp 1667941163
transform 1 0 37996 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_405
timestamp 1667941163
transform 1 0 38364 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1667941163
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1667941163
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1667941163
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1667941163
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1667941163
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1667941163
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_81
timestamp 1667941163
transform 1 0 8556 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_90
timestamp 1667941163
transform 1 0 9384 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_98
timestamp 1667941163
transform 1 0 10120 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_103
timestamp 1667941163
transform 1 0 10580 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_110
timestamp 1667941163
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_119
timestamp 1667941163
transform 1 0 12052 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_128
timestamp 1667941163
transform 1 0 12880 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_135
timestamp 1667941163
transform 1 0 13524 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_147
timestamp 1667941163
transform 1 0 14628 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_159
timestamp 1667941163
transform 1 0 15732 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1667941163
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1667941163
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1667941163
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1667941163
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1667941163
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1667941163
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1667941163
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1667941163
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1667941163
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1667941163
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1667941163
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1667941163
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1667941163
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1667941163
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1667941163
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1667941163
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1667941163
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1667941163
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1667941163
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1667941163
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1667941163
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1667941163
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1667941163
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_53
timestamp 1667941163
transform 1 0 5980 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_59
timestamp 1667941163
transform 1 0 6532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_71
timestamp 1667941163
transform 1 0 7636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1667941163
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1667941163
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_109
timestamp 1667941163
transform 1 0 11132 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_116
timestamp 1667941163
transform 1 0 11776 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_128
timestamp 1667941163
transform 1 0 12880 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1667941163
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1667941163
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1667941163
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1667941163
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1667941163
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1667941163
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1667941163
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1667941163
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1667941163
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1667941163
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1667941163
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_277
timestamp 1667941163
transform 1 0 26588 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_285
timestamp 1667941163
transform 1 0 27324 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_290
timestamp 1667941163
transform 1 0 27784 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_302
timestamp 1667941163
transform 1 0 28888 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1667941163
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1667941163
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1667941163
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1667941163
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1667941163
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1667941163
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1667941163
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_8
timestamp 1667941163
transform 1 0 1840 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_20
timestamp 1667941163
transform 1 0 2944 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_32
timestamp 1667941163
transform 1 0 4048 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_44
timestamp 1667941163
transform 1 0 5152 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1667941163
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1667941163
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1667941163
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1667941163
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1667941163
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_117
timestamp 1667941163
transform 1 0 11868 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_121
timestamp 1667941163
transform 1 0 12236 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_133
timestamp 1667941163
transform 1 0 13340 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_145
timestamp 1667941163
transform 1 0 14444 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_157
timestamp 1667941163
transform 1 0 15548 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_165
timestamp 1667941163
transform 1 0 16284 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1667941163
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1667941163
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1667941163
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1667941163
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1667941163
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_230
timestamp 1667941163
transform 1 0 22264 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_242
timestamp 1667941163
transform 1 0 23368 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_254
timestamp 1667941163
transform 1 0 24472 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_266
timestamp 1667941163
transform 1 0 25576 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_278
timestamp 1667941163
transform 1 0 26680 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1667941163
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1667941163
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1667941163
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1667941163
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1667941163
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1667941163
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1667941163
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_401
timestamp 1667941163
transform 1 0 37996 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1667941163
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_9
timestamp 1667941163
transform 1 0 1932 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_21
timestamp 1667941163
transform 1 0 3036 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1667941163
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1667941163
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1667941163
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1667941163
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1667941163
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1667941163
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1667941163
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_109
timestamp 1667941163
transform 1 0 11132 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_115
timestamp 1667941163
transform 1 0 11684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_127
timestamp 1667941163
transform 1 0 12788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1667941163
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1667941163
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1667941163
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1667941163
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1667941163
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1667941163
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1667941163
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_224
timestamp 1667941163
transform 1 0 21712 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_236
timestamp 1667941163
transform 1 0 22816 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_248
timestamp 1667941163
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1667941163
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1667941163
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1667941163
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1667941163
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1667941163
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_314
timestamp 1667941163
transform 1 0 29992 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_326
timestamp 1667941163
transform 1 0 31096 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_338
timestamp 1667941163
transform 1 0 32200 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_350
timestamp 1667941163
transform 1 0 33304 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_362
timestamp 1667941163
transform 1 0 34408 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1667941163
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1667941163
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_405
timestamp 1667941163
transform 1 0 38364 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1667941163
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1667941163
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1667941163
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1667941163
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1667941163
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_62
timestamp 1667941163
transform 1 0 6808 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_74
timestamp 1667941163
transform 1 0 7912 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_86
timestamp 1667941163
transform 1 0 9016 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_98
timestamp 1667941163
transform 1 0 10120 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1667941163
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1667941163
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_137
timestamp 1667941163
transform 1 0 13708 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_141
timestamp 1667941163
transform 1 0 14076 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_148
timestamp 1667941163
transform 1 0 14720 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_160
timestamp 1667941163
transform 1 0 15824 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1667941163
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1667941163
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1667941163
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1667941163
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1667941163
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_237
timestamp 1667941163
transform 1 0 22908 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_241
timestamp 1667941163
transform 1 0 23276 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_245
timestamp 1667941163
transform 1 0 23644 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_257
timestamp 1667941163
transform 1 0 24748 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_269
timestamp 1667941163
transform 1 0 25852 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_276
timestamp 1667941163
transform 1 0 26496 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1667941163
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_305
timestamp 1667941163
transform 1 0 29164 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_312
timestamp 1667941163
transform 1 0 29808 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_324
timestamp 1667941163
transform 1 0 30912 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1667941163
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1667941163
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1667941163
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1667941163
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_402
timestamp 1667941163
transform 1 0 38088 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_406
timestamp 1667941163
transform 1 0 38456 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_9
timestamp 1667941163
transform 1 0 1932 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_21
timestamp 1667941163
transform 1 0 3036 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1667941163
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_34
timestamp 1667941163
transform 1 0 4232 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_46
timestamp 1667941163
transform 1 0 5336 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_58
timestamp 1667941163
transform 1 0 6440 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_70
timestamp 1667941163
transform 1 0 7544 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_82
timestamp 1667941163
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_97
timestamp 1667941163
transform 1 0 10028 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_104
timestamp 1667941163
transform 1 0 10672 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_116
timestamp 1667941163
transform 1 0 11776 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_128
timestamp 1667941163
transform 1 0 12880 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1667941163
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1667941163
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1667941163
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1667941163
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1667941163
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1667941163
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_221
timestamp 1667941163
transform 1 0 21436 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_228
timestamp 1667941163
transform 1 0 22080 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_237
timestamp 1667941163
transform 1 0 22908 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_249
timestamp 1667941163
transform 1 0 24012 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1667941163
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1667941163
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_289
timestamp 1667941163
transform 1 0 27692 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_295
timestamp 1667941163
transform 1 0 28244 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1667941163
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1667941163
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1667941163
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1667941163
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1667941163
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1667941163
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_377
timestamp 1667941163
transform 1 0 35788 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_384
timestamp 1667941163
transform 1 0 36432 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_396
timestamp 1667941163
transform 1 0 37536 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_52_405
timestamp 1667941163
transform 1 0 38364 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1667941163
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1667941163
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1667941163
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1667941163
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1667941163
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_62
timestamp 1667941163
transform 1 0 6808 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1667941163
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1667941163
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1667941163
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1667941163
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1667941163
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1667941163
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1667941163
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1667941163
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1667941163
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1667941163
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_174
timestamp 1667941163
transform 1 0 17112 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_186
timestamp 1667941163
transform 1 0 18216 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_198
timestamp 1667941163
transform 1 0 19320 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_210
timestamp 1667941163
transform 1 0 20424 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1667941163
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1667941163
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1667941163
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1667941163
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1667941163
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1667941163
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1667941163
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1667941163
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1667941163
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1667941163
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_344
timestamp 1667941163
transform 1 0 32752 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_356
timestamp 1667941163
transform 1 0 33856 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_368
timestamp 1667941163
transform 1 0 34960 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_380
timestamp 1667941163
transform 1 0 36064 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1667941163
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1667941163
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1667941163
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1667941163
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1667941163
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_65
timestamp 1667941163
transform 1 0 7084 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_73
timestamp 1667941163
transform 1 0 7820 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1667941163
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1667941163
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1667941163
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1667941163
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1667941163
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1667941163
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1667941163
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1667941163
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1667941163
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1667941163
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1667941163
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1667941163
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_221
timestamp 1667941163
transform 1 0 21436 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_229
timestamp 1667941163
transform 1 0 22172 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1667941163
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1667941163
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1667941163
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_265
timestamp 1667941163
transform 1 0 25484 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_270
timestamp 1667941163
transform 1 0 25944 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_282
timestamp 1667941163
transform 1 0 27048 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_288
timestamp 1667941163
transform 1 0 27600 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_295
timestamp 1667941163
transform 1 0 28244 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1667941163
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_328
timestamp 1667941163
transform 1 0 31280 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_340
timestamp 1667941163
transform 1 0 32384 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_352
timestamp 1667941163
transform 1 0 33488 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_392
timestamp 1667941163
transform 1 0 37168 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_404
timestamp 1667941163
transform 1 0 38272 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_9
timestamp 1667941163
transform 1 0 1932 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_21
timestamp 1667941163
transform 1 0 3036 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_33
timestamp 1667941163
transform 1 0 4140 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_45
timestamp 1667941163
transform 1 0 5244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_53
timestamp 1667941163
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1667941163
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1667941163
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1667941163
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1667941163
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1667941163
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1667941163
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1667941163
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1667941163
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1667941163
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1667941163
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1667941163
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1667941163
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1667941163
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1667941163
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1667941163
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1667941163
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1667941163
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1667941163
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1667941163
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1667941163
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1667941163
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_305
timestamp 1667941163
transform 1 0 29164 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_309
timestamp 1667941163
transform 1 0 29532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_313
timestamp 1667941163
transform 1 0 29900 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_325
timestamp 1667941163
transform 1 0 31004 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_333
timestamp 1667941163
transform 1 0 31740 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1667941163
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1667941163
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1667941163
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1667941163
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_401
timestamp 1667941163
transform 1 0 37996 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1667941163
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_9
timestamp 1667941163
transform 1 0 1932 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_16
timestamp 1667941163
transform 1 0 2576 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1667941163
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1667941163
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1667941163
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1667941163
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1667941163
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1667941163
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1667941163
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1667941163
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1667941163
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1667941163
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1667941163
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1667941163
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1667941163
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1667941163
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1667941163
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1667941163
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1667941163
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1667941163
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1667941163
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1667941163
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1667941163
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1667941163
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1667941163
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_333
timestamp 1667941163
transform 1 0 31740 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_340
timestamp 1667941163
transform 1 0 32384 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_352
timestamp 1667941163
transform 1 0 33488 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_389
timestamp 1667941163
transform 1 0 36892 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_405
timestamp 1667941163
transform 1 0 38364 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1667941163
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1667941163
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1667941163
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1667941163
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1667941163
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1667941163
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1667941163
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1667941163
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1667941163
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1667941163
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1667941163
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_149
timestamp 1667941163
transform 1 0 14812 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_57_158
timestamp 1667941163
transform 1 0 15640 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_166
timestamp 1667941163
transform 1 0 16376 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1667941163
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1667941163
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1667941163
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1667941163
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1667941163
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_231
timestamp 1667941163
transform 1 0 22356 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_243
timestamp 1667941163
transform 1 0 23460 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_255
timestamp 1667941163
transform 1 0 24564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_267
timestamp 1667941163
transform 1 0 25668 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1667941163
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1667941163
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1667941163
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1667941163
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1667941163
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1667941163
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1667941163
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1667941163
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1667941163
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1667941163
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1667941163
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1667941163
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1667941163
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1667941163
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1667941163
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1667941163
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1667941163
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1667941163
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1667941163
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1667941163
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1667941163
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1667941163
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1667941163
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1667941163
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1667941163
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1667941163
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1667941163
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1667941163
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1667941163
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1667941163
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1667941163
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1667941163
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1667941163
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1667941163
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1667941163
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1667941163
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1667941163
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1667941163
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 1667941163
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_9
timestamp 1667941163
transform 1 0 1932 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_21
timestamp 1667941163
transform 1 0 3036 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_33
timestamp 1667941163
transform 1 0 4140 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_45
timestamp 1667941163
transform 1 0 5244 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_53
timestamp 1667941163
transform 1 0 5980 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_62
timestamp 1667941163
transform 1 0 6808 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_74
timestamp 1667941163
transform 1 0 7912 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_86
timestamp 1667941163
transform 1 0 9016 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_98
timestamp 1667941163
transform 1 0 10120 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_110
timestamp 1667941163
transform 1 0 11224 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1667941163
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1667941163
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1667941163
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1667941163
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1667941163
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1667941163
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1667941163
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1667941163
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1667941163
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1667941163
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1667941163
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1667941163
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1667941163
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1667941163
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1667941163
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1667941163
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1667941163
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1667941163
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1667941163
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1667941163
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1667941163
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1667941163
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1667941163
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1667941163
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1667941163
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1667941163
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1667941163
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1667941163
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1667941163
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1667941163
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1667941163
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1667941163
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1667941163
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1667941163
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1667941163
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_147
timestamp 1667941163
transform 1 0 14628 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_151
timestamp 1667941163
transform 1 0 14996 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_163
timestamp 1667941163
transform 1 0 16100 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_175
timestamp 1667941163
transform 1 0 17204 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_187
timestamp 1667941163
transform 1 0 18308 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1667941163
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1667941163
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1667941163
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1667941163
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1667941163
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1667941163
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1667941163
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1667941163
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1667941163
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1667941163
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1667941163
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1667941163
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1667941163
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1667941163
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1667941163
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1667941163
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1667941163
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_401
timestamp 1667941163
transform 1 0 37996 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_8
timestamp 1667941163
transform 1 0 1840 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_20
timestamp 1667941163
transform 1 0 2944 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_32
timestamp 1667941163
transform 1 0 4048 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_44
timestamp 1667941163
transform 1 0 5152 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1667941163
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1667941163
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1667941163
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1667941163
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1667941163
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1667941163
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1667941163
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1667941163
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1667941163
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1667941163
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1667941163
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1667941163
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1667941163
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1667941163
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1667941163
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1667941163
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1667941163
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1667941163
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1667941163
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1667941163
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1667941163
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1667941163
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_376
timestamp 1667941163
transform 1 0 35696 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_388
timestamp 1667941163
transform 1 0 36800 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_9
timestamp 1667941163
transform 1 0 1932 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_16
timestamp 1667941163
transform 1 0 2576 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1667941163
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1667941163
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1667941163
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1667941163
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1667941163
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1667941163
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1667941163
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1667941163
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1667941163
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1667941163
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1667941163
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1667941163
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1667941163
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1667941163
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1667941163
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1667941163
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1667941163
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1667941163
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1667941163
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1667941163
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1667941163
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1667941163
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1667941163
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1667941163
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1667941163
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1667941163
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1667941163
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1667941163
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1667941163
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_377
timestamp 1667941163
transform 1 0 35788 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_385
timestamp 1667941163
transform 1 0 36524 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_389
timestamp 1667941163
transform 1 0 36892 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_397
timestamp 1667941163
transform 1 0 37628 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_405
timestamp 1667941163
transform 1 0 38364 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_9
timestamp 1667941163
transform 1 0 1932 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_20
timestamp 1667941163
transform 1 0 2944 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1667941163
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1667941163
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1667941163
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1667941163
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1667941163
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_81
timestamp 1667941163
transform 1 0 8556 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_90
timestamp 1667941163
transform 1 0 9384 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_98
timestamp 1667941163
transform 1 0 10120 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_104
timestamp 1667941163
transform 1 0 10672 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1667941163
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1667941163
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1667941163
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1667941163
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1667941163
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1667941163
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_193
timestamp 1667941163
transform 1 0 18860 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_203
timestamp 1667941163
transform 1 0 19780 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_215
timestamp 1667941163
transform 1 0 20884 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1667941163
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_237
timestamp 1667941163
transform 1 0 22908 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_245
timestamp 1667941163
transform 1 0 23644 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_257
timestamp 1667941163
transform 1 0 24748 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_269
timestamp 1667941163
transform 1 0 25852 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_277
timestamp 1667941163
transform 1 0 26588 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_286
timestamp 1667941163
transform 1 0 27416 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_298
timestamp 1667941163
transform 1 0 28520 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_310
timestamp 1667941163
transform 1 0 29624 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_322
timestamp 1667941163
transform 1 0 30728 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_334
timestamp 1667941163
transform 1 0 31832 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1667941163
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_361
timestamp 1667941163
transform 1 0 34316 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_369
timestamp 1667941163
transform 1 0 35052 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_374
timestamp 1667941163
transform 1 0 35512 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_382
timestamp 1667941163
transform 1 0 36248 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_390
timestamp 1667941163
transform 1 0 36984 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_399
timestamp 1667941163
transform 1 0 37812 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_403
timestamp 1667941163
transform 1 0 38180 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_9
timestamp 1667941163
transform 1 0 1932 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_20
timestamp 1667941163
transform 1 0 2944 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_41
timestamp 1667941163
transform 1 0 4876 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_48
timestamp 1667941163
transform 1 0 5520 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_62
timestamp 1667941163
transform 1 0 6808 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_69
timestamp 1667941163
transform 1 0 7452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_81
timestamp 1667941163
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_97
timestamp 1667941163
transform 1 0 10028 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_105
timestamp 1667941163
transform 1 0 10764 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_111
timestamp 1667941163
transform 1 0 11316 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_118
timestamp 1667941163
transform 1 0 11960 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_126
timestamp 1667941163
transform 1 0 12696 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_138
timestamp 1667941163
transform 1 0 13800 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_147
timestamp 1667941163
transform 1 0 14628 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_154
timestamp 1667941163
transform 1 0 15272 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_166
timestamp 1667941163
transform 1 0 16376 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_175
timestamp 1667941163
transform 1 0 17204 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_183
timestamp 1667941163
transform 1 0 17940 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_188
timestamp 1667941163
transform 1 0 18400 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_205
timestamp 1667941163
transform 1 0 19964 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_210
timestamp 1667941163
transform 1 0 20424 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_222
timestamp 1667941163
transform 1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_233
timestamp 1667941163
transform 1 0 22540 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_244
timestamp 1667941163
transform 1 0 23552 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_258
timestamp 1667941163
transform 1 0 24840 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_266
timestamp 1667941163
transform 1 0 25576 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_272
timestamp 1667941163
transform 1 0 26128 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_287
timestamp 1667941163
transform 1 0 27508 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_294
timestamp 1667941163
transform 1 0 28152 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_306
timestamp 1667941163
transform 1 0 29256 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_314
timestamp 1667941163
transform 1 0 29992 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_321
timestamp 1667941163
transform 1 0 30636 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_329
timestamp 1667941163
transform 1 0 31372 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_335
timestamp 1667941163
transform 1 0 31924 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_342
timestamp 1667941163
transform 1 0 32568 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_350
timestamp 1667941163
transform 1 0 33304 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_362
timestamp 1667941163
transform 1 0 34408 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_371
timestamp 1667941163
transform 1 0 35236 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_379
timestamp 1667941163
transform 1 0 35972 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_385
timestamp 1667941163
transform 1 0 36524 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_391
timestamp 1667941163
transform 1 0 37076 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_393
timestamp 1667941163
transform 1 0 37260 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_405
timestamp 1667941163
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0390_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 28888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0391_
timestamp 1667941163
transform 1 0 28428 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0392_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 30084 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0393_
timestamp 1667941163
transform 1 0 30728 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0394_
timestamp 1667941163
transform 1 0 28612 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0395_
timestamp 1667941163
transform 1 0 29716 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0396_
timestamp 1667941163
transform 1 0 10580 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0397_
timestamp 1667941163
transform 1 0 1748 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0398_
timestamp 1667941163
transform 1 0 1564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0399_
timestamp 1667941163
transform 1 0 1932 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0400_
timestamp 1667941163
transform 1 0 3036 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0401_
timestamp 1667941163
transform 1 0 1748 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0402_
timestamp 1667941163
transform 1 0 2300 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0403_
timestamp 1667941163
transform 1 0 28980 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0404_
timestamp 1667941163
transform 1 0 17204 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0405_
timestamp 1667941163
transform 1 0 22356 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0406_
timestamp 1667941163
transform 1 0 24564 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0407_
timestamp 1667941163
transform 1 0 29532 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0408_
timestamp 1667941163
transform 1 0 29900 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0409_
timestamp 1667941163
transform 1 0 27140 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0410_
timestamp 1667941163
transform 1 0 14444 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0411_
timestamp 1667941163
transform 1 0 17756 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0412_
timestamp 1667941163
transform 1 0 14536 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0413_
timestamp 1667941163
transform 1 0 28612 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0414_
timestamp 1667941163
transform 1 0 29716 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0415_
timestamp 1667941163
transform 1 0 30820 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0416_
timestamp 1667941163
transform 1 0 26312 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0417_
timestamp 1667941163
transform 1 0 26312 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0418_
timestamp 1667941163
transform 1 0 26036 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0419_
timestamp 1667941163
transform 1 0 30728 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0420_
timestamp 1667941163
transform 1 0 31372 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0421_
timestamp 1667941163
transform 1 0 10488 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0422_
timestamp 1667941163
transform 1 0 15732 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0423_
timestamp 1667941163
transform 1 0 13984 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0424_
timestamp 1667941163
transform 1 0 14536 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0425_
timestamp 1667941163
transform 1 0 10028 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0426_
timestamp 1667941163
transform 1 0 10212 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0427_
timestamp 1667941163
transform 1 0 16376 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0428_
timestamp 1667941163
transform 1 0 14628 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0429_
timestamp 1667941163
transform 1 0 15180 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0430_
timestamp 1667941163
transform 1 0 28336 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0431_
timestamp 1667941163
transform 1 0 29256 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0432_
timestamp 1667941163
transform 1 0 17848 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0433_
timestamp 1667941163
transform 1 0 16836 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0434_
timestamp 1667941163
transform 1 0 29716 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0435_
timestamp 1667941163
transform 1 0 29256 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0436_
timestamp 1667941163
transform 1 0 27784 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0437_
timestamp 1667941163
transform 1 0 29532 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0438_
timestamp 1667941163
transform 1 0 29716 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0439_
timestamp 1667941163
transform 1 0 24564 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0440_
timestamp 1667941163
transform 1 0 17756 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0441_
timestamp 1667941163
transform 1 0 22448 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0442_
timestamp 1667941163
transform 1 0 22908 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0443_
timestamp 1667941163
transform 1 0 25668 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0444_
timestamp 1667941163
transform 1 0 25024 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0445_
timestamp 1667941163
transform 1 0 21988 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0446_
timestamp 1667941163
transform 1 0 22448 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0447_
timestamp 1667941163
transform 1 0 23092 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0448_
timestamp 1667941163
transform 1 0 27784 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0449_
timestamp 1667941163
transform 1 0 21252 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0450_
timestamp 1667941163
transform 1 0 23644 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0451_
timestamp 1667941163
transform 1 0 23000 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0452_
timestamp 1667941163
transform 1 0 30452 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0453_
timestamp 1667941163
transform 1 0 29900 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0454_
timestamp 1667941163
transform 1 0 29072 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0455_
timestamp 1667941163
transform 1 0 31004 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0456_
timestamp 1667941163
transform 1 0 31280 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0457_
timestamp 1667941163
transform 1 0 12604 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0458_
timestamp 1667941163
transform 1 0 11776 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0459_
timestamp 1667941163
transform 1 0 10304 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0460_
timestamp 1667941163
transform 1 0 11500 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0461_
timestamp 1667941163
transform 1 0 10396 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0462_
timestamp 1667941163
transform 1 0 10948 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0463_
timestamp 1667941163
transform 1 0 11684 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0464_
timestamp 1667941163
transform 1 0 11316 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0465_
timestamp 1667941163
transform 1 0 13248 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0466_
timestamp 1667941163
transform 1 0 26128 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0467_
timestamp 1667941163
transform 1 0 27140 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0468_
timestamp 1667941163
transform 1 0 27140 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0469_
timestamp 1667941163
transform 1 0 27324 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0470_
timestamp 1667941163
transform 1 0 24196 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0471_
timestamp 1667941163
transform 1 0 24840 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0472_
timestamp 1667941163
transform 1 0 18308 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0473_
timestamp 1667941163
transform 1 0 20608 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0474_
timestamp 1667941163
transform 1 0 21252 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0475_
timestamp 1667941163
transform 1 0 18032 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0476_
timestamp 1667941163
transform 1 0 18124 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0477_
timestamp 1667941163
transform 1 0 14812 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0478_
timestamp 1667941163
transform 1 0 6164 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0479_
timestamp 1667941163
transform 1 0 21804 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0480_
timestamp 1667941163
transform 1 0 18676 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0481_
timestamp 1667941163
transform 1 0 20056 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0482_
timestamp 1667941163
transform 1 0 27140 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0483_
timestamp 1667941163
transform 1 0 32292 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0484_
timestamp 1667941163
transform 1 0 13432 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0485_
timestamp 1667941163
transform 1 0 18492 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0486_
timestamp 1667941163
transform 1 0 21068 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0487_
timestamp 1667941163
transform 1 0 24656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0488_
timestamp 1667941163
transform 1 0 20516 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0489_
timestamp 1667941163
transform 1 0 27784 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0490_
timestamp 1667941163
transform 1 0 22356 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0491_
timestamp 1667941163
transform 1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0492_
timestamp 1667941163
transform 1 0 23736 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0493_
timestamp 1667941163
transform 1 0 33580 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0494_
timestamp 1667941163
transform 1 0 29716 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0495_
timestamp 1667941163
transform 1 0 21068 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0496_
timestamp 1667941163
transform 1 0 25668 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0497_
timestamp 1667941163
transform 1 0 16928 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0498_
timestamp 1667941163
transform 1 0 4232 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0499_
timestamp 1667941163
transform 1 0 14076 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0500_
timestamp 1667941163
transform 1 0 6256 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0501_
timestamp 1667941163
transform 1 0 21712 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0502_
timestamp 1667941163
transform 1 0 18676 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0503_
timestamp 1667941163
transform 1 0 20516 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0504_
timestamp 1667941163
transform 1 0 8004 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0505_
timestamp 1667941163
transform 1 0 11040 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0506_
timestamp 1667941163
transform 1 0 17572 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0507_
timestamp 1667941163
transform 1 0 10856 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0508_
timestamp 1667941163
transform 1 0 16100 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0509_
timestamp 1667941163
transform 1 0 10396 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0510_
timestamp 1667941163
transform 1 0 10672 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0511_
timestamp 1667941163
transform 1 0 10120 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0512_
timestamp 1667941163
transform 1 0 11868 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0513_
timestamp 1667941163
transform 1 0 10304 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0514_
timestamp 1667941163
transform 1 0 8464 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0515_
timestamp 1667941163
transform 1 0 11776 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0516_
timestamp 1667941163
transform 1 0 14536 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0517_
timestamp 1667941163
transform 1 0 29072 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0518_
timestamp 1667941163
transform 1 0 26312 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0519_
timestamp 1667941163
transform 1 0 28704 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0520_
timestamp 1667941163
transform 1 0 8372 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0521_
timestamp 1667941163
transform 1 0 29716 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0522_
timestamp 1667941163
transform 1 0 27968 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0523_
timestamp 1667941163
transform 1 0 23828 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0524_
timestamp 1667941163
transform 1 0 8372 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0525_
timestamp 1667941163
transform 1 0 30360 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0526_
timestamp 1667941163
transform 1 0 28060 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0527_
timestamp 1667941163
transform 1 0 27140 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0528_
timestamp 1667941163
transform 1 0 7084 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0529_
timestamp 1667941163
transform 1 0 9108 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0530_
timestamp 1667941163
transform 1 0 26220 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0531_
timestamp 1667941163
transform 1 0 26956 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0532_
timestamp 1667941163
transform 1 0 9016 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0533_
timestamp 1667941163
transform 1 0 10304 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0534_
timestamp 1667941163
transform 1 0 20608 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0535_
timestamp 1667941163
transform 1 0 19504 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0536_
timestamp 1667941163
transform 1 0 18584 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0537_
timestamp 1667941163
transform 1 0 9660 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0538_
timestamp 1667941163
transform 1 0 24564 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0539_
timestamp 1667941163
transform 1 0 24932 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0540_
timestamp 1667941163
transform 1 0 21988 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0541_
timestamp 1667941163
transform 1 0 9108 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0542_
timestamp 1667941163
transform 1 0 23184 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0543_
timestamp 1667941163
transform 1 0 24564 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0544_
timestamp 1667941163
transform 1 0 9108 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0545_
timestamp 1667941163
transform 1 0 17572 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0546_
timestamp 1667941163
transform 1 0 23368 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0547_
timestamp 1667941163
transform 1 0 9752 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0548_
timestamp 1667941163
transform 1 0 9752 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0549_
timestamp 1667941163
transform 1 0 9752 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0550_
timestamp 1667941163
transform 1 0 19964 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0551_
timestamp 1667941163
transform 1 0 22448 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0552_
timestamp 1667941163
transform 1 0 9752 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0553_
timestamp 1667941163
transform 1 0 30360 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0554_
timestamp 1667941163
transform 1 0 24288 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0555_
timestamp 1667941163
transform 1 0 27416 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0556_
timestamp 1667941163
transform 1 0 14260 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0557_
timestamp 1667941163
transform 1 0 11500 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0558_
timestamp 1667941163
transform 1 0 29716 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0559_
timestamp 1667941163
transform 1 0 24564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0560_
timestamp 1667941163
transform 1 0 24932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0561_
timestamp 1667941163
transform 1 0 7820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0562_
timestamp 1667941163
transform 1 0 25208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0563_
timestamp 1667941163
transform 1 0 16836 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0564_
timestamp 1667941163
transform 1 0 9108 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0565_
timestamp 1667941163
transform 1 0 23000 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0566_
timestamp 1667941163
transform 1 0 18492 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0567_
timestamp 1667941163
transform 1 0 4876 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0568_
timestamp 1667941163
transform 1 0 23828 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0569_
timestamp 1667941163
transform 1 0 25576 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0570_
timestamp 1667941163
transform 1 0 25484 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0571_
timestamp 1667941163
transform 1 0 22448 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0572_
timestamp 1667941163
transform 1 0 19688 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0573_
timestamp 1667941163
transform 1 0 15180 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0574_
timestamp 1667941163
transform 1 0 9936 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0575_
timestamp 1667941163
transform 1 0 19780 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0576_
timestamp 1667941163
transform 1 0 11868 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0577_
timestamp 1667941163
transform 1 0 7728 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0578_
timestamp 1667941163
transform 1 0 5796 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0579_
timestamp 1667941163
transform 1 0 8004 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0580_
timestamp 1667941163
transform 1 0 14260 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0581_
timestamp 1667941163
transform 1 0 12328 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0582_
timestamp 1667941163
transform 1 0 7636 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0583_
timestamp 1667941163
transform 1 0 9292 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0584_
timestamp 1667941163
transform 1 0 8372 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0585_
timestamp 1667941163
transform 1 0 4968 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0586_
timestamp 1667941163
transform 1 0 16192 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0587_
timestamp 1667941163
transform 1 0 17848 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0588_
timestamp 1667941163
transform 1 0 16744 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0589_
timestamp 1667941163
transform 1 0 23552 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0590_
timestamp 1667941163
transform 1 0 30268 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0591_
timestamp 1667941163
transform 1 0 26312 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0592_
timestamp 1667941163
transform 1 0 12236 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0593_
timestamp 1667941163
transform 1 0 28980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0594_
timestamp 1667941163
transform 1 0 26220 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0595_
timestamp 1667941163
transform 1 0 22448 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0596_
timestamp 1667941163
transform 1 0 22264 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0597_
timestamp 1667941163
transform 1 0 2300 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0598_
timestamp 1667941163
transform 1 0 10948 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0599_
timestamp 1667941163
transform 1 0 17112 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0600_
timestamp 1667941163
transform 1 0 17020 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0601_
timestamp 1667941163
transform 1 0 7728 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0602_
timestamp 1667941163
transform 1 0 17204 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0603_
timestamp 1667941163
transform 1 0 10948 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0604_
timestamp 1667941163
transform 1 0 12236 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0605_
timestamp 1667941163
transform 1 0 9108 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0606_
timestamp 1667941163
transform 1 0 7176 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0607_
timestamp 1667941163
transform 1 0 18400 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0608_
timestamp 1667941163
transform 1 0 5152 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0609_
timestamp 1667941163
transform 1 0 16100 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0610_
timestamp 1667941163
transform 1 0 16100 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0611_
timestamp 1667941163
transform 1 0 16836 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0612_
timestamp 1667941163
transform 1 0 8372 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0613_
timestamp 1667941163
transform 1 0 21160 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0614_
timestamp 1667941163
transform 1 0 20424 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0615_
timestamp 1667941163
transform 1 0 21712 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0616_
timestamp 1667941163
transform 1 0 10672 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0617_
timestamp 1667941163
transform 1 0 16652 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0618_
timestamp 1667941163
transform 1 0 20792 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0619_
timestamp 1667941163
transform 1 0 10580 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0620_
timestamp 1667941163
transform 1 0 14260 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0621_
timestamp 1667941163
transform 1 0 19412 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0622_
timestamp 1667941163
transform 1 0 27692 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0623_
timestamp 1667941163
transform 1 0 7728 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0624_
timestamp 1667941163
transform 1 0 37352 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0625_
timestamp 1667941163
transform 1 0 25668 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0626_
timestamp 1667941163
transform 1 0 31648 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0627_
timestamp 1667941163
transform 1 0 3956 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0628_
timestamp 1667941163
transform 1 0 7912 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0629_
timestamp 1667941163
transform 1 0 31096 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0630_
timestamp 1667941163
transform 1 0 36156 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0631_
timestamp 1667941163
transform 1 0 30360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0632_
timestamp 1667941163
transform 1 0 28336 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0633_
timestamp 1667941163
transform 1 0 6900 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0634_
timestamp 1667941163
transform 1 0 22540 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0635_
timestamp 1667941163
transform 1 0 30360 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0636_
timestamp 1667941163
transform 1 0 30360 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0637_
timestamp 1667941163
transform 1 0 3956 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0638_
timestamp 1667941163
transform 1 0 7176 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0639_
timestamp 1667941163
transform 1 0 15824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0640_
timestamp 1667941163
transform 1 0 11040 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0641_
timestamp 1667941163
transform 1 0 5612 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0642_
timestamp 1667941163
transform 1 0 23368 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0643_
timestamp 1667941163
transform 1 0 34868 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0644_
timestamp 1667941163
transform 1 0 11408 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0645_
timestamp 1667941163
transform 1 0 29716 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0646_
timestamp 1667941163
transform 1 0 2300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0647_
timestamp 1667941163
transform 1 0 16836 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0648_
timestamp 1667941163
transform 1 0 3680 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0649_
timestamp 1667941163
transform 1 0 27508 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0650_
timestamp 1667941163
transform 1 0 28704 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0651_
timestamp 1667941163
transform 1 0 22540 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0652_
timestamp 1667941163
transform 1 0 10948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0653_
timestamp 1667941163
transform 1 0 34224 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0654_
timestamp 1667941163
transform 1 0 22264 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0655_
timestamp 1667941163
transform 1 0 26220 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0656_
timestamp 1667941163
transform 1 0 6532 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0657_
timestamp 1667941163
transform 1 0 6532 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0658_
timestamp 1667941163
transform 1 0 28520 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1667941163
transform 1 0 14076 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0660_
timestamp 1667941163
transform 1 0 15824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0661_
timestamp 1667941163
transform 1 0 28612 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0662_
timestamp 1667941163
transform 1 0 30636 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0663_
timestamp 1667941163
transform 1 0 21436 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1667941163
transform 1 0 6532 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0665_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 22356 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0666_
timestamp 1667941163
transform 1 0 8280 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0667_
timestamp 1667941163
transform 1 0 6532 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0668_
timestamp 1667941163
transform 1 0 27324 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0669_
timestamp 1667941163
transform 1 0 32936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0670_
timestamp 1667941163
transform 1 0 30360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0671_
timestamp 1667941163
transform 1 0 30360 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0672_
timestamp 1667941163
transform 1 0 6440 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0673_
timestamp 1667941163
transform 1 0 27784 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1667941163
transform 1 0 8004 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0675_
timestamp 1667941163
transform 1 0 9292 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0676_
timestamp 1667941163
transform 1 0 23000 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 1667941163
transform 1 0 6256 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0678_
timestamp 1667941163
transform 1 0 35420 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0679_
timestamp 1667941163
transform 1 0 10396 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0680_
timestamp 1667941163
transform 1 0 14444 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0681_
timestamp 1667941163
transform 1 0 22632 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1667941163
transform 1 0 5060 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0683_
timestamp 1667941163
transform 1 0 9108 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0684_
timestamp 1667941163
transform 1 0 18308 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0685_
timestamp 1667941163
transform 1 0 25208 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1667941163
transform 1 0 5336 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0687_
timestamp 1667941163
transform 1 0 31004 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0688_
timestamp 1667941163
transform 1 0 32292 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1667941163
transform 1 0 15916 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0690_
timestamp 1667941163
transform 1 0 3956 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1667941163
transform 1 0 9108 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0692_
timestamp 1667941163
transform 1 0 32292 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1667941163
transform 1 0 33488 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0694_
timestamp 1667941163
transform 1 0 24564 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0695_
timestamp 1667941163
transform 1 0 25760 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0696_
timestamp 1667941163
transform 1 0 29716 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0697_
timestamp 1667941163
transform 1 0 11960 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0698_
timestamp 1667941163
transform 1 0 29532 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1667941163
transform 1 0 21804 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0700_
timestamp 1667941163
transform 1 0 7728 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0701_
timestamp 1667941163
transform 1 0 29716 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0702_
timestamp 1667941163
transform 1 0 25852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0703_
timestamp 1667941163
transform 1 0 15364 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0704_
timestamp 1667941163
transform 1 0 13800 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1667941163
transform 1 0 6256 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0706_
timestamp 1667941163
transform 1 0 6532 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0707_
timestamp 1667941163
transform 1 0 27140 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0708_
timestamp 1667941163
transform 1 0 22448 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0709_
timestamp 1667941163
transform 1 0 28520 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0710_
timestamp 1667941163
transform 1 0 29716 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0711_
timestamp 1667941163
transform 1 0 28612 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0712_
timestamp 1667941163
transform 1 0 8464 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1667941163
transform 1 0 27876 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0714_
timestamp 1667941163
transform 1 0 10672 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1667941163
transform 1 0 15088 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1667941163
transform 1 0 27968 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1667941163
transform 1 0 30084 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1667941163
transform 1 0 21988 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0719_
timestamp 1667941163
transform 1 0 29716 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1667941163
transform 1 0 11684 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1667941163
transform 1 0 30176 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0722_
timestamp 1667941163
transform 1 0 31464 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0723_
timestamp 1667941163
transform 1 0 3588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1667941163
transform 1 0 2576 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0725_
timestamp 1667941163
transform 1 0 24564 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1667941163
transform 1 0 33488 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0727_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6532 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0728_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14720 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0729_
timestamp 1667941163
transform 1 0 15456 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1667941163
transform 1 0 3864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1667941163
transform 1 0 2576 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1667941163
transform 1 0 6164 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1667941163
transform 1 0 6440 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1667941163
transform 1 0 6808 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1667941163
transform 1 0 13524 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0736_
timestamp 1667941163
transform 1 0 17664 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1667941163
transform 1 0 2576 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1667941163
transform 1 0 1932 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1667941163
transform 1 0 3220 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _0740_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16100 0 1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1667941163
transform 1 0 5980 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1667941163
transform 1 0 2576 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1667941163
transform 1 0 5796 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1667941163
transform 1 0 5796 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1667941163
transform 1 0 5796 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1667941163
transform 1 0 12696 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1667941163
transform 1 0 20608 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1667941163
transform 1 0 3956 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1667941163
transform 1 0 27140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1667941163
transform 1 0 26772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0751_
timestamp 1667941163
transform 1 0 11868 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1667941163
transform 1 0 6808 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0753_
timestamp 1667941163
transform 1 0 16008 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1667941163
transform 1 0 3588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0755_
timestamp 1667941163
transform 1 0 3220 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0756_
timestamp 1667941163
transform 1 0 5152 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1667941163
transform 1 0 5152 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 1667941163
transform 1 0 5336 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0759_
timestamp 1667941163
transform 1 0 3864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0760_
timestamp 1667941163
transform 1 0 5152 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1667941163
transform 1 0 10120 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0762_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 11316 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1667941163
transform 1 0 4876 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 1667941163
transform 1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1667941163
transform 1 0 3220 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0766_
timestamp 1667941163
transform 1 0 3312 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1667941163
transform 1 0 9660 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1667941163
transform 1 0 2300 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0769_
timestamp 1667941163
transform 1 0 7084 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1667941163
transform 1 0 22540 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1667941163
transform 1 0 15272 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1667941163
transform 1 0 5796 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0773_
timestamp 1667941163
transform 1 0 14260 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1667941163
transform 1 0 29072 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0775_
timestamp 1667941163
transform 1 0 29716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1667941163
transform 1 0 31004 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 1667941163
transform 1 0 31556 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1667941163
transform 1 0 28428 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1667941163
transform 1 0 2116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1667941163
transform 1 0 4508 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1667941163
transform 1 0 5796 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1667941163
transform 1 0 5520 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0783_
timestamp 1667941163
transform 1 0 5152 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0784_
timestamp 1667941163
transform 1 0 12052 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0785_
timestamp 1667941163
transform 1 0 10948 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0786_
timestamp 1667941163
transform 1 0 5520 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1667941163
transform 1 0 4508 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 1667941163
transform 1 0 16836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1667941163
transform 1 0 5796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0790_
timestamp 1667941163
transform 1 0 5796 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0791_
timestamp 1667941163
transform 1 0 12052 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 1667941163
transform 1 0 10948 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1667941163
transform 1 0 16100 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0794_
timestamp 1667941163
transform 1 0 22816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0795_
timestamp 1667941163
transform 1 0 12788 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1667941163
transform 1 0 2944 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0797_
timestamp 1667941163
transform 1 0 4600 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1667941163
transform 1 0 2668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0799_
timestamp 1667941163
transform 1 0 4692 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1667941163
transform 1 0 2576 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1667941163
transform 1 0 27140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0802_
timestamp 1667941163
transform 1 0 11684 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0803_
timestamp 1667941163
transform 1 0 8372 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0804_
timestamp 1667941163
transform 1 0 5152 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0805_
timestamp 1667941163
transform 1 0 4232 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0806_
timestamp 1667941163
transform 1 0 14812 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0807_
timestamp 1667941163
transform 1 0 7084 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1667941163
transform 1 0 3220 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0809_
timestamp 1667941163
transform 1 0 23828 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0810_
timestamp 1667941163
transform 1 0 16560 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0811_
timestamp 1667941163
transform 1 0 14904 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1667941163
transform 1 0 4232 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0813_
timestamp 1667941163
transform 1 0 3220 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0814_
timestamp 1667941163
transform 1 0 12236 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0815_
timestamp 1667941163
transform 1 0 29624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1667941163
transform 1 0 30912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0817_
timestamp 1667941163
transform 1 0 16836 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0818_
timestamp 1667941163
transform 1 0 31004 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1667941163
transform 1 0 28060 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1667941163
transform 1 0 28520 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0821_
timestamp 1667941163
transform 1 0 24656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1667941163
transform 1 0 10304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0823_
timestamp 1667941163
transform 1 0 6532 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0824_
timestamp 1667941163
transform 1 0 3220 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0825_
timestamp 1667941163
transform 1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0826_
timestamp 1667941163
transform 1 0 28428 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0827_
timestamp 1667941163
transform 1 0 31188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0828_
timestamp 1667941163
transform 1 0 10120 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0829_
timestamp 1667941163
transform 1 0 19780 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1667941163
transform 1 0 18676 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1667941163
transform 1 0 12880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0832_
timestamp 1667941163
transform 1 0 4508 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1667941163
transform 1 0 3220 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1667941163
transform 1 0 10948 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1667941163
transform 1 0 18952 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1667941163
transform 1 0 18032 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1667941163
transform 1 0 4876 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0838_
timestamp 1667941163
transform 1 0 10764 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0839_
timestamp 1667941163
transform 1 0 13248 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0840_
timestamp 1667941163
transform 1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1667941163
transform 1 0 23184 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1667941163
transform 1 0 22356 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0843_
timestamp 1667941163
transform 1 0 23644 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0844_
timestamp 1667941163
transform 1 0 25668 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0845_
timestamp 1667941163
transform 1 0 23736 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0846_
timestamp 1667941163
transform 1 0 5796 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0847_
timestamp 1667941163
transform 1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0848_
timestamp 1667941163
transform 1 0 25024 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0849_
timestamp 1667941163
transform 1 0 9108 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0850_
timestamp 1667941163
transform 1 0 26128 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0851_
timestamp 1667941163
transform 1 0 21252 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0852_
timestamp 1667941163
transform 1 0 23092 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0853_
timestamp 1667941163
transform 1 0 22908 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0854_
timestamp 1667941163
transform 1 0 2300 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0855_
timestamp 1667941163
transform 1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0856_
timestamp 1667941163
transform 1 0 23736 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0857_
timestamp 1667941163
transform 1 0 2576 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _0858_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4600 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0859_
timestamp 1667941163
transform 1 0 4232 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0860_
timestamp 1667941163
transform 1 0 11960 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0861_
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0862_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 12328 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0863_
timestamp 1667941163
transform 1 0 14444 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0864_
timestamp 1667941163
transform 1 0 17112 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0865_
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0866_
timestamp 1667941163
transform 1 0 4232 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0867_
timestamp 1667941163
transform 1 0 9292 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0868_
timestamp 1667941163
transform 1 0 4232 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0869_
timestamp 1667941163
transform 1 0 7176 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0870_
timestamp 1667941163
transform 1 0 11868 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0871_
timestamp 1667941163
transform 1 0 9108 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0872_
timestamp 1667941163
transform 1 0 6808 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0873_
timestamp 1667941163
transform 1 0 13340 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0874_
timestamp 1667941163
transform 1 0 17020 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0875_
timestamp 1667941163
transform 1 0 14536 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0876_
timestamp 1667941163
transform 1 0 17112 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0877_
timestamp 1667941163
transform 1 0 19688 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0878_
timestamp 1667941163
transform 1 0 14260 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0879_
timestamp 1667941163
transform 1 0 13340 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0880_
timestamp 1667941163
transform 1 0 11776 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0881_
timestamp 1667941163
transform 1 0 6716 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0882_
timestamp 1667941163
transform 1 0 9660 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0883_
timestamp 1667941163
transform 1 0 9108 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0884_
timestamp 1667941163
transform 1 0 4232 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0885_
timestamp 1667941163
transform 1 0 7728 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0886_
timestamp 1667941163
transform 1 0 11868 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0887_
timestamp 1667941163
transform 1 0 11316 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0888_
timestamp 1667941163
transform 1 0 11684 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0889_
timestamp 1667941163
transform 1 0 6716 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0890_
timestamp 1667941163
transform 1 0 14536 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0891_
timestamp 1667941163
transform 1 0 9384 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0892_
timestamp 1667941163
transform 1 0 11960 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0893_
timestamp 1667941163
transform 1 0 4508 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0894_
timestamp 1667941163
transform 1 0 12052 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0895_
timestamp 1667941163
transform 1 0 19412 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0896_
timestamp 1667941163
transform 1 0 16560 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0897_
timestamp 1667941163
transform 1 0 11040 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0898_
timestamp 1667941163
transform 1 0 19504 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0899_
timestamp 1667941163
transform 1 0 19504 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0900_
timestamp 1667941163
transform 1 0 21988 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0901_
timestamp 1667941163
transform 1 0 17112 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0902_
timestamp 1667941163
transform 1 0 16928 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0903_
timestamp 1667941163
transform 1 0 6716 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0904_
timestamp 1667941163
transform 1 0 8648 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0905_
timestamp 1667941163
transform 1 0 11868 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0906_
timestamp 1667941163
transform 1 0 14444 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0907_
timestamp 1667941163
transform 1 0 11960 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0908_
timestamp 1667941163
transform 1 0 11684 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0909_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 10396 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0910_
timestamp 1667941163
transform 1 0 9108 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0911_
timestamp 1667941163
transform 1 0 16836 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0912_
timestamp 1667941163
transform 1 0 9292 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0913_
timestamp 1667941163
transform 1 0 6808 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0914_
timestamp 1667941163
transform 1 0 9476 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0915_
timestamp 1667941163
transform 1 0 14260 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0916_
timestamp 1667941163
transform 1 0 15916 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0917_
timestamp 1667941163
transform 1 0 19596 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0918_
timestamp 1667941163
transform 1 0 14536 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0919_
timestamp 1667941163
transform 1 0 14260 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0920_
timestamp 1667941163
transform 1 0 6808 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0921_
timestamp 1667941163
transform 1 0 7084 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0922_
timestamp 1667941163
transform 1 0 7820 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0923_
timestamp 1667941163
transform 1 0 19412 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0924_
timestamp 1667941163
transform 1 0 14352 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0925_
timestamp 1667941163
transform 1 0 12512 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0926_
timestamp 1667941163
transform 1 0 6808 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0927_
timestamp 1667941163
transform 1 0 7268 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0928_
timestamp 1667941163
transform 1 0 7912 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0929_
timestamp 1667941163
transform 1 0 11684 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0930_
timestamp 1667941163
transform 1 0 17112 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0931_
timestamp 1667941163
transform 1 0 14628 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0932_
timestamp 1667941163
transform 1 0 13984 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0933_
timestamp 1667941163
transform 1 0 6808 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0934_
timestamp 1667941163
transform 1 0 8556 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0935_
timestamp 1667941163
transform 1 0 12880 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0936_
timestamp 1667941163
transform 1 0 17112 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0937_
timestamp 1667941163
transform 1 0 17020 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0938_
timestamp 1667941163
transform 1 0 19412 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0939_
timestamp 1667941163
transform 1 0 21712 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0940_
timestamp 1667941163
transform 1 0 19688 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0941_
timestamp 1667941163
transform 1 0 17204 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0942_
timestamp 1667941163
transform 1 0 14352 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0943_
timestamp 1667941163
transform 1 0 14168 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0944_
timestamp 1667941163
transform 1 0 9568 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0945_
timestamp 1667941163
transform 1 0 9384 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0946_
timestamp 1667941163
transform 1 0 18308 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0947_
timestamp 1667941163
transform 1 0 19228 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0948_
timestamp 1667941163
transform 1 0 17204 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0949_
timestamp 1667941163
transform 1 0 16744 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0950_
timestamp 1667941163
transform 1 0 19228 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0951_
timestamp 1667941163
transform 1 0 6808 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0952_
timestamp 1667941163
transform 1 0 7084 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0953_
timestamp 1667941163
transform 1 0 14168 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0954_
timestamp 1667941163
transform 1 0 16928 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0955_
timestamp 1667941163
transform 1 0 16008 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0956_
timestamp 1667941163
transform 1 0 6716 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0957_
timestamp 1667941163
transform 1 0 11684 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0958_
timestamp 1667941163
transform 1 0 19964 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0959_
timestamp 1667941163
transform 1 0 19044 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0960_
timestamp 1667941163
transform 1 0 16836 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0961_
timestamp 1667941163
transform 1 0 19964 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0962_
timestamp 1667941163
transform 1 0 19412 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0963_
timestamp 1667941163
transform 1 0 19412 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0964_
timestamp 1667941163
transform 1 0 7728 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0965_
timestamp 1667941163
transform 1 0 19412 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0966_
timestamp 1667941163
transform 1 0 16836 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0967_
timestamp 1667941163
transform 1 0 13984 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0968_
timestamp 1667941163
transform 1 0 17480 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0969_
timestamp 1667941163
transform 1 0 19688 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0970_
timestamp 1667941163
transform 1 0 18768 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0971_
timestamp 1667941163
transform 1 0 19780 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0972_
timestamp 1667941163
transform 1 0 6716 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0973_
timestamp 1667941163
transform 1 0 4508 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0974_
timestamp 1667941163
transform 1 0 19780 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0975_
timestamp 1667941163
transform 1 0 11684 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _1002_
timestamp 1667941163
transform 1 0 22080 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1003_
timestamp 1667941163
transform 1 0 34316 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1004_
timestamp 1667941163
transform 1 0 30728 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1005_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 28060 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1006_
timestamp 1667941163
transform 1 0 3864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1007_
timestamp 1667941163
transform 1 0 6256 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1008_
timestamp 1667941163
transform 1 0 29992 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1009_
timestamp 1667941163
transform 1 0 32936 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1010_
timestamp 1667941163
transform 1 0 27140 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1011_
timestamp 1667941163
transform 1 0 34960 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1012_
timestamp 1667941163
transform 1 0 34868 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1013_
timestamp 1667941163
transform 1 0 35144 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1014_
timestamp 1667941163
transform 1 0 14720 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1015_
timestamp 1667941163
transform 1 0 32476 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1016_
timestamp 1667941163
transform 1 0 29624 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1017_
timestamp 1667941163
transform 1 0 27968 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1018_
timestamp 1667941163
transform 1 0 33672 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1019_
timestamp 1667941163
transform 1 0 32108 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1020_
timestamp 1667941163
transform 1 0 3864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1021_
timestamp 1667941163
transform 1 0 15088 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1022_
timestamp 1667941163
transform 1 0 36616 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1023_
timestamp 1667941163
transform 1 0 27140 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1024_
timestamp 1667941163
transform 1 0 16836 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1025_
timestamp 1667941163
transform 1 0 19412 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1026_
timestamp 1667941163
transform 1 0 31004 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1027_
timestamp 1667941163
transform 1 0 2300 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1028_
timestamp 1667941163
transform 1 0 17388 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1029_
timestamp 1667941163
transform 1 0 32752 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1030_
timestamp 1667941163
transform 1 0 36616 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1031_
timestamp 1667941163
transform 1 0 10856 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1032_
timestamp 1667941163
transform 1 0 23276 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1033_
timestamp 1667941163
transform 1 0 27324 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1034_
timestamp 1667941163
transform 1 0 37352 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1035_
timestamp 1667941163
transform 1 0 28336 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1036_
timestamp 1667941163
transform 1 0 19320 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1037_
timestamp 1667941163
transform 1 0 2944 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1038_
timestamp 1667941163
transform 1 0 4508 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1039_
timestamp 1667941163
transform 1 0 4140 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1040_
timestamp 1667941163
transform 1 0 15456 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1041_
timestamp 1667941163
transform 1 0 3956 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1042_
timestamp 1667941163
transform 1 0 7084 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1043_
timestamp 1667941163
transform 1 0 37812 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1044_
timestamp 1667941163
transform 1 0 24564 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1045_
timestamp 1667941163
transform 1 0 36892 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1046_
timestamp 1667941163
transform 1 0 37812 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1047_
timestamp 1667941163
transform 1 0 9016 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1048_
timestamp 1667941163
transform 1 0 21988 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1049_
timestamp 1667941163
transform 1 0 4508 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1050_
timestamp 1667941163
transform 1 0 1932 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1051_
timestamp 1667941163
transform 1 0 23828 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1052_
timestamp 1667941163
transform 1 0 1748 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1053_
timestamp 1667941163
transform 1 0 22264 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1054_
timestamp 1667941163
transform 1 0 10396 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1055_
timestamp 1667941163
transform 1 0 20056 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1056_
timestamp 1667941163
transform 1 0 14996 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1057_
timestamp 1667941163
transform 1 0 37812 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1058_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14444 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1059_
timestamp 1667941163
transform 1 0 10764 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1060_
timestamp 1667941163
transform 1 0 26128 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1060__142 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 27784 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1061_
timestamp 1667941163
transform 1 0 18308 0 -1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1062_
timestamp 1667941163
transform 1 0 12972 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1063_
timestamp 1667941163
transform 1 0 10120 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1064_
timestamp 1667941163
transform 1 0 21068 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1065_
timestamp 1667941163
transform 1 0 17020 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1066_
timestamp 1667941163
transform 1 0 11868 0 -1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1067_
timestamp 1667941163
transform 1 0 21988 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1068_
timestamp 1667941163
transform 1 0 20976 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1069_
timestamp 1667941163
transform 1 0 22264 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1070_
timestamp 1667941163
transform 1 0 8648 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1071_
timestamp 1667941163
transform 1 0 18308 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1072__143
timestamp 1667941163
transform 1 0 4508 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1072_
timestamp 1667941163
transform 1 0 7452 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1073_
timestamp 1667941163
transform 1 0 7452 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1074_
timestamp 1667941163
transform 1 0 15180 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1075_
timestamp 1667941163
transform 1 0 16284 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1076_
timestamp 1667941163
transform 1 0 8280 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1077_
timestamp 1667941163
transform 1 0 12144 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1078_
timestamp 1667941163
transform 1 0 14720 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1079_
timestamp 1667941163
transform 1 0 9108 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1080_
timestamp 1667941163
transform 1 0 14536 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1081_
timestamp 1667941163
transform 1 0 17848 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1082_
timestamp 1667941163
transform 1 0 22816 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1083_
timestamp 1667941163
transform 1 0 23092 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1084_
timestamp 1667941163
transform 1 0 27140 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1084__144
timestamp 1667941163
transform 1 0 27784 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1085_
timestamp 1667941163
transform 1 0 17388 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1086_
timestamp 1667941163
transform 1 0 17480 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1087_
timestamp 1667941163
transform 1 0 12328 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1088_
timestamp 1667941163
transform 1 0 24196 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1089_
timestamp 1667941163
transform 1 0 12972 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1090_
timestamp 1667941163
transform 1 0 24564 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1091_
timestamp 1667941163
transform 1 0 23552 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1092_
timestamp 1667941163
transform 1 0 2760 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1093_
timestamp 1667941163
transform 1 0 22908 0 1 2176
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1094_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6256 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1095_
timestamp 1667941163
transform 1 0 11684 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1096_
timestamp 1667941163
transform 1 0 5244 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1096__145
timestamp 1667941163
transform 1 0 5612 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1097_
timestamp 1667941163
transform 1 0 22632 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1098_
timestamp 1667941163
transform 1 0 23184 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1099_
timestamp 1667941163
transform 1 0 21160 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1100_
timestamp 1667941163
transform 1 0 12420 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1101_
timestamp 1667941163
transform 1 0 13248 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1102_
timestamp 1667941163
transform 1 0 7268 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1103_
timestamp 1667941163
transform 1 0 6624 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1104_
timestamp 1667941163
transform 1 0 4140 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1105_
timestamp 1667941163
transform 1 0 5244 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1106_
timestamp 1667941163
transform 1 0 20332 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1107_
timestamp 1667941163
transform 1 0 23092 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1108_
timestamp 1667941163
transform 1 0 25300 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1108__146
timestamp 1667941163
transform 1 0 26220 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1109_
timestamp 1667941163
transform 1 0 15916 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1110_
timestamp 1667941163
transform 1 0 19228 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1111_
timestamp 1667941163
transform 1 0 11224 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1112_
timestamp 1667941163
transform 1 0 25576 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1113_
timestamp 1667941163
transform 1 0 25760 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1114_
timestamp 1667941163
transform 1 0 4048 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1115_
timestamp 1667941163
transform 1 0 23092 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1116_
timestamp 1667941163
transform 1 0 15180 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1117_
timestamp 1667941163
transform 1 0 23828 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1118_
timestamp 1667941163
transform 1 0 24840 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1119_
timestamp 1667941163
transform 1 0 24564 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1120__147
timestamp 1667941163
transform 1 0 28704 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1120_
timestamp 1667941163
transform 1 0 26496 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1121_
timestamp 1667941163
transform 1 0 8188 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1122_
timestamp 1667941163
transform 1 0 15180 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1123_
timestamp 1667941163
transform 1 0 23552 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1124_
timestamp 1667941163
transform 1 0 12512 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1125_
timestamp 1667941163
transform 1 0 14536 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1126_
timestamp 1667941163
transform 1 0 25208 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1127_
timestamp 1667941163
transform 1 0 24840 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1128_
timestamp 1667941163
transform 1 0 6808 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1129_
timestamp 1667941163
transform 1 0 23552 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1130_
timestamp 1667941163
transform 1 0 12604 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1131_
timestamp 1667941163
transform 1 0 13248 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1132_
timestamp 1667941163
transform 1 0 8372 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1133_
timestamp 1667941163
transform 1 0 14260 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1133__148
timestamp 1667941163
transform 1 0 9476 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1134_
timestamp 1667941163
transform 1 0 14628 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1135_
timestamp 1667941163
transform 1 0 20700 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1136_
timestamp 1667941163
transform 1 0 10120 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1137_
timestamp 1667941163
transform 1 0 24564 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1138_
timestamp 1667941163
transform 1 0 13248 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1139_
timestamp 1667941163
transform 1 0 24012 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1140_
timestamp 1667941163
transform 1 0 19872 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1141_
timestamp 1667941163
transform 1 0 22908 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1142_
timestamp 1667941163
transform 1 0 12604 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1143_
timestamp 1667941163
transform 1 0 13064 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1144_
timestamp 1667941163
transform 1 0 17480 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1145_
timestamp 1667941163
transform 1 0 19412 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1145__149
timestamp 1667941163
transform 1 0 19596 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1146_
timestamp 1667941163
transform 1 0 21988 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1147_
timestamp 1667941163
transform 1 0 24656 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1148_
timestamp 1667941163
transform 1 0 10396 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1149_
timestamp 1667941163
transform 1 0 26128 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1150_
timestamp 1667941163
transform 1 0 10028 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1151_
timestamp 1667941163
transform 1 0 20240 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1152_
timestamp 1667941163
transform 1 0 23368 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1153_
timestamp 1667941163
transform 1 0 27140 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1154_
timestamp 1667941163
transform 1 0 25852 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1155_
timestamp 1667941163
transform 1 0 25760 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1156_
timestamp 1667941163
transform 1 0 9568 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1157__150
timestamp 1667941163
transform 1 0 25668 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1157_
timestamp 1667941163
transform 1 0 24472 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1158_
timestamp 1667941163
transform 1 0 6900 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1159_
timestamp 1667941163
transform 1 0 26404 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1160_
timestamp 1667941163
transform 1 0 12052 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1161_
timestamp 1667941163
transform 1 0 24656 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1162_
timestamp 1667941163
transform 1 0 25852 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1163_
timestamp 1667941163
transform 1 0 24840 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1164_
timestamp 1667941163
transform 1 0 25484 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1165_
timestamp 1667941163
transform 1 0 23828 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1166_
timestamp 1667941163
transform 1 0 12328 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1167_
timestamp 1667941163
transform 1 0 11684 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1168_
timestamp 1667941163
transform 1 0 11316 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1169__151
timestamp 1667941163
transform 1 0 9476 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1169_
timestamp 1667941163
transform 1 0 9660 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1170_
timestamp 1667941163
transform 1 0 14628 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1171_
timestamp 1667941163
transform 1 0 12788 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1172_
timestamp 1667941163
transform 1 0 16468 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1173_
timestamp 1667941163
transform 1 0 9936 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1174_
timestamp 1667941163
transform 1 0 12880 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1175_
timestamp 1667941163
transform 1 0 10212 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1176_
timestamp 1667941163
transform 1 0 7084 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1177_
timestamp 1667941163
transform 1 0 23092 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1178_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17480 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1179_
timestamp 1667941163
transform 1 0 19596 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1180__152
timestamp 1667941163
transform 1 0 22448 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1180_
timestamp 1667941163
transform 1 0 22080 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1181_
timestamp 1667941163
transform 1 0 4416 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1182_
timestamp 1667941163
transform 1 0 15916 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1183_
timestamp 1667941163
transform 1 0 25024 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1184_
timestamp 1667941163
transform 1 0 16928 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1185_
timestamp 1667941163
transform 1 0 4048 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1186_
timestamp 1667941163
transform 1 0 25024 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1187_
timestamp 1667941163
transform 1 0 25760 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1188__153
timestamp 1667941163
transform 1 0 32292 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1188_
timestamp 1667941163
transform 1 0 27140 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1189_
timestamp 1667941163
transform 1 0 24104 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1190_
timestamp 1667941163
transform 1 0 24564 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1191_
timestamp 1667941163
transform 1 0 21344 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1192_
timestamp 1667941163
transform 1 0 22540 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1193_
timestamp 1667941163
transform 1 0 23092 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1194_
timestamp 1667941163
transform 1 0 19596 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1195_
timestamp 1667941163
transform 1 0 22632 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1196__154
timestamp 1667941163
transform 1 0 19412 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1196_
timestamp 1667941163
transform 1 0 18768 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1197_
timestamp 1667941163
transform 1 0 14260 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1198_
timestamp 1667941163
transform 1 0 26956 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _1199_
timestamp 1667941163
transform 1 0 24564 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1200_
timestamp 1667941163
transform 1 0 19412 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1201_
timestamp 1667941163
transform 1 0 24564 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1202_
timestamp 1667941163
transform 1 0 18216 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1203_
timestamp 1667941163
transform 1 0 19780 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1203__155
timestamp 1667941163
transform 1 0 20332 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1204_
timestamp 1667941163
transform 1 0 10396 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1205_
timestamp 1667941163
transform 1 0 17112 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1206_
timestamp 1667941163
transform 1 0 18124 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1207_
timestamp 1667941163
transform 1 0 22540 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1208_
timestamp 1667941163
transform 1 0 22724 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1209__156
timestamp 1667941163
transform 1 0 20056 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1209_
timestamp 1667941163
transform 1 0 20056 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1210_
timestamp 1667941163
transform 1 0 25852 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1211_
timestamp 1667941163
transform 1 0 26864 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1212_
timestamp 1667941163
transform 1 0 18584 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1213_
timestamp 1667941163
transform 1 0 25760 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1214_
timestamp 1667941163
transform 1 0 12880 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1215_
timestamp 1667941163
transform 1 0 13064 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1215__157
timestamp 1667941163
transform 1 0 11316 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1216_
timestamp 1667941163
transform 1 0 11776 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1217_
timestamp 1667941163
transform 1 0 12788 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1218_
timestamp 1667941163
transform 1 0 11960 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1219_
timestamp 1667941163
transform 1 0 11684 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1220_
timestamp 1667941163
transform 1 0 29256 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1221__158
timestamp 1667941163
transform 1 0 30728 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1221_
timestamp 1667941163
transform 1 0 30636 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1222_
timestamp 1667941163
transform 1 0 23184 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1223_
timestamp 1667941163
transform 1 0 27140 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1224_
timestamp 1667941163
transform 1 0 28520 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1225_
timestamp 1667941163
transform 1 0 21988 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1226_
timestamp 1667941163
transform 1 0 24380 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1227__159
timestamp 1667941163
transform 1 0 23092 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1227_
timestamp 1667941163
transform 1 0 23092 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1228_
timestamp 1667941163
transform 1 0 24564 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1229_
timestamp 1667941163
transform 1 0 24564 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1230_
timestamp 1667941163
transform 1 0 21988 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1231_
timestamp 1667941163
transform 1 0 16744 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1232_
timestamp 1667941163
transform 1 0 28428 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1233__160
timestamp 1667941163
transform 1 0 29808 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1233_
timestamp 1667941163
transform 1 0 28704 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1234_
timestamp 1667941163
transform 1 0 16836 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1235_
timestamp 1667941163
transform 1 0 27968 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1236_
timestamp 1667941163
transform 1 0 26680 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1237_
timestamp 1667941163
transform 1 0 27692 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1238_
timestamp 1667941163
transform 1 0 13064 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1239__161
timestamp 1667941163
transform 1 0 14720 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1239_
timestamp 1667941163
transform 1 0 14628 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1240_
timestamp 1667941163
transform 1 0 14352 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1241_
timestamp 1667941163
transform 1 0 11960 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1242_
timestamp 1667941163
transform 1 0 15272 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1243_
timestamp 1667941163
transform 1 0 14536 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1244__162
timestamp 1667941163
transform 1 0 29348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1244_
timestamp 1667941163
transform 1 0 29256 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1245_
timestamp 1667941163
transform 1 0 24564 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1246_
timestamp 1667941163
transform 1 0 29716 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1247_
timestamp 1667941163
transform 1 0 25668 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1248__163
timestamp 1667941163
transform 1 0 29256 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1248_
timestamp 1667941163
transform 1 0 28428 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1249_
timestamp 1667941163
transform 1 0 15088 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1250_
timestamp 1667941163
transform 1 0 27140 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1251_
timestamp 1667941163
transform 1 0 15456 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1252__164
timestamp 1667941163
transform 1 0 27876 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1252_
timestamp 1667941163
transform 1 0 28152 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1253_
timestamp 1667941163
transform 1 0 25300 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1254_
timestamp 1667941163
transform 1 0 29716 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1255_
timestamp 1667941163
transform 1 0 17848 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1256__165
timestamp 1667941163
transform 1 0 2392 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1256_
timestamp 1667941163
transform 1 0 2392 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1257_
timestamp 1667941163
transform 1 0 2208 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1258_
timestamp 1667941163
transform 1 0 2484 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1259_
timestamp 1667941163
transform 1 0 1932 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1260_
timestamp 1667941163
transform 1 0 29716 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1260__166
timestamp 1667941163
transform 1 0 29256 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1261_
timestamp 1667941163
transform 1 0 27324 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1262_
timestamp 1667941163
transform 1 0 28336 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1263_
timestamp 1667941163
transform 1 0 27508 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 11960 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk
timestamp 1667941163
transform 1 0 6532 0 -1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1667941163
transform 1 0 5428 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1667941163
transform 1 0 9844 0 -1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1667941163
transform 1 0 10304 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1667941163
transform 1 0 7176 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1667941163
transform 1 0 9108 0 1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1667941163
transform 1 0 10212 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1667941163
transform 1 0 10212 0 -1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1667941163
transform 1 0 12788 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1667941163
transform 1 0 15364 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1667941163
transform 1 0 16928 0 -1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1667941163
transform 1 0 21988 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1667941163
transform 1 0 14628 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1667941163
transform 1 0 14904 0 -1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1667941163
transform 1 0 17940 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1667941163
transform 1 0 19412 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1667941163
transform 1 0 1564 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1667941163
transform 1 0 1564 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1667941163
transform 1 0 5244 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1667941163
transform 1 0 1932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1667941163
transform 1 0 35512 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1667941163
transform 1 0 32936 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1667941163
transform 1 0 1564 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1667941163
transform 1 0 1564 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1667941163
transform 1 0 18124 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1667941163
transform 1 0 2300 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1667941163
transform 1 0 4784 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1667941163
transform 1 0 25852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1667941163
transform 1 0 6532 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1667941163
transform 1 0 31648 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1667941163
transform 1 0 9108 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1667941163
transform 1 0 16468 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1667941163
transform 1 0 1564 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1667941163
transform 1 0 2208 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1667941163
transform 1 0 27876 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1667941163
transform 1 0 4508 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1667941163
transform 1 0 38088 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1667941163
transform 1 0 38088 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1667941163
transform 1 0 2944 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1667941163
transform 1 0 2852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1667941163
transform 1 0 38088 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1667941163
transform 1 0 14996 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1667941163
transform 1 0 38088 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1667941163
transform 1 0 38088 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1667941163
transform 1 0 32292 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1667941163
transform 1 0 3588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1667941163
transform 1 0 37260 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37444 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1667941163
transform 1 0 24564 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1667941163
transform 1 0 12328 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input35
timestamp 1667941163
transform 1 0 37444 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input36
timestamp 1667941163
transform 1 0 9108 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1667941163
transform 1 0 11684 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input38
timestamp 1667941163
transform 1 0 22632 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1667941163
transform 1 0 2300 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1667941163
transform 1 0 2668 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1667941163
transform 1 0 37996 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input42
timestamp 1667941163
transform 1 0 3956 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1667941163
transform 1 0 36708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1667941163
transform 1 0 1564 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45
timestamp 1667941163
transform 1 0 37444 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1667941163
transform 1 0 1564 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1667941163
transform 1 0 3956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1667941163
transform 1 0 1564 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1667941163
transform 1 0 16008 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50
timestamp 1667941163
transform 1 0 1564 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input51
timestamp 1667941163
transform 1 0 2024 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1667941163
transform 1 0 1564 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input53
timestamp 1667941163
transform 1 0 1564 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1667941163
transform 1 0 1564 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input55
timestamp 1667941163
transform 1 0 37444 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input56
timestamp 1667941163
transform 1 0 9108 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1667941163
transform 1 0 1564 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input58
timestamp 1667941163
transform 1 0 24564 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input59
timestamp 1667941163
transform 1 0 37444 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1667941163
transform 1 0 14260 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1667941163
transform 1 0 33580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1667941163
transform 1 0 3588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1667941163
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1667941163
transform 1 0 37996 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1667941163
transform 1 0 37996 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1667941163
transform 1 0 38088 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1667941163
transform 1 0 32292 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input68
timestamp 1667941163
transform 1 0 1564 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1667941163
transform 1 0 11960 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1667941163
transform 1 0 35236 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1667941163
transform 1 0 38088 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1667941163
transform 1 0 1564 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1667941163
transform 1 0 1564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1667941163
transform 1 0 3956 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1667941163
transform 1 0 21988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1667941163
transform 1 0 38088 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1667941163
transform 1 0 28520 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1667941163
transform 1 0 30360 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1667941163
transform 1 0 29716 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1667941163
transform 1 0 3312 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1667941163
transform 1 0 7176 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1667941163
transform 1 0 32292 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1667941163
transform 1 0 1564 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output84 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 29716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1667941163
transform 1 0 36156 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1667941163
transform 1 0 37996 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1667941163
transform 1 0 33580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1667941163
transform 1 0 1564 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1667941163
transform 1 0 1564 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1667941163
transform 1 0 20056 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1667941163
transform 1 0 37996 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1667941163
transform 1 0 35880 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1667941163
transform 1 0 19412 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1667941163
transform 1 0 34868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1667941163
transform 1 0 31004 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1667941163
transform 1 0 34868 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1667941163
transform 1 0 35880 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1667941163
transform 1 0 16008 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1667941163
transform 1 0 37996 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1667941163
transform 1 0 37996 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1667941163
transform 1 0 37996 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1667941163
transform 1 0 27784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1667941163
transform 1 0 1564 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1667941163
transform 1 0 32936 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1667941163
transform 1 0 1564 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1667941163
transform 1 0 30452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1667941163
transform 1 0 37996 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1667941163
transform 1 0 37996 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1667941163
transform 1 0 27140 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1667941163
transform 1 0 36616 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1667941163
transform 1 0 37444 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1667941163
transform 1 0 1564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1667941163
transform 1 0 5244 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1667941163
transform 1 0 37996 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1667941163
transform 1 0 1564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1667941163
transform 1 0 37996 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1667941163
transform 1 0 37996 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1667941163
transform 1 0 16836 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1667941163
transform 1 0 3128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1667941163
transform 1 0 37996 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1667941163
transform 1 0 37996 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1667941163
transform 1 0 37996 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1667941163
transform 1 0 1564 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1667941163
transform 1 0 37996 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1667941163
transform 1 0 37996 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1667941163
transform 1 0 36616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1667941163
transform 1 0 37996 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1667941163
transform 1 0 1564 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1667941163
transform 1 0 1564 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1667941163
transform 1 0 1564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1667941163
transform 1 0 2392 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1667941163
transform 1 0 1564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1667941163
transform 1 0 1564 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1667941163
transform 1 0 10396 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1667941163
transform 1 0 23276 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1667941163
transform 1 0 1564 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1667941163
transform 1 0 6532 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1667941163
transform 1 0 1656 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1667941163
transform 1 0 1564 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1667941163
transform 1 0 21160 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  sb_4__1__141
timestamp 1667941163
transform 1 0 38088 0 -1 4352
box -38 -48 314 592
<< labels >>
flabel metal3 s 200 19048 800 19168 0 FreeSans 480 0 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
port 0 nsew signal input
flabel metal3 s 200 7488 800 7608 0 FreeSans 480 0 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
port 1 nsew signal input
flabel metal2 s 5170 39200 5226 39800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 2 nsew signal input
flabel metal3 s 200 5448 800 5568 0 FreeSans 480 0 0 0 bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
port 3 nsew signal input
flabel metal2 s 35438 200 35494 800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
port 4 nsew signal input
flabel metal2 s 25778 200 25834 800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
port 5 nsew signal input
flabel metal3 s 200 22448 800 22568 0 FreeSans 480 0 0 0 bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_
port 6 nsew signal input
flabel metal3 s 200 6808 800 6928 0 FreeSans 480 0 0 0 bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_
port 7 nsew signal input
flabel metal2 s 18050 39200 18106 39800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_
port 8 nsew signal input
flabel metal3 s 200 38768 800 38888 0 FreeSans 480 0 0 0 bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_
port 9 nsew signal input
flabel metal2 s 12898 200 12954 800 0 FreeSans 224 90 0 0 ccff_head
port 10 nsew signal input
flabel metal2 s 28998 200 29054 800 0 FreeSans 224 90 0 0 ccff_tail
port 11 nsew signal tristate
flabel metal2 s 25778 39200 25834 39800 0 FreeSans 224 90 0 0 chanx_left_in[0]
port 12 nsew signal input
flabel metal2 s 5814 39200 5870 39800 0 FreeSans 224 90 0 0 chanx_left_in[10]
port 13 nsew signal input
flabel metal2 s 24490 200 24546 800 0 FreeSans 224 90 0 0 chanx_left_in[11]
port 14 nsew signal input
flabel metal2 s 9034 39200 9090 39800 0 FreeSans 224 90 0 0 chanx_left_in[12]
port 15 nsew signal input
flabel metal2 s 19982 200 20038 800 0 FreeSans 224 90 0 0 chanx_left_in[13]
port 16 nsew signal input
flabel metal3 s 200 17008 800 17128 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 17 nsew signal input
flabel metal3 s 200 2048 800 2168 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 18 nsew signal input
flabel metal2 s 27710 39200 27766 39800 0 FreeSans 224 90 0 0 chanx_left_in[16]
port 19 nsew signal input
flabel metal2 s 11610 200 11666 800 0 FreeSans 224 90 0 0 chanx_left_in[17]
port 20 nsew signal input
flabel metal3 s 39200 31968 39800 32088 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 21 nsew signal input
flabel metal3 s 39200 27208 39800 27328 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 22 nsew signal input
flabel metal2 s 9678 200 9734 800 0 FreeSans 224 90 0 0 chanx_left_in[2]
port 23 nsew signal input
flabel metal3 s 200 688 800 808 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 24 nsew signal input
flabel metal3 s 39200 8848 39800 8968 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 25 nsew signal input
flabel metal2 s 14830 39200 14886 39800 0 FreeSans 224 90 0 0 chanx_left_in[5]
port 26 nsew signal input
flabel metal3 s 39200 30608 39800 30728 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 27 nsew signal input
flabel metal3 s 39200 28568 39800 28688 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 28 nsew signal input
flabel metal2 s 32218 39200 32274 39800 0 FreeSans 224 90 0 0 chanx_left_in[8]
port 29 nsew signal input
flabel metal2 s 18050 200 18106 800 0 FreeSans 224 90 0 0 chanx_left_in[9]
port 30 nsew signal input
flabel metal2 s 36082 39200 36138 39800 0 FreeSans 224 90 0 0 chanx_left_out[0]
port 31 nsew signal tristate
flabel metal3 s 39200 12248 39800 12368 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 32 nsew signal tristate
flabel metal2 s 33506 200 33562 800 0 FreeSans 224 90 0 0 chanx_left_out[11]
port 33 nsew signal tristate
flabel metal3 s 200 30608 800 30728 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 34 nsew signal tristate
flabel metal3 s 200 15648 800 15768 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 35 nsew signal tristate
flabel metal3 s 39200 2048 39800 2168 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 36 nsew signal tristate
flabel metal2 s 19982 39200 20038 39800 0 FreeSans 224 90 0 0 chanx_left_out[15]
port 37 nsew signal tristate
flabel metal3 s 39200 35368 39800 35488 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 38 nsew signal tristate
flabel metal3 s 39200 8 39800 128 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 39 nsew signal tristate
flabel metal2 s 19338 39200 19394 39800 0 FreeSans 224 90 0 0 chanx_left_out[18]
port 40 nsew signal tristate
flabel metal2 s 34150 200 34206 800 0 FreeSans 224 90 0 0 chanx_left_out[1]
port 41 nsew signal tristate
flabel metal2 s 30930 39200 30986 39800 0 FreeSans 224 90 0 0 chanx_left_out[2]
port 42 nsew signal tristate
flabel metal2 s 34150 39200 34206 39800 0 FreeSans 224 90 0 0 chanx_left_out[3]
port 43 nsew signal tristate
flabel metal3 s 39200 37408 39800 37528 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 44 nsew signal tristate
flabel metal2 s 16118 39200 16174 39800 0 FreeSans 224 90 0 0 chanx_left_out[5]
port 45 nsew signal tristate
flabel metal3 s 39200 10888 39800 11008 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 46 nsew signal tristate
flabel metal3 s 39200 13608 39800 13728 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 47 nsew signal tristate
flabel metal3 s 39200 19048 39800 19168 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 48 nsew signal tristate
flabel metal2 s 27710 200 27766 800 0 FreeSans 224 90 0 0 chanx_left_out[9]
port 49 nsew signal tristate
flabel metal3 s 39200 38768 39800 38888 0 FreeSans 480 0 0 0 chany_bottom_in[0]
port 50 nsew signal input
flabel metal3 s 39200 32648 39800 32768 0 FreeSans 480 0 0 0 chany_bottom_in[10]
port 51 nsew signal input
flabel metal2 s 24490 39200 24546 39800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 52 nsew signal input
flabel metal2 s 12254 39200 12310 39800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 53 nsew signal input
flabel metal3 s 39200 23808 39800 23928 0 FreeSans 480 0 0 0 chany_bottom_in[13]
port 54 nsew signal input
flabel metal2 s 8390 39200 8446 39800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 55 nsew signal input
flabel metal2 s 11610 39200 11666 39800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 56 nsew signal input
flabel metal2 s 22558 39200 22614 39800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 57 nsew signal input
flabel metal2 s 10322 200 10378 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 58 nsew signal input
flabel metal2 s 2594 39200 2650 39800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 59 nsew signal input
flabel metal3 s 39200 14968 39800 15088 0 FreeSans 480 0 0 0 chany_bottom_in[1]
port 60 nsew signal input
flabel metal2 s 3882 39200 3938 39800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 61 nsew signal input
flabel metal3 s 39200 688 39800 808 0 FreeSans 480 0 0 0 chany_bottom_in[3]
port 62 nsew signal input
flabel metal3 s 200 14288 800 14408 0 FreeSans 480 0 0 0 chany_bottom_in[4]
port 63 nsew signal input
flabel metal3 s 39200 7488 39800 7608 0 FreeSans 480 0 0 0 chany_bottom_in[5]
port 64 nsew signal input
flabel metal3 s 200 28568 800 28688 0 FreeSans 480 0 0 0 chany_bottom_in[6]
port 65 nsew signal input
flabel metal2 s 16762 200 16818 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 66 nsew signal input
flabel metal3 s 200 21088 800 21208 0 FreeSans 480 0 0 0 chany_bottom_in[8]
port 67 nsew signal input
flabel metal2 s 16118 200 16174 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 68 nsew signal input
flabel metal3 s 200 24488 800 24608 0 FreeSans 480 0 0 0 chany_bottom_out[0]
port 69 nsew signal tristate
flabel metal2 s 32862 39200 32918 39800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 70 nsew signal tristate
flabel metal3 s 200 32648 800 32768 0 FreeSans 480 0 0 0 chany_bottom_out[11]
port 71 nsew signal tristate
flabel metal2 s 30286 200 30342 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 72 nsew signal tristate
flabel metal3 s 39200 25168 39800 25288 0 FreeSans 480 0 0 0 chany_bottom_out[13]
port 73 nsew signal tristate
flabel metal3 s 39200 5448 39800 5568 0 FreeSans 480 0 0 0 chany_bottom_out[14]
port 74 nsew signal tristate
flabel metal2 s 26422 39200 26478 39800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 75 nsew signal tristate
flabel metal2 s 39302 39200 39358 39800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 76 nsew signal tristate
flabel metal2 s 37370 39200 37426 39800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 77 nsew signal tristate
flabel metal2 s 662 200 718 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 78 nsew signal tristate
flabel metal2 s 5170 200 5226 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 79 nsew signal tristate
flabel metal2 s 38658 200 38714 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 80 nsew signal tristate
flabel metal3 s 200 13608 800 13728 0 FreeSans 480 0 0 0 chany_bottom_out[3]
port 81 nsew signal tristate
flabel metal3 s 39200 21768 39800 21888 0 FreeSans 480 0 0 0 chany_bottom_out[4]
port 82 nsew signal tristate
flabel metal3 s 39200 15648 39800 15768 0 FreeSans 480 0 0 0 chany_bottom_out[5]
port 83 nsew signal tristate
flabel metal2 s 16762 39200 16818 39800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 84 nsew signal tristate
flabel metal2 s 3238 200 3294 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 85 nsew signal tristate
flabel metal3 s 39200 3408 39800 3528 0 FreeSans 480 0 0 0 chany_bottom_out[8]
port 86 nsew signal tristate
flabel metal3 s 39200 17008 39800 17128 0 FreeSans 480 0 0 0 chany_bottom_out[9]
port 87 nsew signal tristate
flabel metal3 s 200 27208 800 27328 0 FreeSans 480 0 0 0 chany_top_in[0]
port 88 nsew signal input
flabel metal2 s 1950 39200 2006 39800 0 FreeSans 224 90 0 0 chany_top_in[10]
port 89 nsew signal input
flabel metal3 s 200 25848 800 25968 0 FreeSans 480 0 0 0 chany_top_in[11]
port 90 nsew signal input
flabel metal3 s 200 20408 800 20528 0 FreeSans 480 0 0 0 chany_top_in[12]
port 91 nsew signal input
flabel metal3 s 200 39448 800 39568 0 FreeSans 480 0 0 0 chany_top_in[13]
port 92 nsew signal input
flabel metal2 s 38658 39200 38714 39800 0 FreeSans 224 90 0 0 chany_top_in[14]
port 93 nsew signal input
flabel metal2 s 8390 200 8446 800 0 FreeSans 224 90 0 0 chany_top_in[15]
port 94 nsew signal input
flabel metal3 s 200 17688 800 17808 0 FreeSans 480 0 0 0 chany_top_in[16]
port 95 nsew signal input
flabel metal2 s 23202 200 23258 800 0 FreeSans 224 90 0 0 chany_top_in[17]
port 96 nsew signal input
flabel metal2 s 37370 200 37426 800 0 FreeSans 224 90 0 0 chany_top_in[18]
port 97 nsew signal input
flabel metal2 s 13542 39200 13598 39800 0 FreeSans 224 90 0 0 chany_top_in[1]
port 98 nsew signal input
flabel metal2 s 30930 200 30986 800 0 FreeSans 224 90 0 0 chany_top_in[2]
port 99 nsew signal input
flabel metal2 s 3882 200 3938 800 0 FreeSans 224 90 0 0 chany_top_in[3]
port 100 nsew signal input
flabel metal2 s 14830 200 14886 800 0 FreeSans 224 90 0 0 chany_top_in[4]
port 101 nsew signal input
flabel metal3 s 39200 4088 39800 4208 0 FreeSans 480 0 0 0 chany_top_in[5]
port 102 nsew signal input
flabel metal3 s 39200 29248 39800 29368 0 FreeSans 480 0 0 0 chany_top_in[6]
port 103 nsew signal input
flabel metal3 s 39200 20408 39800 20528 0 FreeSans 480 0 0 0 chany_top_in[7]
port 104 nsew signal input
flabel metal2 s 32218 200 32274 800 0 FreeSans 224 90 0 0 chany_top_in[8]
port 105 nsew signal input
flabel metal3 s 200 23808 800 23928 0 FreeSans 480 0 0 0 chany_top_in[9]
port 106 nsew signal input
flabel metal3 s 39200 10208 39800 10328 0 FreeSans 480 0 0 0 chany_top_out[0]
port 107 nsew signal tristate
flabel metal3 s 200 31968 800 32088 0 FreeSans 480 0 0 0 chany_top_out[10]
port 108 nsew signal tristate
flabel metal3 s 39200 22448 39800 22568 0 FreeSans 480 0 0 0 chany_top_out[11]
port 109 nsew signal tristate
flabel metal3 s 39200 34008 39800 34128 0 FreeSans 480 0 0 0 chany_top_out[12]
port 110 nsew signal tristate
flabel metal2 s 36726 200 36782 800 0 FreeSans 224 90 0 0 chany_top_out[13]
port 111 nsew signal tristate
flabel metal3 s 39200 36048 39800 36168 0 FreeSans 480 0 0 0 chany_top_out[14]
port 112 nsew signal tristate
flabel metal3 s 200 12248 800 12368 0 FreeSans 480 0 0 0 chany_top_out[15]
port 113 nsew signal tristate
flabel metal3 s 200 34008 800 34128 0 FreeSans 480 0 0 0 chany_top_out[16]
port 114 nsew signal tristate
flabel metal3 s 200 3408 800 3528 0 FreeSans 480 0 0 0 chany_top_out[17]
port 115 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 chany_top_out[18]
port 116 nsew signal tristate
flabel metal3 s 200 4088 800 4208 0 FreeSans 480 0 0 0 chany_top_out[1]
port 117 nsew signal tristate
flabel metal3 s 200 37408 800 37528 0 FreeSans 480 0 0 0 chany_top_out[2]
port 118 nsew signal tristate
flabel metal2 s 10322 39200 10378 39800 0 FreeSans 224 90 0 0 chany_top_out[3]
port 119 nsew signal tristate
flabel metal2 s 23202 39200 23258 39800 0 FreeSans 224 90 0 0 chany_top_out[4]
port 120 nsew signal tristate
flabel metal3 s 200 29248 800 29368 0 FreeSans 480 0 0 0 chany_top_out[5]
port 121 nsew signal tristate
flabel metal2 s 6458 200 6514 800 0 FreeSans 224 90 0 0 chany_top_out[6]
port 122 nsew signal tristate
flabel metal2 s 1950 200 2006 800 0 FreeSans 224 90 0 0 chany_top_out[7]
port 123 nsew signal tristate
flabel metal3 s 200 8848 800 8968 0 FreeSans 480 0 0 0 chany_top_out[8]
port 124 nsew signal tristate
flabel metal2 s 21270 39200 21326 39800 0 FreeSans 224 90 0 0 chany_top_out[9]
port 125 nsew signal tristate
flabel metal2 s 19338 200 19394 800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 126 nsew signal input
flabel metal2 s 35438 39200 35494 39800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 127 nsew signal input
flabel metal3 s 39200 6808 39800 6928 0 FreeSans 480 0 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
port 128 nsew signal input
flabel metal3 s 200 36048 800 36168 0 FreeSans 480 0 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
port 129 nsew signal input
flabel metal3 s 200 10888 800 11008 0 FreeSans 480 0 0 0 pReset
port 130 nsew signal input
flabel metal2 s 7102 200 7158 800 0 FreeSans 224 90 0 0 prog_clk
port 131 nsew signal input
flabel metal2 s 13542 200 13598 800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
port 132 nsew signal input
flabel metal2 s 21270 200 21326 800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
port 133 nsew signal input
flabel metal3 s 39200 25848 39800 25968 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 134 nsew signal input
flabel metal2 s 22558 200 22614 800 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
port 135 nsew signal input
flabel metal2 s 29642 39200 29698 39800 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
port 136 nsew signal input
flabel metal2 s 28998 39200 29054 39800 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
port 137 nsew signal input
flabel metal2 s 662 39200 718 39800 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_
port 138 nsew signal input
flabel metal2 s 7102 39200 7158 39800 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_
port 139 nsew signal input
flabel metal2 s 27066 200 27122 800 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_
port 140 nsew signal input
flabel metal3 s 200 10208 800 10328 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_
port 141 nsew signal input
flabel metal3 s 200 35368 800 35488 0 FreeSans 480 0 0 0 vccd1
port 142 nsew signal bidirectional
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 142 nsew signal bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 142 nsew signal bidirectional
flabel metal3 s 39200 18368 39800 18488 0 FreeSans 480 0 0 0 vssd1
port 143 nsew signal bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 143 nsew signal bidirectional
rlabel metal1 19964 37536 19964 37536 0 vccd1
rlabel metal1 19964 36992 19964 36992 0 vssd1
rlabel metal1 22310 10438 22310 10438 0 _0000_
rlabel metal1 16376 14246 16376 14246 0 _0001_
rlabel metal1 7360 12954 7360 12954 0 _0002_
rlabel metal2 21666 4709 21666 4709 0 _0003_
rlabel metal1 21121 4522 21121 4522 0 _0004_
rlabel metal1 30728 3910 30728 3910 0 _0005_
rlabel metal2 31694 2176 31694 2176 0 _0006_
rlabel metal2 22034 5151 22034 5151 0 _0007_
rlabel metal2 6578 5916 6578 5916 0 _0008_
rlabel metal1 6578 6154 6578 6154 0 _0009_
rlabel metal1 12528 7446 12528 7446 0 _0010_
rlabel metal1 13846 6732 13846 6732 0 _0011_
rlabel metal2 12742 6018 12742 6018 0 _0012_
rlabel metal2 12466 7548 12466 7548 0 _0013_
rlabel metal1 8326 11526 8326 11526 0 _0014_
rlabel metal1 4600 7242 4600 7242 0 _0015_
rlabel metal1 17572 7174 17572 7174 0 _0016_
rlabel metal1 8951 7310 8951 7310 0 _0017_
rlabel metal1 6256 15878 6256 15878 0 _0018_
rlabel metal1 11546 10778 11546 10778 0 _0019_
rlabel metal2 14858 11594 14858 11594 0 _0020_
rlabel metal1 16468 14790 16468 14790 0 _0021_
rlabel metal1 21167 8874 21167 8874 0 _0022_
rlabel metal2 15134 3859 15134 3859 0 _0023_
rlabel metal2 13386 3638 13386 3638 0 _0024_
rlabel metal1 2898 3910 2898 3910 0 _0025_
rlabel metal2 7958 4981 7958 4981 0 _0026_
rlabel metal2 8602 3213 8602 3213 0 _0027_
rlabel metal1 20838 3543 20838 3543 0 _0028_
rlabel metal1 13754 9384 13754 9384 0 _0029_
rlabel metal2 11914 15113 11914 15113 0 _0030_
rlabel metal1 5290 13192 5290 13192 0 _0031_
rlabel metal2 7544 12580 7544 12580 0 _0032_
rlabel metal1 7728 12614 7728 12614 0 _0033_
rlabel metal2 13570 7327 13570 7327 0 _0034_
rlabel metal1 18538 7895 18538 7895 0 _0035_
rlabel metal1 16429 7786 16429 7786 0 _0036_
rlabel metal2 15318 8126 15318 8126 0 _0037_
rlabel metal2 4370 6817 4370 6817 0 _0038_
rlabel metal1 4784 5542 4784 5542 0 _0039_
rlabel via2 12374 8517 12374 8517 0 _0040_
rlabel metal2 29762 2669 29762 2669 0 _0041_
rlabel metal1 18821 3094 18821 3094 0 _0042_
rlabel metal1 20838 2523 20838 2523 0 _0043_
rlabel metal1 24019 4522 24019 4522 0 _0044_
rlabel metal2 22034 6069 22034 6069 0 _0045_
rlabel metal1 20378 6392 20378 6392 0 _0046_
rlabel metal1 10534 2958 10534 2958 0 _0047_
rlabel metal1 9522 5032 9522 5032 0 _0048_
rlabel metal1 4784 4454 4784 4454 0 _0049_
rlabel metal1 2162 4012 2162 4012 0 _0050_
rlabel metal1 28290 4182 28290 4182 0 _0051_
rlabel metal1 20654 2951 20654 2951 0 _0052_
rlabel metal1 19550 14246 19550 14246 0 _0053_
rlabel metal1 18584 14246 18584 14246 0 _0054_
rlabel metal2 20010 11424 20010 11424 0 _0055_
rlabel metal1 4922 15334 4922 15334 0 _0056_
rlabel metal1 3542 7378 3542 7378 0 _0057_
rlabel metal1 13938 6324 13938 6324 0 _0058_
rlabel metal1 18538 14790 18538 14790 0 _0059_
rlabel metal1 17894 14246 17894 14246 0 _0060_
rlabel metal1 6072 14314 6072 14314 0 _0061_
rlabel metal1 11454 10642 11454 10642 0 _0062_
rlabel metal2 22034 7310 22034 7310 0 _0063_
rlabel metal2 21022 8296 21022 8296 0 _0064_
rlabel metal1 20102 12920 20102 12920 0 _0065_
rlabel metal1 21788 12138 21788 12138 0 _0066_
rlabel metal1 21466 9554 21466 9554 0 _0067_
rlabel metal1 22409 12886 22409 12886 0 _0068_
rlabel metal1 7951 12886 7951 12886 0 _0069_
rlabel metal1 21620 15334 21620 15334 0 _0070_
rlabel metal1 21206 8432 21206 8432 0 _0071_
rlabel metal1 14398 11832 14398 11832 0 _0072_
rlabel metal2 18906 7174 18906 7174 0 _0073_
rlabel metal2 21390 5780 21390 5780 0 _0074_
rlabel metal1 21206 13940 21206 13940 0 _0075_
rlabel metal1 22908 9146 22908 9146 0 _0076_
rlabel metal1 3128 9486 3128 9486 0 _0077_
rlabel metal2 5842 6936 5842 6936 0 _0078_
rlabel metal2 23874 4063 23874 4063 0 _0079_
rlabel metal2 12466 5185 12466 5185 0 _0080_
rlabel metal1 4830 9418 4830 9418 0 _0081_
rlabel metal1 5803 2346 5803 2346 0 _0082_
rlabel metal2 12558 4233 12558 4233 0 _0083_
rlabel metal2 8326 14773 8326 14773 0 _0084_
rlabel via2 13110 9605 13110 9605 0 _0085_
rlabel metal1 14529 12886 14529 12886 0 _0086_
rlabel metal1 17848 15878 17848 15878 0 _0087_
rlabel metal2 9890 6936 9890 6936 0 _0088_
rlabel metal1 2415 9962 2415 9962 0 _0089_
rlabel metal1 4462 10098 4462 10098 0 _0090_
rlabel metal2 6118 6494 6118 6494 0 _0091_
rlabel metal1 4646 4726 4646 4726 0 _0092_
rlabel metal1 10718 13362 10718 13362 0 _0093_
rlabel metal1 9768 13226 9768 13226 0 _0094_
rlabel metal1 6946 13226 6946 13226 0 _0095_
rlabel metal1 13156 10778 13156 10778 0 _0096_
rlabel metal2 20746 4284 20746 4284 0 _0097_
rlabel metal2 12650 4148 12650 4148 0 _0098_
rlabel metal1 19327 5610 19327 5610 0 _0099_
rlabel metal1 26772 5882 26772 5882 0 _0100_
rlabel metal2 6946 14144 6946 14144 0 _0101_
rlabel metal1 15594 9350 15594 9350 0 _0102_
rlabel metal1 12190 4488 12190 4488 0 _0103_
rlabel metal1 5474 2074 5474 2074 0 _0104_
rlabel metal1 5336 15334 5336 15334 0 _0105_
rlabel metal1 5198 7242 5198 7242 0 _0106_
rlabel metal1 5520 8058 5520 8058 0 _0107_
rlabel metal1 3910 14790 3910 14790 0 _0108_
rlabel metal1 6394 12750 6394 12750 0 _0109_
rlabel metal2 12742 9690 12742 9690 0 _0110_
rlabel metal1 5244 13838 5244 13838 0 _0111_
rlabel metal1 5290 6834 5290 6834 0 _0112_
rlabel metal2 15318 2176 15318 2176 0 _0113_
rlabel metal1 6946 2278 6946 2278 0 _0114_
rlabel metal1 12574 2346 12574 2346 0 _0115_
rlabel metal1 3634 8840 3634 8840 0 _0116_
rlabel metal1 9430 12648 9430 12648 0 _0117_
rlabel metal1 2622 4658 2622 4658 0 _0118_
rlabel metal1 5244 7854 5244 7854 0 _0119_
rlabel metal2 15318 15028 15318 15028 0 _0120_
rlabel metal1 14490 14314 14490 14314 0 _0121_
rlabel metal1 16698 7378 16698 7378 0 _0122_
rlabel metal1 2622 7820 2622 7820 0 _0123_
rlabel metal2 12558 13447 12558 13447 0 _0124_
rlabel metal2 21390 13124 21390 13124 0 _0125_
rlabel metal2 4922 14926 4922 14926 0 _0126_
rlabel metal1 23966 8466 23966 8466 0 _0127_
rlabel metal1 30958 16048 30958 16048 0 _0128_
rlabel metal2 28658 19652 28658 19652 0 _0129_
rlabel metal2 3266 7378 3266 7378 0 _0130_
rlabel metal1 2162 15674 2162 15674 0 _0131_
rlabel metal1 24794 21590 24794 21590 0 _0132_
rlabel metal1 29854 18394 29854 18394 0 _0133_
rlabel metal1 17158 18598 17158 18598 0 _0134_
rlabel metal2 29946 15674 29946 15674 0 _0135_
rlabel metal2 26266 15164 26266 15164 0 _0136_
rlabel metal1 31602 9520 31602 9520 0 _0137_
rlabel metal2 14030 26486 14030 26486 0 _0138_
rlabel metal2 10074 26758 10074 26758 0 _0139_
rlabel metal1 15042 26554 15042 26554 0 _0140_
rlabel metal1 17664 19482 17664 19482 0 _0141_
rlabel metal2 29486 10812 29486 10812 0 _0142_
rlabel metal2 29946 14042 29946 14042 0 _0143_
rlabel metal2 22494 25738 22494 25738 0 _0144_
rlabel metal1 25484 20026 25484 20026 0 _0145_
rlabel metal1 23322 26996 23322 26996 0 _0146_
rlabel metal1 23460 19346 23460 19346 0 _0147_
rlabel metal2 30498 12036 30498 12036 0 _0148_
rlabel metal2 31510 14348 31510 14348 0 _0149_
rlabel metal2 10350 28356 10350 28356 0 _0150_
rlabel metal1 10810 27574 10810 27574 0 _0151_
rlabel metal2 13018 27166 13018 27166 0 _0152_
rlabel metal2 27554 18938 27554 18938 0 _0153_
rlabel metal1 24794 24786 24794 24786 0 _0154_
rlabel metal1 21482 26316 21482 26316 0 _0155_
rlabel metal1 15180 14994 15180 14994 0 _0156_
rlabel metal1 2484 9554 2484 9554 0 _0157_
rlabel metal1 2300 10030 2300 10030 0 _0158_
rlabel metal2 14674 16218 14674 16218 0 _0159_
rlabel metal2 10994 15742 10994 15742 0 _0160_
rlabel metal1 27094 7786 27094 7786 0 _0161_
rlabel metal2 19550 25704 19550 25704 0 _0162_
rlabel metal1 13800 24854 13800 24854 0 _0163_
rlabel metal2 10350 23800 10350 23800 0 _0164_
rlabel metal2 21298 25432 21298 25432 0 _0165_
rlabel metal2 17250 23902 17250 23902 0 _0166_
rlabel metal2 10810 25704 10810 25704 0 _0167_
rlabel metal2 20562 14756 20562 14756 0 _0168_
rlabel metal1 21252 17850 21252 17850 0 _0169_
rlabel metal2 21850 13736 21850 13736 0 _0170_
rlabel metal1 7084 15062 7084 15062 0 _0171_
rlabel metal2 18538 14280 18538 14280 0 _0172_
rlabel metal2 7682 15640 7682 15640 0 _0173_
rlabel metal1 8096 19754 8096 19754 0 _0174_
rlabel metal1 16192 23766 16192 23766 0 _0175_
rlabel metal1 16376 17306 16376 17306 0 _0176_
rlabel metal1 8878 20502 8878 20502 0 _0177_
rlabel metal2 12374 21896 12374 21896 0 _0178_
rlabel metal1 14812 18326 14812 18326 0 _0179_
rlabel metal1 8878 15402 8878 15402 0 _0180_
rlabel metal1 15134 24854 15134 24854 0 _0181_
rlabel metal1 17940 24854 17940 24854 0 _0182_
rlabel metal2 22402 12002 22402 12002 0 _0183_
rlabel metal2 22586 4692 22586 4692 0 _0184_
rlabel metal2 26358 14144 26358 14144 0 _0185_
rlabel metal2 17618 15470 17618 15470 0 _0186_
rlabel metal1 17480 18938 17480 18938 0 _0187_
rlabel metal2 12558 19040 12558 19040 0 _0188_
rlabel metal1 25070 3094 25070 3094 0 _0189_
rlabel metal2 12282 18190 12282 18190 0 _0190_
rlabel metal1 25070 18666 25070 18666 0 _0191_
rlabel metal2 23690 9384 23690 9384 0 _0192_
rlabel metal2 2990 5848 2990 5848 0 _0193_
rlabel metal1 26772 2006 26772 2006 0 _0194_
rlabel metal1 8372 18938 8372 18938 0 _0195_
rlabel metal1 9844 17782 9844 17782 0 _0196_
rlabel metal1 7268 20570 7268 20570 0 _0197_
rlabel metal1 22862 24072 22862 24072 0 _0198_
rlabel metal2 23414 23528 23414 23528 0 _0199_
rlabel metal1 21390 19720 21390 19720 0 _0200_
rlabel metal2 12650 24344 12650 24344 0 _0201_
rlabel metal1 13938 22678 13938 22678 0 _0202_
rlabel metal2 7498 21726 7498 21726 0 _0203_
rlabel metal2 7866 19176 7866 19176 0 _0204_
rlabel metal2 5106 19618 5106 19618 0 _0205_
rlabel metal2 5474 18462 5474 18462 0 _0206_
rlabel metal1 20562 15368 20562 15368 0 _0207_
rlabel metal2 23322 4590 23322 4590 0 _0208_
rlabel metal1 25576 10778 25576 10778 0 _0209_
rlabel metal2 13110 14110 13110 14110 0 _0210_
rlabel metal2 19918 20196 19918 20196 0 _0211_
rlabel metal1 11454 17544 11454 17544 0 _0212_
rlabel metal1 25760 14042 25760 14042 0 _0213_
rlabel metal2 25990 18088 25990 18088 0 _0214_
rlabel metal2 4278 17374 4278 17374 0 _0215_
rlabel metal1 23230 10234 23230 10234 0 _0216_
rlabel metal2 15318 19992 15318 19992 0 _0217_
rlabel metal1 21666 10200 21666 10200 0 _0218_
rlabel metal2 25070 8738 25070 8738 0 _0219_
rlabel metal1 24748 8058 24748 8058 0 _0220_
rlabel metal2 29302 4828 29302 4828 0 _0221_
rlabel metal2 8418 20366 8418 20366 0 _0222_
rlabel metal1 15640 21590 15640 21590 0 _0223_
rlabel metal1 24978 7990 24978 7990 0 _0224_
rlabel metal2 12926 18088 12926 18088 0 _0225_
rlabel metal1 14582 20570 14582 20570 0 _0226_
rlabel metal2 27554 6120 27554 6120 0 _0227_
rlabel metal2 30498 4267 30498 4267 0 _0228_
rlabel metal2 7958 17816 7958 17816 0 _0229_
rlabel metal1 23920 6358 23920 6358 0 _0230_
rlabel metal2 9890 13974 9890 13974 0 _0231_
rlabel metal1 14030 15062 14030 15062 0 _0232_
rlabel metal1 9062 16150 9062 16150 0 _0233_
rlabel metal2 14490 16626 14490 16626 0 _0234_
rlabel metal1 14858 18632 14858 18632 0 _0235_
rlabel metal1 21482 17136 21482 17136 0 _0236_
rlabel metal1 9798 16490 9798 16490 0 _0237_
rlabel metal1 24656 13226 24656 13226 0 _0238_
rlabel metal2 13478 16558 13478 16558 0 _0239_
rlabel metal1 23874 16762 23874 16762 0 _0240_
rlabel metal2 20102 16558 20102 16558 0 _0241_
rlabel metal2 23138 6120 23138 6120 0 _0242_
rlabel metal2 12834 19822 12834 19822 0 _0243_
rlabel metal2 13294 19992 13294 19992 0 _0244_
rlabel metal1 17756 21930 17756 21930 0 _0245_
rlabel metal1 19642 21624 19642 21624 0 _0246_
rlabel metal1 22172 22746 22172 22746 0 _0247_
rlabel metal2 25070 22882 25070 22882 0 _0248_
rlabel metal1 10120 17238 10120 17238 0 _0249_
rlabel metal1 26450 18666 26450 18666 0 _0250_
rlabel metal2 9982 20400 9982 20400 0 _0251_
rlabel metal2 20470 21080 20470 21080 0 _0252_
rlabel metal2 23598 21726 23598 21726 0 _0253_
rlabel metal1 26864 22202 26864 22202 0 _0254_
rlabel metal1 28198 2550 28198 2550 0 _0255_
rlabel metal2 28934 3706 28934 3706 0 _0256_
rlabel metal2 9798 16609 9798 16609 0 _0257_
rlabel metal2 24702 15198 24702 15198 0 _0258_
rlabel metal2 7130 17544 7130 17544 0 _0259_
rlabel metal1 26484 6698 26484 6698 0 _0260_
rlabel metal1 11546 16150 11546 16150 0 _0261_
rlabel metal1 24978 4182 24978 4182 0 _0262_
rlabel metal2 27554 4590 27554 4590 0 _0263_
rlabel metal1 25070 6664 25070 6664 0 _0264_
rlabel metal1 26956 5270 26956 5270 0 _0265_
rlabel metal1 25254 7446 25254 7446 0 _0266_
rlabel metal2 12466 19074 12466 19074 0 _0267_
rlabel metal1 11224 18326 11224 18326 0 _0268_
rlabel metal1 11776 23494 11776 23494 0 _0269_
rlabel metal2 9890 23086 9890 23086 0 _0270_
rlabel metal2 14858 23256 14858 23256 0 _0271_
rlabel metal2 13018 23256 13018 23256 0 _0272_
rlabel metal1 16698 20808 16698 20808 0 _0273_
rlabel metal1 10580 22406 10580 22406 0 _0274_
rlabel metal2 13110 19176 13110 19176 0 _0275_
rlabel metal2 10810 20264 10810 20264 0 _0276_
rlabel metal1 7820 22474 7820 22474 0 _0277_
rlabel metal2 17710 21046 17710 21046 0 _0278_
rlabel metal2 15042 15062 15042 15062 0 _0279_
rlabel metal2 19550 15385 19550 15385 0 _0280_
rlabel metal2 22310 16864 22310 16864 0 _0281_
rlabel metal1 4646 20808 4646 20808 0 _0282_
rlabel metal1 15180 18122 15180 18122 0 _0283_
rlabel metal2 23690 17170 23690 17170 0 _0284_
rlabel metal1 17112 16762 17112 16762 0 _0285_
rlabel metal1 4508 17850 4508 17850 0 _0286_
rlabel metal1 25300 11050 25300 11050 0 _0287_
rlabel metal2 25990 3672 25990 3672 0 _0288_
rlabel via2 30406 3077 30406 3077 0 _0289_
rlabel metal2 24334 13566 24334 13566 0 _0290_
rlabel metal1 24794 3400 24794 3400 0 _0291_
rlabel metal1 21390 14042 21390 14042 0 _0292_
rlabel metal2 22770 3502 22770 3502 0 _0293_
rlabel metal1 23322 13192 23322 13192 0 _0294_
rlabel metal2 20654 19108 20654 19108 0 _0295_
rlabel metal1 22034 16150 22034 16150 0 _0296_
rlabel metal1 18814 16762 18814 16762 0 _0297_
rlabel metal1 14030 18394 14030 18394 0 _0298_
rlabel metal2 27462 3298 27462 3298 0 _0299_
rlabel metal2 24794 12036 24794 12036 0 _0300_
rlabel metal1 19826 16490 19826 16490 0 _0301_
rlabel metal1 27048 4998 27048 4998 0 _0302_
rlabel metal1 18630 18394 18630 18394 0 _0303_
rlabel metal1 21206 22950 21206 22950 0 _0304_
rlabel metal1 8464 14586 8464 14586 0 _0305_
rlabel metal1 16012 15878 16012 15878 0 _0306_
rlabel metal1 18262 18394 18262 18394 0 _0307_
rlabel metal1 19136 14042 19136 14042 0 _0308_
rlabel metal2 22954 24718 22954 24718 0 _0309_
rlabel metal1 20332 23698 20332 23698 0 _0310_
rlabel metal1 26726 18938 26726 18938 0 _0311_
rlabel metal1 26680 22406 26680 22406 0 _0312_
rlabel metal2 18814 23868 18814 23868 0 _0313_
rlabel metal1 26634 20366 26634 20366 0 _0314_
rlabel metal2 12098 27438 12098 27438 0 _0315_
rlabel metal2 13294 26588 13294 26588 0 _0316_
rlabel metal1 11776 26962 11776 26962 0 _0317_
rlabel metal1 12880 27506 12880 27506 0 _0318_
rlabel metal1 11960 24786 11960 24786 0 _0319_
rlabel metal2 11914 27676 11914 27676 0 _0320_
rlabel metal2 29486 11934 29486 11934 0 _0321_
rlabel metal1 31096 12818 31096 12818 0 _0322_
rlabel metal2 23046 19992 23046 19992 0 _0323_
rlabel metal2 27922 11560 27922 11560 0 _0324_
rlabel metal2 29210 13124 29210 13124 0 _0325_
rlabel metal2 21390 19924 21390 19924 0 _0326_
rlabel metal1 24840 20434 24840 20434 0 _0327_
rlabel metal1 23230 26758 23230 26758 0 _0328_
rlabel metal2 24794 24684 24794 24684 0 _0329_
rlabel metal2 24702 19652 24702 19652 0 _0330_
rlabel metal1 22172 24922 22172 24922 0 _0331_
rlabel metal1 17020 23154 17020 23154 0 _0332_
rlabel metal2 29302 10948 29302 10948 0 _0333_
rlabel metal2 29762 13668 29762 13668 0 _0334_
rlabel metal2 17066 19006 17066 19006 0 _0335_
rlabel metal1 28336 12410 28336 12410 0 _0336_
rlabel metal1 27416 13362 27416 13362 0 _0337_
rlabel metal1 28658 18326 28658 18326 0 _0338_
rlabel metal2 12834 26622 12834 26622 0 _0339_
rlabel metal1 15042 25874 15042 25874 0 _0340_
rlabel metal2 14582 25500 14582 25500 0 _0341_
rlabel metal2 12190 25466 12190 25466 0 _0342_
rlabel metal1 16008 26418 16008 26418 0 _0343_
rlabel metal2 14766 23902 14766 23902 0 _0344_
rlabel metal2 29486 8908 29486 8908 0 _0345_
rlabel metal2 26082 15300 26082 15300 0 _0346_
rlabel metal1 30452 9010 30452 9010 0 _0347_
rlabel metal1 26174 12750 26174 12750 0 _0348_
rlabel metal1 28842 14994 28842 14994 0 _0349_
rlabel via1 15318 17595 15318 17595 0 _0350_
rlabel metal1 27324 13906 27324 13906 0 _0351_
rlabel metal2 15686 16830 15686 16830 0 _0352_
rlabel metal1 28566 17170 28566 17170 0 _0353_
rlabel metal1 25162 18258 25162 18258 0 _0354_
rlabel metal1 29532 18802 29532 18802 0 _0355_
rlabel metal1 17664 19346 17664 19346 0 _0356_
rlabel metal2 2622 15436 2622 15436 0 _0357_
rlabel metal2 2898 7820 2898 7820 0 _0358_
rlabel metal2 2714 14620 2714 14620 0 _0359_
rlabel metal1 1932 5338 1932 5338 0 _0360_
rlabel metal2 29946 18088 29946 18088 0 _0361_
rlabel metal1 29164 15538 29164 15538 0 _0362_
rlabel metal2 28566 17272 28566 17272 0 _0363_
rlabel metal2 28566 15844 28566 15844 0 _0364_
rlabel metal3 1234 19108 1234 19108 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
rlabel metal3 1234 7548 1234 7548 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
rlabel metal1 5336 37230 5336 37230 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal3 1142 5508 1142 5508 0 bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 35466 1894 35466 1894 0 bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 31970 3196 31970 3196 0 bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal3 1234 22508 1234 22508 0 bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal3 1050 6868 1050 6868 0 bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_
rlabel metal1 18216 37230 18216 37230 0 bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal3 1786 38828 1786 38828 0 bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_
rlabel metal2 5106 5508 5106 5508 0 ccff_head
rlabel metal2 29026 1520 29026 1520 0 ccff_tail
rlabel metal1 25944 37230 25944 37230 0 chanx_left_in[0]
rlabel metal1 6302 37230 6302 37230 0 chanx_left_in[10]
rlabel metal1 31878 3468 31878 3468 0 chanx_left_in[11]
rlabel metal1 9200 36754 9200 36754 0 chanx_left_in[12]
rlabel metal1 16698 3434 16698 3434 0 chanx_left_in[13]
rlabel metal3 1234 17068 1234 17068 0 chanx_left_in[14]
rlabel metal3 1280 2108 1280 2108 0 chanx_left_in[15]
rlabel metal1 27922 37230 27922 37230 0 chanx_left_in[16]
rlabel metal2 11638 1761 11638 1761 0 chanx_left_in[17]
rlabel metal2 38318 32215 38318 32215 0 chanx_left_in[18]
rlabel metal2 38318 27353 38318 27353 0 chanx_left_in[1]
rlabel metal2 9706 2370 9706 2370 0 chanx_left_in[2]
rlabel metal3 1211 748 1211 748 0 chanx_left_in[3]
rlabel via2 38318 8925 38318 8925 0 chanx_left_in[4]
rlabel metal2 15180 37230 15180 37230 0 chanx_left_in[5]
rlabel via2 38318 30685 38318 30685 0 chanx_left_in[6]
rlabel metal2 38318 28883 38318 28883 0 chanx_left_in[7]
rlabel metal1 32384 37230 32384 37230 0 chanx_left_in[8]
rlabel metal2 18078 1418 18078 1418 0 chanx_left_in[9]
rlabel metal1 36248 37094 36248 37094 0 chanx_left_out[0]
rlabel metal2 38226 12461 38226 12461 0 chanx_left_out[10]
rlabel metal2 33534 1520 33534 1520 0 chanx_left_out[11]
rlabel metal3 1234 30668 1234 30668 0 chanx_left_out[12]
rlabel metal3 1234 15708 1234 15708 0 chanx_left_out[13]
rlabel metal1 20148 37094 20148 37094 0 chanx_left_out[15]
rlabel via2 38226 35445 38226 35445 0 chanx_left_out[16]
rlabel metal1 36616 2550 36616 2550 0 chanx_left_out[17]
rlabel metal1 19504 36890 19504 36890 0 chanx_left_out[18]
rlabel metal2 34178 1520 34178 1520 0 chanx_left_out[1]
rlabel metal1 31096 37094 31096 37094 0 chanx_left_out[2]
rlabel metal1 34822 37094 34822 37094 0 chanx_left_out[3]
rlabel metal1 36156 36890 36156 36890 0 chanx_left_out[4]
rlabel metal1 16192 37094 16192 37094 0 chanx_left_out[5]
rlabel metal2 38226 11101 38226 11101 0 chanx_left_out[6]
rlabel via2 38226 13685 38226 13685 0 chanx_left_out[7]
rlabel via2 38226 19125 38226 19125 0 chanx_left_out[8]
rlabel metal2 27738 1520 27738 1520 0 chanx_left_out[9]
rlabel metal1 37306 36142 37306 36142 0 chany_bottom_in[0]
rlabel metal2 37490 32793 37490 32793 0 chany_bottom_in[10]
rlabel metal1 24656 37230 24656 37230 0 chany_bottom_in[11]
rlabel metal2 12374 37230 12374 37230 0 chany_bottom_in[12]
rlabel metal2 37490 24021 37490 24021 0 chany_bottom_in[13]
rlabel metal1 8786 37298 8786 37298 0 chany_bottom_in[14]
rlabel metal1 11776 37230 11776 37230 0 chany_bottom_in[15]
rlabel metal1 22632 37298 22632 37298 0 chany_bottom_in[16]
rlabel metal1 2530 11220 2530 11220 0 chany_bottom_in[17]
rlabel metal1 2852 36754 2852 36754 0 chany_bottom_in[18]
rlabel metal2 38134 15215 38134 15215 0 chany_bottom_in[1]
rlabel metal1 3956 37298 3956 37298 0 chany_bottom_in[2]
rlabel metal1 37398 3026 37398 3026 0 chany_bottom_in[3]
rlabel metal3 1234 14348 1234 14348 0 chany_bottom_in[4]
rlabel metal2 37490 7701 37490 7701 0 chany_bottom_in[5]
rlabel metal3 1234 28628 1234 28628 0 chany_bottom_in[6]
rlabel metal2 14582 3961 14582 3961 0 chany_bottom_in[7]
rlabel metal3 1188 21148 1188 21148 0 chany_bottom_in[8]
rlabel metal2 16146 1894 16146 1894 0 chany_bottom_in[9]
rlabel metal3 1234 24548 1234 24548 0 chany_bottom_out[0]
rlabel metal2 33028 37094 33028 37094 0 chany_bottom_out[10]
rlabel metal3 1234 32708 1234 32708 0 chany_bottom_out[11]
rlabel metal2 30314 1520 30314 1520 0 chany_bottom_out[12]
rlabel metal2 38226 25177 38226 25177 0 chany_bottom_out[13]
rlabel via2 38226 5525 38226 5525 0 chany_bottom_out[14]
rlabel metal1 26910 37094 26910 37094 0 chany_bottom_out[15]
rlabel metal2 36846 37128 36846 37128 0 chany_bottom_out[16]
rlabel metal1 37536 36890 37536 36890 0 chany_bottom_out[17]
rlabel metal2 690 1792 690 1792 0 chany_bottom_out[18]
rlabel metal1 5336 3910 5336 3910 0 chany_bottom_out[1]
rlabel metal2 38686 1792 38686 1792 0 chany_bottom_out[2]
rlabel metal3 1234 13668 1234 13668 0 chany_bottom_out[3]
rlabel via2 38226 21845 38226 21845 0 chany_bottom_out[4]
rlabel metal2 38226 15793 38226 15793 0 chany_bottom_out[5]
rlabel metal1 16928 37094 16928 37094 0 chany_bottom_out[6]
rlabel metal2 3266 1520 3266 1520 0 chany_bottom_out[7]
rlabel metal2 38226 3417 38226 3417 0 chany_bottom_out[8]
rlabel via2 38226 17051 38226 17051 0 chany_bottom_out[9]
rlabel metal3 1142 27268 1142 27268 0 chany_top_in[0]
rlabel metal1 2024 37298 2024 37298 0 chany_top_in[10]
rlabel metal3 1188 25908 1188 25908 0 chany_top_in[11]
rlabel metal3 1142 20468 1142 20468 0 chany_top_in[12]
rlabel metal3 1832 39508 1832 39508 0 chany_top_in[13]
rlabel metal1 38088 37298 38088 37298 0 chany_top_in[14]
rlabel metal2 8418 823 8418 823 0 chany_top_in[15]
rlabel metal3 1142 17748 1142 17748 0 chany_top_in[16]
rlabel metal2 23230 1554 23230 1554 0 chany_top_in[17]
rlabel metal2 37398 1588 37398 1588 0 chany_top_in[18]
rlabel metal1 13984 37230 13984 37230 0 chany_top_in[1]
rlabel metal2 33810 3740 33810 3740 0 chany_top_in[2]
rlabel metal1 3864 8466 3864 8466 0 chany_top_in[3]
rlabel metal1 14168 2822 14168 2822 0 chany_top_in[4]
rlabel metal2 38134 4335 38134 4335 0 chany_top_in[5]
rlabel metal2 38134 29427 38134 29427 0 chany_top_in[6]
rlabel via2 38318 20451 38318 20451 0 chany_top_in[7]
rlabel metal2 32246 1588 32246 1588 0 chany_top_in[8]
rlabel metal3 1142 23868 1142 23868 0 chany_top_in[9]
rlabel metal2 38226 10353 38226 10353 0 chany_top_out[0]
rlabel metal3 1234 32028 1234 32028 0 chany_top_out[10]
rlabel via2 38226 22491 38226 22491 0 chany_top_out[11]
rlabel metal2 38226 34221 38226 34221 0 chany_top_out[12]
rlabel metal2 36754 1520 36754 1520 0 chany_top_out[13]
rlabel metal2 38226 36057 38226 36057 0 chany_top_out[14]
rlabel metal3 1234 12308 1234 12308 0 chany_top_out[15]
rlabel metal3 1234 34068 1234 34068 0 chany_top_out[16]
rlabel metal3 1234 3468 1234 3468 0 chany_top_out[17]
rlabel metal2 46 1656 46 1656 0 chany_top_out[18]
rlabel metal3 1234 4148 1234 4148 0 chany_top_out[1]
rlabel metal2 1794 36907 1794 36907 0 chany_top_out[2]
rlabel metal1 10488 37094 10488 37094 0 chany_top_out[3]
rlabel metal1 23368 36890 23368 36890 0 chany_top_out[4]
rlabel metal3 1234 29308 1234 29308 0 chany_top_out[5]
rlabel metal1 6624 2822 6624 2822 0 chany_top_out[6]
rlabel metal2 1978 1520 1978 1520 0 chany_top_out[7]
rlabel metal3 1234 8908 1234 8908 0 chany_top_out[8]
rlabel metal1 21344 37094 21344 37094 0 chany_top_out[9]
rlabel metal1 13478 7854 13478 7854 0 clknet_0_prog_clk
rlabel metal1 6900 2482 6900 2482 0 clknet_4_0_0_prog_clk
rlabel metal1 17020 4590 17020 4590 0 clknet_4_10_0_prog_clk
rlabel metal2 20010 7684 20010 7684 0 clknet_4_11_0_prog_clk
rlabel metal2 15502 9826 15502 9826 0 clknet_4_12_0_prog_clk
rlabel metal1 15364 11662 15364 11662 0 clknet_4_13_0_prog_clk
rlabel metal1 17112 9554 17112 9554 0 clknet_4_14_0_prog_clk
rlabel metal1 16744 12750 16744 12750 0 clknet_4_15_0_prog_clk
rlabel metal1 6532 7922 6532 7922 0 clknet_4_1_0_prog_clk
rlabel metal1 8602 2482 8602 2482 0 clknet_4_2_0_prog_clk
rlabel metal1 11914 5678 11914 5678 0 clknet_4_3_0_prog_clk
rlabel metal2 6854 8772 6854 8772 0 clknet_4_4_0_prog_clk
rlabel metal2 9200 13362 9200 13362 0 clknet_4_5_0_prog_clk
rlabel metal1 8878 7922 8878 7922 0 clknet_4_6_0_prog_clk
rlabel metal1 7958 11798 7958 11798 0 clknet_4_7_0_prog_clk
rlabel metal1 13800 3434 13800 3434 0 clknet_4_8_0_prog_clk
rlabel metal1 15410 7922 15410 7922 0 clknet_4_9_0_prog_clk
rlabel metal2 19366 1639 19366 1639 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel metal2 35466 37988 35466 37988 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal3 38786 6868 38786 6868 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
rlabel metal3 1234 36108 1234 36108 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
rlabel metal3 7866 12444 7866 12444 0 mem_bottom_track_1.DFFR_0_.D
rlabel metal2 5842 17765 5842 17765 0 mem_bottom_track_1.DFFR_0_.Q
rlabel metal1 13432 11526 13432 11526 0 mem_bottom_track_1.DFFR_1_.Q
rlabel metal1 14168 21998 14168 21998 0 mem_bottom_track_1.DFFR_2_.Q
rlabel metal2 13570 19125 13570 19125 0 mem_bottom_track_1.DFFR_3_.Q
rlabel metal1 9200 12954 9200 12954 0 mem_bottom_track_1.DFFR_4_.Q
rlabel metal2 9476 15572 9476 15572 0 mem_bottom_track_1.DFFR_5_.Q
rlabel metal1 9338 17612 9338 17612 0 mem_bottom_track_1.DFFR_6_.Q
rlabel metal2 11362 14620 11362 14620 0 mem_bottom_track_1.DFFR_7_.Q
rlabel metal2 16330 2210 16330 2210 0 mem_bottom_track_17.DFFR_0_.D
rlabel metal1 13984 7514 13984 7514 0 mem_bottom_track_17.DFFR_0_.Q
rlabel metal1 11592 19822 11592 19822 0 mem_bottom_track_17.DFFR_1_.Q
rlabel metal2 14306 20383 14306 20383 0 mem_bottom_track_17.DFFR_2_.Q
rlabel metal1 18354 2482 18354 2482 0 mem_bottom_track_17.DFFR_3_.Q
rlabel metal1 23598 2958 23598 2958 0 mem_bottom_track_17.DFFR_4_.Q
rlabel metal1 21850 4726 21850 4726 0 mem_bottom_track_17.DFFR_5_.Q
rlabel metal2 21298 4930 21298 4930 0 mem_bottom_track_17.DFFR_6_.Q
rlabel metal1 29762 5236 29762 5236 0 mem_bottom_track_17.DFFR_7_.Q
rlabel via2 18906 4165 18906 4165 0 mem_bottom_track_25.DFFR_0_.Q
rlabel metal1 8556 17646 8556 17646 0 mem_bottom_track_25.DFFR_1_.Q
rlabel metal1 25438 15606 25438 15606 0 mem_bottom_track_25.DFFR_2_.Q
rlabel metal1 14536 3434 14536 3434 0 mem_bottom_track_25.DFFR_3_.Q
rlabel metal2 16054 4471 16054 4471 0 mem_bottom_track_25.DFFR_4_.Q
rlabel metal2 19550 4947 19550 4947 0 mem_bottom_track_25.DFFR_5_.Q
rlabel metal1 12558 20808 12558 20808 0 mem_bottom_track_33.DFFR_0_.Q
rlabel metal1 14766 23698 14766 23698 0 mem_bottom_track_33.DFFR_1_.Q
rlabel metal2 8004 16660 8004 16660 0 mem_bottom_track_33.DFFR_2_.Q
rlabel metal1 12650 13736 12650 13736 0 mem_bottom_track_33.DFFR_3_.Q
rlabel metal1 14444 8874 14444 8874 0 mem_bottom_track_33.DFFR_4_.Q
rlabel metal2 13202 15997 13202 15997 0 mem_bottom_track_33.DFFR_5_.Q
rlabel metal1 15502 19346 15502 19346 0 mem_bottom_track_9.DFFR_0_.Q
rlabel via2 19734 13243 19734 13243 0 mem_bottom_track_9.DFFR_1_.Q
rlabel metal1 19826 19890 19826 19890 0 mem_bottom_track_9.DFFR_2_.Q
rlabel metal3 8832 12580 8832 12580 0 mem_bottom_track_9.DFFR_3_.Q
rlabel metal2 18262 7905 18262 7905 0 mem_bottom_track_9.DFFR_4_.Q
rlabel metal2 18722 2329 18722 2329 0 mem_bottom_track_9.DFFR_5_.Q
rlabel metal1 15180 2482 15180 2482 0 mem_bottom_track_9.DFFR_6_.Q
rlabel metal3 18975 18020 18975 18020 0 mem_left_track_1.DFFR_0_.Q
rlabel metal1 7774 14994 7774 14994 0 mem_left_track_1.DFFR_1_.Q
rlabel metal2 14260 12716 14260 12716 0 mem_left_track_1.DFFR_2_.Q
rlabel metal1 16882 16558 16882 16558 0 mem_left_track_1.DFFR_3_.Q
rlabel metal1 17940 7922 17940 7922 0 mem_left_track_1.DFFR_4_.Q
rlabel metal2 19136 17238 19136 17238 0 mem_left_track_1.DFFR_5_.Q
rlabel metal1 26174 22576 26174 22576 0 mem_left_track_11.DFFR_0_.D
rlabel metal2 12604 17238 12604 17238 0 mem_left_track_11.DFFR_0_.Q
rlabel metal1 13386 11730 13386 11730 0 mem_left_track_11.DFFR_1_.Q
rlabel metal1 19458 11832 19458 11832 0 mem_left_track_13.DFFR_0_.Q
rlabel metal1 20194 7310 20194 7310 0 mem_left_track_13.DFFR_1_.Q
rlabel metal1 14674 17646 14674 17646 0 mem_left_track_15.DFFR_0_.Q
rlabel metal1 20148 9962 20148 9962 0 mem_left_track_15.DFFR_1_.Q
rlabel metal1 17250 19312 17250 19312 0 mem_left_track_17.DFFR_0_.Q
rlabel metal1 20470 14042 20470 14042 0 mem_left_track_17.DFFR_1_.Q
rlabel metal2 21758 16014 21758 16014 0 mem_left_track_19.DFFR_0_.Q
rlabel metal2 21574 11730 21574 11730 0 mem_left_track_19.DFFR_1_.Q
rlabel metal1 21482 13770 21482 13770 0 mem_left_track_21.DFFR_0_.Q
rlabel metal1 20056 12750 20056 12750 0 mem_left_track_21.DFFR_1_.Q
rlabel metal1 18078 19380 18078 19380 0 mem_left_track_23.DFFR_0_.Q
rlabel metal1 21022 11696 21022 11696 0 mem_left_track_23.DFFR_1_.Q
rlabel metal2 13156 19516 13156 19516 0 mem_left_track_25.DFFR_0_.Q
rlabel metal1 9614 12614 9614 12614 0 mem_left_track_25.DFFR_1_.Q
rlabel metal1 2208 5678 2208 5678 0 mem_left_track_27.DFFR_0_.Q
rlabel metal1 1748 14994 1748 14994 0 mem_left_track_27.DFFR_1_.Q
rlabel metal1 21114 13872 21114 13872 0 mem_left_track_3.DFFR_0_.Q
rlabel metal1 21574 6154 21574 6154 0 mem_left_track_3.DFFR_1_.Q
rlabel metal1 22126 3502 22126 3502 0 mem_left_track_3.DFFR_2_.Q
rlabel metal1 20194 2278 20194 2278 0 mem_left_track_3.DFFR_3_.Q
rlabel metal1 19458 2822 19458 2822 0 mem_left_track_3.DFFR_4_.Q
rlabel metal1 32062 2924 32062 2924 0 mem_left_track_3.DFFR_5_.Q
rlabel metal1 20240 5610 20240 5610 0 mem_left_track_37.DFFR_0_.Q
rlabel metal1 21436 2822 21436 2822 0 mem_left_track_5.DFFR_0_.Q
rlabel metal1 20424 18734 20424 18734 0 mem_left_track_5.DFFR_1_.Q
rlabel metal2 31878 4420 31878 4420 0 mem_left_track_5.DFFR_2_.Q
rlabel metal2 14766 12852 14766 12852 0 mem_left_track_5.DFFR_3_.Q
rlabel metal1 16882 16490 16882 16490 0 mem_left_track_5.DFFR_4_.Q
rlabel metal2 16468 15538 16468 15538 0 mem_left_track_5.DFFR_5_.Q
rlabel metal1 16560 13838 16560 13838 0 mem_left_track_7.DFFR_0_.Q
rlabel metal1 7491 9146 7491 9146 0 mem_left_track_7.DFFR_1_.Q
rlabel metal3 14743 15300 14743 15300 0 mem_left_track_7.DFFR_2_.Q
rlabel metal1 17664 11186 17664 11186 0 mem_left_track_7.DFFR_3_.Q
rlabel metal1 18768 18258 18768 18258 0 mem_left_track_7.DFFR_4_.Q
rlabel metal1 20194 17612 20194 17612 0 mem_left_track_7.DFFR_5_.Q
rlabel metal1 24794 23528 24794 23528 0 mem_left_track_9.DFFR_0_.Q
rlabel metal1 21712 13294 21712 13294 0 mem_top_track_0.DFFR_0_.Q
rlabel metal2 19412 19652 19412 19652 0 mem_top_track_0.DFFR_1_.Q
rlabel metal2 16330 15708 16330 15708 0 mem_top_track_0.DFFR_2_.Q
rlabel metal2 14122 9248 14122 9248 0 mem_top_track_0.DFFR_3_.Q
rlabel metal2 20470 14433 20470 14433 0 mem_top_track_0.DFFR_4_.Q
rlabel metal1 13616 3910 13616 3910 0 mem_top_track_0.DFFR_5_.Q
rlabel metal1 7544 16082 7544 16082 0 mem_top_track_0.DFFR_6_.Q
rlabel metal1 17657 6970 17657 6970 0 mem_top_track_0.DFFR_7_.Q
rlabel metal1 17664 16558 17664 16558 0 mem_top_track_16.DFFR_0_.D
rlabel metal1 16192 16762 16192 16762 0 mem_top_track_16.DFFR_0_.Q
rlabel metal1 9246 20910 9246 20910 0 mem_top_track_16.DFFR_1_.Q
rlabel metal2 16882 24004 16882 24004 0 mem_top_track_16.DFFR_2_.Q
rlabel metal2 7498 5321 7498 5321 0 mem_top_track_16.DFFR_3_.Q
rlabel metal1 8602 15538 8602 15538 0 mem_top_track_16.DFFR_4_.Q
rlabel metal1 5106 14994 5106 14994 0 mem_top_track_16.DFFR_5_.Q
rlabel metal1 8970 4012 8970 4012 0 mem_top_track_16.DFFR_6_.Q
rlabel metal1 6716 2346 6716 2346 0 mem_top_track_16.DFFR_7_.Q
rlabel metal2 2346 3468 2346 3468 0 mem_top_track_24.DFFR_0_.Q
rlabel metal1 14950 2278 14950 2278 0 mem_top_track_24.DFFR_1_.Q
rlabel metal1 12351 19346 12351 19346 0 mem_top_track_24.DFFR_2_.Q
rlabel metal2 15732 12716 15732 12716 0 mem_top_track_24.DFFR_3_.Q
rlabel metal1 19458 6630 19458 6630 0 mem_top_track_24.DFFR_4_.Q
rlabel metal1 18952 5746 18952 5746 0 mem_top_track_24.DFFR_5_.Q
rlabel metal1 17342 4488 17342 4488 0 mem_top_track_24.DFFR_6_.Q
rlabel metal1 19780 8874 19780 8874 0 mem_top_track_24.DFFR_7_.Q
rlabel metal1 20792 21522 20792 21522 0 mem_top_track_32.DFFR_0_.Q
rlabel metal1 16054 18190 16054 18190 0 mem_top_track_32.DFFR_1_.Q
rlabel metal1 25024 22610 25024 22610 0 mem_top_track_32.DFFR_2_.Q
rlabel metal1 9062 19822 9062 19822 0 mem_top_track_32.DFFR_3_.Q
rlabel metal1 9844 18258 9844 18258 0 mem_top_track_32.DFFR_4_.Q
rlabel metal1 18216 6834 18216 6834 0 mem_top_track_8.DFFR_0_.Q
rlabel metal1 9982 18734 9982 18734 0 mem_top_track_8.DFFR_1_.Q
rlabel metal1 22494 16524 22494 16524 0 mem_top_track_8.DFFR_2_.Q
rlabel metal1 9154 17238 9154 17238 0 mem_top_track_8.DFFR_3_.Q
rlabel metal1 14674 6834 14674 6834 0 mem_top_track_8.DFFR_4_.Q
rlabel metal1 5566 18190 5566 18190 0 mux_bottom_track_1.INVTX1_0_.out
rlabel metal2 12558 25874 12558 25874 0 mux_bottom_track_1.INVTX1_1_.out
rlabel metal1 15962 21964 15962 21964 0 mux_bottom_track_1.INVTX1_2_.out
rlabel metal1 7360 31110 7360 31110 0 mux_bottom_track_1.INVTX1_3_.out
rlabel metal1 4048 12954 4048 12954 0 mux_bottom_track_1.INVTX1_4_.out
rlabel metal1 23322 24242 23322 24242 0 mux_bottom_track_1.INVTX1_5_.out
rlabel metal1 24748 23154 24748 23154 0 mux_bottom_track_1.INVTX1_6_.out
rlabel metal2 21298 20434 21298 20434 0 mux_bottom_track_1.INVTX1_7_.out
rlabel metal1 23552 30022 23552 30022 0 mux_bottom_track_1.INVTX1_8_.out
rlabel metal1 13800 22542 13800 22542 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 23552 23630 23552 23630 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 7038 19958 7038 19958 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 5888 23698 5888 23698 0 mux_bottom_track_1.out
rlabel metal1 26726 5746 26726 5746 0 mux_bottom_track_17.INVTX1_0_.out
rlabel metal2 15594 17102 15594 17102 0 mux_bottom_track_17.INVTX1_1_.out
rlabel metal1 14398 21590 14398 21590 0 mux_bottom_track_17.INVTX1_2_.out
rlabel metal2 25346 6256 25346 6256 0 mux_bottom_track_17.INVTX1_3_.out
rlabel metal1 6808 18326 6808 18326 0 mux_bottom_track_17.INVTX1_4_.out
rlabel metal1 7176 19754 7176 19754 0 mux_bottom_track_17.INVTX1_5_.out
rlabel metal1 15456 21454 15456 21454 0 mux_bottom_track_17.INVTX1_6_.out
rlabel metal1 23092 6154 23092 6154 0 mux_bottom_track_17.INVTX1_7_.out
rlabel metal1 30728 24582 30728 24582 0 mux_bottom_track_17.INVTX1_8_.out
rlabel metal1 13892 16490 13892 16490 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 17204 21454 17204 21454 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 33005 7378 33005 7378 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 36340 6290 36340 6290 0 mux_bottom_track_17.out
rlabel metal1 22908 12954 22908 12954 0 mux_bottom_track_25.INVTX1_0_.out
rlabel metal2 13754 17595 13754 17595 0 mux_bottom_track_25.INVTX1_1_.out
rlabel metal2 1978 7106 1978 7106 0 mux_bottom_track_25.INVTX1_2_.out
rlabel metal1 25622 5100 25622 5100 0 mux_bottom_track_25.INVTX1_3_.out
rlabel metal2 7038 17612 7038 17612 0 mux_bottom_track_25.INVTX1_4_.out
rlabel metal1 20838 17272 20838 17272 0 mux_bottom_track_25.INVTX1_5_.out
rlabel metal1 24564 17034 24564 17034 0 mux_bottom_track_25.INVTX1_6_.out
rlabel metal2 8510 16286 8510 16286 0 mux_bottom_track_25.INVTX1_7_.out
rlabel metal3 13087 15300 13087 15300 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal4 12604 13328 12604 13328 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 15226 15487 15226 15487 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 32430 2907 32430 2907 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 33074 3842 33074 3842 0 mux_bottom_track_25.out
rlabel metal2 25806 20706 25806 20706 0 mux_bottom_track_33.INVTX1_0_.out
rlabel metal1 22126 20332 22126 20332 0 mux_bottom_track_33.INVTX1_1_.out
rlabel metal1 9660 21930 9660 21930 0 mux_bottom_track_33.INVTX1_2_.out
rlabel metal1 6394 16218 6394 16218 0 mux_bottom_track_33.INVTX1_3_.out
rlabel metal1 20608 30634 20608 30634 0 mux_bottom_track_33.INVTX1_4_.out
rlabel metal2 13110 27370 13110 27370 0 mux_bottom_track_33.INVTX1_5_.out
rlabel metal1 10258 20536 10258 20536 0 mux_bottom_track_33.INVTX1_6_.out
rlabel metal1 10350 15402 10350 15402 0 mux_bottom_track_33.INVTX1_7_.out
rlabel via2 23782 21029 23782 21029 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 13478 23358 13478 23358 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 11270 20366 11270 20366 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 24978 35666 24978 35666 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 36846 35972 36846 35972 0 mux_bottom_track_33.out
rlabel metal1 23276 13362 23276 13362 0 mux_bottom_track_9.INVTX1_0_.out
rlabel metal1 25714 14484 25714 14484 0 mux_bottom_track_9.INVTX1_1_.out
rlabel metal1 27738 28390 27738 28390 0 mux_bottom_track_9.INVTX1_2_.out
rlabel metal1 4508 17102 4508 17102 0 mux_bottom_track_9.INVTX1_3_.out
rlabel metal1 15410 20366 15410 20366 0 mux_bottom_track_9.INVTX1_4_.out
rlabel via2 2438 3077 2438 3077 0 mux_bottom_track_9.INVTX1_5_.out
rlabel metal1 27508 23494 27508 23494 0 mux_bottom_track_9.INVTX1_6_.out
rlabel metal1 12190 18768 12190 18768 0 mux_bottom_track_9.INVTX1_7_.out
rlabel metal2 23230 3604 23230 3604 0 mux_bottom_track_9.INVTX1_8_.out
rlabel metal1 13662 17782 13662 17782 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 16698 20366 16698 20366 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 34868 21998 34868 21998 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 36294 21998 36294 21998 0 mux_bottom_track_9.out
rlabel metal3 4715 20740 4715 20740 0 mux_left_track_1.INVTX1_1_.out
rlabel metal1 16146 19482 16146 19482 0 mux_left_track_1.INVTX1_2_.out
rlabel metal1 29716 13362 29716 13362 0 mux_left_track_1.INVTX1_3_.out
rlabel metal1 21666 14450 21666 14450 0 mux_left_track_1.INVTX1_4_.out
rlabel metal1 19872 14926 19872 14926 0 mux_left_track_1.mux_2level_tapbuf_basis_input2_mem2_0_out
rlabel metal2 4830 18768 4830 18768 0 mux_left_track_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 31050 31858 31050 31858 0 mux_left_track_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 31142 32436 31142 32436 0 mux_left_track_1.out
rlabel metal1 11914 25806 11914 25806 0 mux_left_track_11.INVTX1_1_.out
rlabel metal1 6716 34510 6716 34510 0 mux_left_track_11.INVTX1_2_.out
rlabel metal2 12466 27268 12466 27268 0 mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 13064 26214 13064 26214 0 mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 13478 28900 13478 28900 0 mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 14444 35054 14444 35054 0 mux_left_track_11.out
rlabel metal2 22126 15708 22126 15708 0 mux_left_track_13.INVTX1_1_.out
rlabel metal1 26404 12954 26404 12954 0 mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 30406 8704 30406 8704 0 mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 33166 10098 33166 10098 0 mux_left_track_13.out
rlabel metal1 14306 18190 14306 18190 0 mux_left_track_15.INVTX1_1_.out
rlabel metal2 16146 16082 16146 16082 0 mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 28336 14790 28336 14790 0 mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 32476 14382 32476 14382 0 mux_left_track_15.out
rlabel metal1 25530 18190 25530 18190 0 mux_left_track_17.INVTX1_1_.out
rlabel metal1 29762 18700 29762 18700 0 mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 30222 17782 30222 17782 0 mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 35190 18564 35190 18564 0 mux_left_track_17.out
rlabel metal2 23322 20910 23322 20910 0 mux_left_track_19.INVTX1_1_.out
rlabel metal1 25346 20298 25346 20298 0 mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 29302 13158 29302 13158 0 mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 27646 8993 27646 8993 0 mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 27370 6290 27370 6290 0 mux_left_track_19.out
rlabel metal1 24610 24276 24610 24276 0 mux_left_track_21.INVTX1_1_.out
rlabel metal1 24932 24310 24932 24310 0 mux_left_track_21.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 24104 25670 24104 25670 0 mux_left_track_21.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 26404 19958 26404 19958 0 mux_left_track_21.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 31326 16252 31326 16252 0 mux_left_track_21.out
rlabel metal2 14766 17680 14766 17680 0 mux_left_track_23.INVTX1_1_.out
rlabel metal1 27186 13294 27186 13294 0 mux_left_track_23.INVTX1_2_.out
rlabel metal1 28106 18156 28106 18156 0 mux_left_track_23.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 27508 13498 27508 13498 0 mux_left_track_23.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 28842 12614 28842 12614 0 mux_left_track_23.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 30222 7548 30222 7548 0 mux_left_track_23.out
rlabel metal1 14950 24718 14950 24718 0 mux_left_track_25.INVTX1_1_.out
rlabel metal2 28106 30464 28106 30464 0 mux_left_track_25.INVTX1_2_.out
rlabel metal1 14720 24378 14720 24378 0 mux_left_track_25.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 15318 26112 15318 26112 0 mux_left_track_25.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 12650 26010 12650 26010 0 mux_left_track_25.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 9522 26282 9522 26282 0 mux_left_track_25.out
rlabel metal2 2254 6494 2254 6494 0 mux_left_track_27.INVTX1_1_.out
rlabel metal1 2576 7514 2576 7514 0 mux_left_track_27.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 3082 14688 3082 14688 0 mux_left_track_27.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 3910 14042 3910 14042 0 mux_left_track_27.out
rlabel metal2 24702 13804 24702 13804 0 mux_left_track_3.INVTX1_1_.out
rlabel metal2 33626 4318 33626 4318 0 mux_left_track_3.INVTX1_2_.out
rlabel metal1 23782 14450 23782 14450 0 mux_left_track_3.mux_2level_tapbuf_basis_input2_mem2_0_out
rlabel metal1 23506 13396 23506 13396 0 mux_left_track_3.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 32338 4658 32338 4658 0 mux_left_track_3.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 33718 4114 33718 4114 0 mux_left_track_3.out
rlabel metal2 33626 17374 33626 17374 0 mux_left_track_37.INVTX1_0_.out
rlabel metal2 28198 16354 28198 16354 0 mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 26036 25262 26036 25262 0 mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 23506 33490 23506 33490 0 mux_left_track_37.out
rlabel metal1 11730 29002 11730 29002 0 mux_left_track_5.INVTX1_1_.out
rlabel via1 27094 3587 27094 3587 0 mux_left_track_5.INVTX1_2_.out
rlabel metal1 22862 16014 22862 16014 0 mux_left_track_5.mux_2level_tapbuf_basis_input2_mem2_0_out
rlabel metal2 19550 16864 19550 16864 0 mux_left_track_5.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 24472 24378 24472 24378 0 mux_left_track_5.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 26404 24786 26404 24786 0 mux_left_track_5.out
rlabel metal1 12765 17102 12765 17102 0 mux_left_track_7.INVTX1_1_.out
rlabel metal1 17434 20366 17434 20366 0 mux_left_track_7.INVTX1_2_.out
rlabel metal1 18032 20842 18032 20842 0 mux_left_track_7.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 23506 23256 23506 23256 0 mux_left_track_7.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 29670 31348 29670 31348 0 mux_left_track_7.out
rlabel metal1 26450 18802 26450 18802 0 mux_left_track_9.INVTX1_1_.out
rlabel metal1 17066 33286 17066 33286 0 mux_left_track_9.INVTX1_2_.out
rlabel metal1 26726 20570 26726 20570 0 mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 20746 24276 20746 24276 0 mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 27554 23392 27554 23392 0 mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 30130 29818 30130 29818 0 mux_left_track_9.out
rlabel metal2 31786 7752 31786 7752 0 mux_top_track_0.INVTX1_0_.out
rlabel metal1 23552 31858 23552 31858 0 mux_top_track_0.INVTX1_1_.out
rlabel metal2 21942 14484 21942 14484 0 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 14260 15538 14260 15538 0 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 37398 11917 37398 11917 0 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 37766 10030 37766 10030 0 mux_top_track_0.out
rlabel metal1 22954 24684 22954 24684 0 mux_top_track_16.INVTX1_0_.out
rlabel metal1 8096 31790 8096 31790 0 mux_top_track_16.INVTX1_1_.out
rlabel metal2 9614 20553 9614 20553 0 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 14306 17323 14306 17323 0 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 7866 14399 7866 14399 0 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 4738 13770 4738 13770 0 mux_top_track_16.out
rlabel metal1 27554 2482 27554 2482 0 mux_top_track_24.INVTX1_0_.out
rlabel metal1 24334 3128 24334 3128 0 mux_top_track_24.INVTX1_1_.out
rlabel metal2 20286 17408 20286 17408 0 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 18630 19448 18630 19448 0 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 36202 22372 36202 22372 0 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 36708 30906 36708 30906 0 mux_top_track_24.out
rlabel metal1 27370 31858 27370 31858 0 mux_top_track_32.INVTX1_0_.out
rlabel metal1 8602 17102 8602 17102 0 mux_top_track_32.INVTX1_1_.out
rlabel metal1 27232 22542 27232 22542 0 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 25438 22984 25438 22984 0 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 20102 21352 20102 21352 0 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 13432 21454 13432 21454 0 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 8464 25942 8464 25942 0 mux_top_track_32.out
rlabel metal2 23046 5916 23046 5916 0 mux_top_track_8.INVTX1_0_.out
rlabel metal1 6992 16694 6992 16694 0 mux_top_track_8.INVTX1_1_.out
rlabel metal1 13432 16014 13432 16014 0 mux_top_track_8.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 20332 15946 20332 15946 0 mux_top_track_8.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 16790 16694 16790 16694 0 mux_top_track_8.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 14720 16150 14720 16150 0 mux_top_track_8.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 22034 31790 22034 31790 0 mux_top_track_8.out
rlabel metal1 1610 18836 1610 18836 0 net1
rlabel metal1 4416 36006 4416 36006 0 net10
rlabel metal2 38042 14076 38042 14076 0 net100
rlabel metal2 36938 19142 36938 19142 0 net101
rlabel metal1 27784 2414 27784 2414 0 net102
rlabel metal1 4324 23562 4324 23562 0 net103
rlabel metal2 25530 32368 25530 32368 0 net104
rlabel metal1 1978 32878 1978 32878 0 net105
rlabel metal1 30774 2414 30774 2414 0 net106
rlabel metal2 22862 24208 22862 24208 0 net107
rlabel metal1 36961 5678 36961 5678 0 net108
rlabel metal2 27186 37060 27186 37060 0 net109
rlabel metal1 10248 3706 10248 3706 0 net11
rlabel metal2 36662 36550 36662 36550 0 net110
rlabel metal1 37766 36754 37766 36754 0 net111
rlabel metal1 1610 3094 1610 3094 0 net112
rlabel metal1 3266 14042 3266 14042 0 net113
rlabel metal1 37996 3026 37996 3026 0 net114
rlabel metal2 1610 11135 1610 11135 0 net115
rlabel metal1 38042 21964 38042 21964 0 net116
rlabel metal2 38042 16252 38042 16252 0 net117
rlabel metal1 16928 37230 16928 37230 0 net118
rlabel via3 3197 2652 3197 2652 0 net119
rlabel metal1 24288 30702 24288 30702 0 net12
rlabel metal2 38042 4794 38042 4794 0 net120
rlabel metal1 36961 17170 36961 17170 0 net121
rlabel metal1 37950 10234 37950 10234 0 net122
rlabel metal2 1978 24548 1978 24548 0 net123
rlabel metal1 37950 21114 37950 21114 0 net124
rlabel metal1 37490 31994 37490 31994 0 net125
rlabel metal1 36662 2448 36662 2448 0 net126
rlabel metal1 37950 36142 37950 36142 0 net127
rlabel metal1 1610 12784 1610 12784 0 net128
rlabel metal1 2346 34578 2346 34578 0 net129
rlabel metal2 6578 36992 6578 36992 0 net13
rlabel via2 2254 3587 2254 3587 0 net130
rlabel metal1 2484 2414 2484 2414 0 net131
rlabel metal3 1771 5372 1771 5372 0 net132
rlabel metal2 1702 28492 1702 28492 0 net133
rlabel metal2 10442 37060 10442 37060 0 net134
rlabel metal1 22816 31994 22816 31994 0 net135
rlabel metal1 1656 19482 1656 19482 0 net136
rlabel metal2 13662 4573 13662 4573 0 net137
rlabel via3 1725 2652 1725 2652 0 net138
rlabel metal1 1610 8976 1610 8976 0 net139
rlabel metal1 31602 3366 31602 3366 0 net14
rlabel metal1 21620 29274 21620 29274 0 net140
rlabel metal1 37766 3910 37766 3910 0 net141
rlabel metal1 27048 7514 27048 7514 0 net142
rlabel metal2 7590 14620 7590 14620 0 net143
rlabel metal1 27554 14042 27554 14042 0 net144
rlabel metal2 5658 21216 5658 21216 0 net145
rlabel metal2 26266 11424 26266 11424 0 net146
rlabel metal1 26542 4522 26542 4522 0 net147
rlabel metal1 14398 16456 14398 16456 0 net148
rlabel metal2 19642 21216 19642 21216 0 net149
rlabel metal1 9476 36550 9476 36550 0 net15
rlabel metal1 24702 14926 24702 14926 0 net150
rlabel metal2 9798 22814 9798 22814 0 net151
rlabel metal2 22218 17374 22218 17374 0 net152
rlabel via1 31786 3349 31786 3349 0 net153
rlabel metal2 18906 17374 18906 17374 0 net154
rlabel metal2 20378 22848 20378 22848 0 net155
rlabel metal2 20102 23868 20102 23868 0 net156
rlabel metal1 12765 25262 12765 25262 0 net157
rlabel metal2 30682 12988 30682 12988 0 net158
rlabel metal2 23138 26044 23138 26044 0 net159
rlabel metal2 22218 4692 22218 4692 0 net16
rlabel metal1 29302 13906 29302 13906 0 net160
rlabel metal1 14720 25874 14720 25874 0 net161
rlabel metal2 29302 8976 29302 8976 0 net162
rlabel metal1 28888 14926 28888 14926 0 net163
rlabel metal2 28198 17340 28198 17340 0 net164
rlabel metal2 2438 15164 2438 15164 0 net165
rlabel metal2 29854 16864 29854 16864 0 net166
rlabel metal2 1610 16796 1610 16796 0 net17
rlabel metal2 2254 9112 2254 9112 0 net18
rlabel metal1 23414 30260 23414 30260 0 net19
rlabel metal1 1564 6630 1564 6630 0 net2
rlabel metal1 10948 3026 10948 3026 0 net20
rlabel metal1 37904 32198 37904 32198 0 net21
rlabel metal1 32522 23698 32522 23698 0 net22
rlabel metal2 2898 4012 2898 4012 0 net23
rlabel metal1 6578 8432 6578 8432 0 net24
rlabel metal2 38134 8636 38134 8636 0 net25
rlabel metal1 14766 30226 14766 30226 0 net26
rlabel metal2 38134 26047 38134 26047 0 net27
rlabel metal1 38042 29002 38042 29002 0 net28
rlabel metal1 31832 37094 31832 37094 0 net29
rlabel metal1 5750 37094 5750 37094 0 net3
rlabel via2 13386 2805 13386 2805 0 net30
rlabel metal1 37398 36006 37398 36006 0 net31
rlabel metal1 38226 20910 38226 20910 0 net32
rlabel metal2 24610 33932 24610 33932 0 net33
rlabel metal2 22494 36589 22494 36589 0 net34
rlabel metal1 37904 30226 37904 30226 0 net35
rlabel metal1 8878 37230 8878 37230 0 net36
rlabel metal1 13570 33490 13570 33490 0 net37
rlabel metal2 22954 31484 22954 31484 0 net38
rlabel metal1 2530 5678 2530 5678 0 net39
rlabel metal2 1978 9316 1978 9316 0 net4
rlabel metal1 2990 36550 2990 36550 0 net40
rlabel metal2 38226 14892 38226 14892 0 net41
rlabel metal1 4278 37196 4278 37196 0 net42
rlabel metal2 34730 3876 34730 3876 0 net43
rlabel metal1 1932 19346 1932 19346 0 net44
rlabel metal1 36823 7922 36823 7922 0 net45
rlabel metal2 2162 24480 2162 24480 0 net46
rlabel metal2 5106 3434 5106 3434 0 net47
rlabel metal2 22126 28407 22126 28407 0 net48
rlabel metal2 16330 3485 16330 3485 0 net49
rlabel metal1 35098 2890 35098 2890 0 net5
rlabel metal2 5658 18887 5658 18887 0 net50
rlabel metal1 2438 37230 2438 37230 0 net51
rlabel metal1 34178 12410 34178 12410 0 net52
rlabel metal2 1886 20706 1886 20706 0 net53
rlabel metal2 1886 36249 1886 36249 0 net54
rlabel metal2 37766 36958 37766 36958 0 net55
rlabel metal1 30728 22610 30728 22610 0 net56
rlabel metal1 1886 18326 1886 18326 0 net57
rlabel metal1 16560 1700 16560 1700 0 net58
rlabel metal2 37766 12002 37766 12002 0 net59
rlabel metal2 32982 4420 32982 4420 0 net6
rlabel metal1 17388 37366 17388 37366 0 net60
rlabel metal1 32614 3672 32614 3672 0 net61
rlabel metal2 4002 8058 4002 8058 0 net62
rlabel metal2 12926 3366 12926 3366 0 net63
rlabel metal1 38042 4794 38042 4794 0 net64
rlabel metal2 38226 28492 38226 28492 0 net65
rlabel metal2 34730 19482 34730 19482 0 net66
rlabel metal1 32798 17170 32798 17170 0 net67
rlabel metal2 1886 24004 1886 24004 0 net68
rlabel via2 12006 2907 12006 2907 0 net69
rlabel metal1 8740 21998 8740 21998 0 net7
rlabel metal1 33718 36550 33718 36550 0 net70
rlabel metal2 34086 9622 34086 9622 0 net71
rlabel metal1 3588 35462 3588 35462 0 net72
rlabel metal1 1610 11016 1610 11016 0 net73
rlabel metal1 18446 11016 18446 11016 0 net74
rlabel metal1 22218 2550 22218 2550 0 net75
rlabel metal1 32844 25262 32844 25262 0 net76
rlabel metal1 28474 2618 28474 2618 0 net77
rlabel metal1 29256 31858 29256 31858 0 net78
rlabel metal2 25714 32028 25714 32028 0 net79
rlabel metal1 1748 8602 1748 8602 0 net8
rlabel metal1 4968 36550 4968 36550 0 net80
rlabel metal1 7590 37094 7590 37094 0 net81
rlabel metal2 32338 3740 32338 3740 0 net82
rlabel metal1 1794 10778 1794 10778 0 net83
rlabel metal2 21574 5593 21574 5593 0 net84
rlabel metal1 36110 37230 36110 37230 0 net85
rlabel metal2 34454 13804 34454 13804 0 net86
rlabel metal1 33534 2414 33534 2414 0 net87
rlabel metal1 1610 30668 1610 30668 0 net88
rlabel metal1 1610 16116 1610 16116 0 net89
rlabel metal1 17664 37094 17664 37094 0 net9
rlabel metal2 20194 26962 20194 26962 0 net90
rlabel metal1 31602 22746 31602 22746 0 net91
rlabel metal1 35742 2414 35742 2414 0 net92
rlabel metal1 20792 33626 20792 33626 0 net93
rlabel metal1 34868 2414 34868 2414 0 net94
rlabel metal1 29532 36890 29532 36890 0 net95
rlabel metal1 34086 37230 34086 37230 0 net96
rlabel metal2 35926 34102 35926 34102 0 net97
rlabel metal1 15410 35258 15410 35258 0 net98
rlabel metal2 36938 10914 36938 10914 0 net99
rlabel metal3 1234 10948 1234 10948 0 pReset
rlabel metal1 7406 2822 7406 2822 0 prog_clk
rlabel metal2 13570 823 13570 823 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
rlabel metal2 21298 1588 21298 1588 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
rlabel metal3 38786 25908 38786 25908 0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 22586 1520 22586 1520 0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 30406 37230 30406 37230 0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 29486 37230 29486 37230 0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 3312 36754 3312 36754 0 top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal1 7268 37230 7268 37230 0 top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_
rlabel metal2 27094 823 27094 823 0 top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal3 1234 10268 1234 10268 0 top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
