magic
tech sky130A
magscale 1 2
timestamp 1674229378
<< viali >>
rect 22753 37417 22787 37451
rect 23949 37417 23983 37451
rect 36737 37417 36771 37451
rect 20177 37349 20211 37383
rect 3157 37281 3191 37315
rect 3433 37281 3467 37315
rect 4169 37281 4203 37315
rect 4445 37281 4479 37315
rect 8309 37281 8343 37315
rect 10609 37281 10643 37315
rect 11713 37281 11747 37315
rect 13185 37281 13219 37315
rect 15117 37281 15151 37315
rect 16865 37281 16899 37315
rect 18705 37281 18739 37315
rect 29929 37281 29963 37315
rect 30389 37281 30423 37315
rect 8585 37213 8619 37247
rect 10885 37213 10919 37247
rect 13461 37213 13495 37247
rect 14841 37213 14875 37247
rect 15853 37213 15887 37247
rect 17049 37213 17083 37247
rect 17601 37213 17635 37247
rect 19441 37213 19475 37247
rect 20913 37213 20947 37247
rect 21373 37213 21407 37247
rect 22017 37213 22051 37247
rect 24777 37213 24811 37247
rect 25329 37213 25363 37247
rect 27169 37213 27203 37247
rect 28917 37213 28951 37247
rect 30665 37213 30699 37247
rect 32321 37213 32355 37247
rect 33609 37213 33643 37247
rect 35541 37213 35575 37247
rect 36921 37213 36955 37247
rect 37473 37213 37507 37247
rect 1685 37077 1719 37111
rect 5917 37077 5951 37111
rect 6837 37077 6871 37111
rect 9137 37077 9171 37111
rect 15669 37077 15703 37111
rect 18153 37077 18187 37111
rect 19625 37077 19659 37111
rect 20729 37077 20763 37111
rect 22201 37077 22235 37111
rect 23305 37077 23339 37111
rect 24685 37077 24719 37111
rect 25513 37077 25547 37111
rect 26525 37077 26559 37111
rect 27353 37077 27387 37111
rect 29101 37077 29135 37111
rect 31769 37077 31803 37111
rect 32505 37077 32539 37111
rect 33793 37077 33827 37111
rect 35725 37077 35759 37111
rect 37657 37077 37691 37111
rect 16037 36873 16071 36907
rect 38209 36873 38243 36907
rect 2329 36805 2363 36839
rect 5733 36805 5767 36839
rect 11713 36805 11747 36839
rect 13461 36805 13495 36839
rect 17693 36805 17727 36839
rect 2053 36737 2087 36771
rect 6929 36737 6963 36771
rect 13737 36737 13771 36771
rect 14473 36737 14507 36771
rect 14933 36737 14967 36771
rect 15853 36737 15887 36771
rect 17049 36737 17083 36771
rect 17785 36737 17819 36771
rect 18889 36737 18923 36771
rect 19533 36737 19567 36771
rect 23397 36737 23431 36771
rect 25421 36737 25455 36771
rect 26065 36737 26099 36771
rect 32505 36737 32539 36771
rect 33149 36737 33183 36771
rect 34345 36737 34379 36771
rect 34989 36737 35023 36771
rect 38025 36737 38059 36771
rect 6009 36669 6043 36703
rect 7205 36669 7239 36703
rect 8677 36669 8711 36703
rect 9137 36669 9171 36703
rect 10885 36669 10919 36703
rect 11161 36669 11195 36703
rect 32597 36669 32631 36703
rect 14289 36601 14323 36635
rect 21097 36601 21131 36635
rect 22017 36601 22051 36635
rect 22569 36601 22603 36635
rect 24041 36601 24075 36635
rect 24593 36601 24627 36635
rect 25605 36601 25639 36635
rect 3801 36533 3835 36567
rect 4261 36533 4295 36567
rect 15025 36533 15059 36567
rect 16865 36533 16899 36567
rect 18797 36533 18831 36567
rect 19441 36533 19475 36567
rect 19993 36533 20027 36567
rect 20545 36533 20579 36567
rect 23581 36533 23615 36567
rect 34437 36533 34471 36567
rect 4432 36329 4466 36363
rect 13185 36329 13219 36363
rect 20545 36329 20579 36363
rect 22201 36329 22235 36363
rect 22753 36329 22787 36363
rect 23305 36329 23339 36363
rect 23857 36329 23891 36363
rect 25145 36329 25179 36363
rect 38209 36329 38243 36363
rect 1685 36193 1719 36227
rect 4169 36193 4203 36227
rect 6377 36193 6411 36227
rect 8125 36193 8159 36227
rect 12357 36193 12391 36227
rect 12633 36193 12667 36227
rect 19441 36193 19475 36227
rect 19993 36193 20027 36227
rect 21097 36193 21131 36227
rect 8401 36125 8435 36159
rect 9873 36125 9907 36159
rect 10149 36125 10183 36159
rect 13369 36125 13403 36159
rect 14657 36125 14691 36159
rect 15301 36125 15335 36159
rect 15761 36125 15795 36159
rect 17969 36125 18003 36159
rect 38025 36125 38059 36159
rect 1961 36057 1995 36091
rect 10609 36057 10643 36091
rect 3433 35989 3467 36023
rect 5917 35989 5951 36023
rect 14565 35989 14599 36023
rect 15209 35989 15243 36023
rect 15853 35989 15887 36023
rect 16405 35989 16439 36023
rect 17509 35989 17543 36023
rect 18521 35989 18555 36023
rect 21649 35989 21683 36023
rect 24593 35989 24627 36023
rect 25697 35989 25731 36023
rect 17693 35785 17727 35819
rect 20085 35785 20119 35819
rect 20637 35785 20671 35819
rect 21189 35785 21223 35819
rect 22017 35785 22051 35819
rect 23121 35785 23155 35819
rect 23673 35785 23707 35819
rect 24777 35785 24811 35819
rect 27537 35785 27571 35819
rect 1685 35717 1719 35751
rect 5089 35717 5123 35751
rect 8677 35717 8711 35751
rect 13185 35717 13219 35751
rect 14013 35717 14047 35751
rect 18981 35717 19015 35751
rect 5365 35649 5399 35683
rect 6009 35649 6043 35683
rect 8953 35649 8987 35683
rect 13461 35649 13495 35683
rect 14473 35649 14507 35683
rect 15485 35649 15519 35683
rect 16313 35649 16347 35683
rect 16865 35649 16899 35683
rect 17785 35649 17819 35683
rect 27445 35649 27479 35683
rect 38025 35649 38059 35683
rect 2881 35581 2915 35615
rect 3157 35581 3191 35615
rect 7205 35581 7239 35615
rect 10885 35581 10919 35615
rect 11161 35581 11195 35615
rect 25329 35581 25363 35615
rect 1869 35513 1903 35547
rect 11713 35513 11747 35547
rect 24225 35513 24259 35547
rect 3617 35445 3651 35479
rect 5917 35445 5951 35479
rect 6653 35445 6687 35479
rect 9413 35445 9447 35479
rect 14565 35445 14599 35479
rect 15669 35445 15703 35479
rect 16221 35445 16255 35479
rect 16957 35445 16991 35479
rect 18521 35445 18555 35479
rect 19533 35445 19567 35479
rect 22569 35445 22603 35479
rect 37473 35445 37507 35479
rect 38209 35445 38243 35479
rect 3433 35241 3467 35275
rect 18061 35241 18095 35275
rect 18705 35241 18739 35275
rect 21097 35241 21131 35275
rect 22201 35241 22235 35275
rect 9367 35173 9401 35207
rect 21649 35173 21683 35207
rect 1685 35105 1719 35139
rect 5457 35105 5491 35139
rect 10885 35105 10919 35139
rect 19993 35105 20027 35139
rect 20545 35105 20579 35139
rect 5733 35037 5767 35071
rect 6285 35037 6319 35071
rect 9137 35037 9171 35071
rect 13553 35037 13587 35071
rect 14289 35037 14323 35071
rect 15393 35037 15427 35071
rect 16129 35037 16163 35071
rect 16221 35037 16255 35071
rect 16865 35037 16899 35071
rect 16957 35037 16991 35071
rect 18797 35037 18831 35071
rect 1961 34969 1995 35003
rect 6561 34969 6595 35003
rect 8309 34969 8343 35003
rect 11161 34969 11195 35003
rect 12909 34969 12943 35003
rect 17785 34969 17819 35003
rect 22753 34969 22787 35003
rect 24593 34969 24627 35003
rect 3985 34901 4019 34935
rect 13645 34901 13679 34935
rect 14381 34901 14415 34935
rect 15485 34901 15519 34935
rect 19533 34901 19567 34935
rect 23305 34901 23339 34935
rect 23857 34901 23891 34935
rect 19165 34697 19199 34731
rect 20361 34697 20395 34731
rect 20821 34697 20855 34731
rect 22569 34697 22603 34731
rect 23673 34697 23707 34731
rect 24225 34697 24259 34731
rect 14105 34629 14139 34663
rect 16221 34629 16255 34663
rect 23121 34629 23155 34663
rect 1777 34561 1811 34595
rect 3985 34561 4019 34595
rect 6745 34561 6779 34595
rect 10977 34561 11011 34595
rect 11713 34561 11747 34595
rect 15485 34561 15519 34595
rect 16129 34561 16163 34595
rect 17325 34561 17359 34595
rect 17969 34561 18003 34595
rect 18429 34561 18463 34595
rect 19257 34561 19291 34595
rect 19717 34561 19751 34595
rect 3525 34493 3559 34527
rect 8493 34493 8527 34527
rect 8953 34493 8987 34527
rect 11989 34493 12023 34527
rect 13461 34493 13495 34527
rect 14013 34493 14047 34527
rect 14473 34493 14507 34527
rect 15577 34493 15611 34527
rect 17049 34493 17083 34527
rect 17877 34493 17911 34527
rect 18521 34493 18555 34527
rect 21373 34493 21407 34527
rect 5733 34425 5767 34459
rect 22017 34425 22051 34459
rect 2040 34357 2074 34391
rect 4248 34357 4282 34391
rect 7002 34357 7036 34391
rect 9216 34357 9250 34391
rect 9400 34153 9434 34187
rect 20177 34153 20211 34187
rect 21281 34153 21315 34187
rect 22937 34153 22971 34187
rect 23489 34153 23523 34187
rect 24593 34153 24627 34187
rect 3433 34017 3467 34051
rect 3985 34017 4019 34051
rect 9137 34017 9171 34051
rect 11161 34017 11195 34051
rect 11621 34017 11655 34051
rect 16497 34017 16531 34051
rect 6285 33949 6319 33983
rect 16773 33949 16807 33983
rect 17233 33949 17267 33983
rect 17509 33949 17543 33983
rect 18153 33949 18187 33983
rect 20269 33949 20303 33983
rect 3157 33881 3191 33915
rect 4261 33881 4295 33915
rect 6561 33881 6595 33915
rect 8309 33881 8343 33915
rect 11897 33881 11931 33915
rect 14473 33881 14507 33915
rect 15393 33881 15427 33915
rect 15485 33881 15519 33915
rect 18429 33881 18463 33915
rect 20729 33881 20763 33915
rect 22385 33881 22419 33915
rect 1685 33813 1719 33847
rect 5733 33813 5767 33847
rect 13369 33813 13403 33847
rect 19441 33813 19475 33847
rect 21833 33813 21867 33847
rect 20729 33609 20763 33643
rect 22017 33609 22051 33643
rect 22661 33609 22695 33643
rect 23121 33609 23155 33643
rect 24225 33609 24259 33643
rect 24777 33609 24811 33643
rect 5733 33541 5767 33575
rect 9413 33541 9447 33575
rect 15761 33541 15795 33575
rect 18797 33541 18831 33575
rect 19533 33541 19567 33575
rect 19625 33541 19659 33575
rect 3525 33473 3559 33507
rect 9137 33473 9171 33507
rect 11713 33473 11747 33507
rect 13737 33473 13771 33507
rect 14657 33473 14691 33507
rect 16313 33473 16347 33507
rect 17325 33473 17359 33507
rect 37565 33473 37599 33507
rect 38209 33473 38243 33507
rect 1777 33405 1811 33439
rect 3249 33405 3283 33439
rect 3985 33405 4019 33439
rect 6009 33405 6043 33439
rect 6837 33405 6871 33439
rect 7113 33405 7147 33439
rect 11161 33405 11195 33439
rect 15669 33405 15703 33439
rect 17141 33405 17175 33439
rect 18613 33405 18647 33439
rect 18889 33405 18923 33439
rect 19809 33405 19843 33439
rect 23673 33337 23707 33371
rect 38025 33337 38059 33371
rect 8585 33269 8619 33303
rect 11976 33269 12010 33303
rect 14749 33269 14783 33303
rect 21189 33269 21223 33303
rect 1685 33065 1719 33099
rect 9689 33065 9723 33099
rect 18061 33065 18095 33099
rect 18705 33065 18739 33099
rect 19533 33065 19567 33099
rect 20177 33065 20211 33099
rect 22017 33065 22051 33099
rect 22569 33065 22603 33099
rect 23581 33065 23615 33099
rect 24593 33065 24627 33099
rect 8401 32997 8435 33031
rect 15209 32997 15243 33031
rect 15945 32997 15979 33031
rect 3433 32929 3467 32963
rect 10885 32929 10919 32963
rect 16497 32929 16531 32963
rect 4077 32861 4111 32895
rect 4813 32861 4847 32895
rect 5825 32861 5859 32895
rect 8309 32861 8343 32895
rect 9597 32861 9631 32895
rect 10241 32861 10275 32895
rect 13553 32861 13587 32895
rect 14473 32861 14507 32895
rect 15301 32861 15335 32895
rect 17049 32861 17083 32895
rect 18153 32861 18187 32895
rect 18797 32861 18831 32895
rect 19625 32861 19659 32895
rect 20269 32861 20303 32895
rect 20913 32861 20947 32895
rect 21373 32861 21407 32895
rect 3157 32793 3191 32827
rect 4261 32793 4295 32827
rect 6101 32793 6135 32827
rect 7849 32793 7883 32827
rect 11161 32793 11195 32827
rect 12909 32793 12943 32827
rect 16405 32793 16439 32827
rect 17325 32793 17359 32827
rect 20821 32793 20855 32827
rect 4905 32725 4939 32759
rect 10333 32725 10367 32759
rect 13645 32725 13679 32759
rect 14565 32725 14599 32759
rect 23121 32725 23155 32759
rect 21097 32521 21131 32555
rect 22661 32521 22695 32555
rect 23121 32521 23155 32555
rect 23673 32521 23707 32555
rect 6009 32453 6043 32487
rect 8309 32453 8343 32487
rect 13185 32453 13219 32487
rect 14105 32453 14139 32487
rect 15485 32453 15519 32487
rect 17877 32453 17911 32487
rect 18429 32453 18463 32487
rect 3525 32385 3559 32419
rect 3985 32385 4019 32419
rect 8585 32385 8619 32419
rect 9321 32385 9355 32419
rect 14657 32385 14691 32419
rect 17049 32385 17083 32419
rect 19901 32385 19935 32419
rect 20361 32385 20395 32419
rect 21005 32385 21039 32419
rect 37565 32385 37599 32419
rect 38209 32385 38243 32419
rect 3249 32317 3283 32351
rect 4261 32317 4295 32351
rect 6561 32317 6595 32351
rect 9597 32317 9631 32351
rect 13461 32317 13495 32351
rect 14013 32317 14047 32351
rect 15393 32317 15427 32351
rect 17785 32317 17819 32351
rect 19257 32317 19291 32351
rect 11069 32249 11103 32283
rect 15945 32249 15979 32283
rect 22109 32249 22143 32283
rect 38025 32249 38059 32283
rect 1777 32181 1811 32215
rect 11713 32181 11747 32215
rect 17141 32181 17175 32215
rect 19809 32181 19843 32215
rect 20453 32181 20487 32215
rect 24225 32181 24259 32215
rect 16865 31977 16899 32011
rect 22477 31977 22511 32011
rect 9505 31909 9539 31943
rect 13001 31909 13035 31943
rect 15853 31909 15887 31943
rect 20729 31909 20763 31943
rect 23489 31909 23523 31943
rect 2605 31841 2639 31875
rect 3985 31841 4019 31875
rect 5457 31841 5491 31875
rect 11253 31841 11287 31875
rect 13645 31841 13679 31875
rect 17509 31841 17543 31875
rect 19441 31841 19475 31875
rect 20085 31841 20119 31875
rect 22937 31841 22971 31875
rect 2881 31773 2915 31807
rect 3433 31773 3467 31807
rect 5733 31773 5767 31807
rect 8493 31773 8527 31807
rect 12265 31773 12299 31807
rect 13093 31773 13127 31807
rect 13553 31783 13587 31817
rect 14749 31773 14783 31807
rect 16957 31773 16991 31807
rect 20821 31773 20855 31807
rect 21281 31773 21315 31807
rect 21833 31773 21867 31807
rect 6469 31705 6503 31739
rect 8217 31705 8251 31739
rect 10977 31705 11011 31739
rect 14657 31705 14691 31739
rect 15302 31705 15336 31739
rect 15393 31705 15427 31739
rect 17601 31705 17635 31739
rect 18521 31705 18555 31739
rect 19993 31705 20027 31739
rect 11805 31637 11839 31671
rect 12357 31637 12391 31671
rect 1685 31433 1719 31467
rect 3433 31433 3467 31467
rect 20361 31433 20395 31467
rect 21005 31433 21039 31467
rect 22109 31433 22143 31467
rect 23121 31433 23155 31467
rect 8401 31365 8435 31399
rect 13461 31365 13495 31399
rect 14565 31365 14599 31399
rect 17049 31365 17083 31399
rect 19625 31365 19659 31399
rect 19717 31365 19751 31399
rect 1869 31297 1903 31331
rect 2421 31297 2455 31331
rect 3341 31297 3375 31331
rect 3985 31297 4019 31331
rect 8677 31297 8711 31331
rect 11161 31297 11195 31331
rect 11713 31297 11747 31331
rect 13737 31297 13771 31331
rect 15117 31297 15151 31331
rect 15761 31297 15795 31331
rect 18613 31297 18647 31331
rect 20453 31297 20487 31331
rect 20913 31297 20947 31331
rect 4261 31229 4295 31263
rect 6653 31229 6687 31263
rect 9137 31229 9171 31263
rect 10885 31229 10919 31263
rect 14473 31229 14507 31263
rect 16957 31229 16991 31263
rect 17877 31229 17911 31263
rect 2605 31161 2639 31195
rect 19165 31161 19199 31195
rect 22569 31161 22603 31195
rect 5733 31093 5767 31127
rect 15853 31093 15887 31127
rect 18521 31093 18555 31127
rect 3341 30889 3375 30923
rect 13645 30889 13679 30923
rect 23029 30889 23063 30923
rect 14749 30821 14783 30855
rect 15945 30821 15979 30855
rect 17785 30821 17819 30855
rect 3985 30753 4019 30787
rect 5457 30753 5491 30787
rect 6561 30753 6595 30787
rect 8309 30753 8343 30787
rect 11989 30753 12023 30787
rect 21281 30753 21315 30787
rect 21925 30753 21959 30787
rect 1869 30685 1903 30719
rect 2329 30685 2363 30719
rect 3249 30685 3283 30719
rect 5733 30685 5767 30719
rect 8585 30685 8619 30719
rect 9597 30685 9631 30719
rect 10241 30685 10275 30719
rect 12265 30685 12299 30719
rect 13093 30685 13127 30719
rect 13737 30685 13771 30719
rect 14657 30685 14691 30719
rect 16681 30685 16715 30719
rect 18521 30685 18555 30719
rect 20821 30685 20855 30719
rect 13001 30617 13035 30651
rect 15393 30617 15427 30651
rect 15485 30617 15519 30651
rect 17233 30617 17267 30651
rect 17325 30617 17359 30651
rect 19533 30617 19567 30651
rect 19625 30617 19659 30651
rect 20177 30617 20211 30651
rect 1685 30549 1719 30583
rect 2421 30549 2455 30583
rect 9689 30549 9723 30583
rect 16589 30549 16623 30583
rect 18429 30549 18463 30583
rect 20729 30549 20763 30583
rect 22385 30549 22419 30583
rect 16221 30345 16255 30379
rect 10425 30277 10459 30311
rect 11989 30277 12023 30311
rect 15485 30277 15519 30311
rect 17049 30277 17083 30311
rect 19533 30277 19567 30311
rect 20361 30277 20395 30311
rect 21465 30277 21499 30311
rect 3801 30209 3835 30243
rect 6009 30209 6043 30243
rect 9873 30209 9907 30243
rect 10333 30209 10367 30243
rect 10977 30209 11011 30243
rect 14473 30209 14507 30243
rect 16313 30209 16347 30243
rect 20913 30209 20947 30243
rect 3525 30141 3559 30175
rect 5733 30141 5767 30175
rect 7021 30141 7055 30175
rect 8769 30141 8803 30175
rect 9045 30141 9079 30175
rect 11713 30141 11747 30175
rect 15577 30141 15611 30175
rect 16957 30141 16991 30175
rect 17877 30141 17911 30175
rect 18981 30141 19015 30175
rect 19625 30141 19659 30175
rect 20269 30141 20303 30175
rect 22017 30141 22051 30175
rect 38025 30141 38059 30175
rect 38301 30141 38335 30175
rect 9781 30073 9815 30107
rect 13461 30073 13495 30107
rect 15025 30073 15059 30107
rect 2053 30005 2087 30039
rect 4261 30005 4295 30039
rect 11069 30005 11103 30039
rect 14381 30005 14415 30039
rect 18429 30005 18463 30039
rect 22661 30005 22695 30039
rect 6745 29801 6779 29835
rect 21097 29801 21131 29835
rect 38301 29801 38335 29835
rect 7389 29733 7423 29767
rect 8033 29733 8067 29767
rect 1961 29665 1995 29699
rect 3433 29665 3467 29699
rect 3985 29665 4019 29699
rect 11989 29665 12023 29699
rect 13277 29665 13311 29699
rect 14657 29665 14691 29699
rect 14933 29665 14967 29699
rect 18153 29665 18187 29699
rect 18797 29665 18831 29699
rect 20177 29665 20211 29699
rect 1685 29597 1719 29631
rect 6653 29597 6687 29631
rect 7289 29591 7323 29625
rect 7941 29597 7975 29631
rect 9321 29597 9355 29631
rect 21189 29597 21223 29631
rect 21833 29597 21867 29631
rect 4261 29529 4295 29563
rect 9965 29529 9999 29563
rect 11713 29529 11747 29563
rect 12633 29529 12667 29563
rect 13185 29529 13219 29563
rect 14841 29529 14875 29563
rect 15669 29529 15703 29563
rect 15761 29529 15795 29563
rect 16313 29529 16347 29563
rect 17049 29529 17083 29563
rect 17141 29529 17175 29563
rect 17693 29529 17727 29563
rect 18705 29529 18739 29563
rect 20361 29529 20395 29563
rect 20453 29529 20487 29563
rect 5733 29461 5767 29495
rect 9413 29461 9447 29495
rect 21741 29461 21775 29495
rect 22385 29461 22419 29495
rect 1685 29257 1719 29291
rect 2237 29257 2271 29291
rect 4997 29257 5031 29291
rect 5917 29257 5951 29291
rect 7941 29257 7975 29291
rect 8585 29257 8619 29291
rect 21189 29257 21223 29291
rect 23397 29257 23431 29291
rect 6653 29189 6687 29223
rect 10057 29189 10091 29223
rect 12633 29189 12667 29223
rect 13737 29189 13771 29223
rect 13829 29189 13863 29223
rect 14473 29189 14507 29223
rect 14565 29189 14599 29223
rect 15761 29189 15795 29223
rect 16313 29189 16347 29223
rect 17693 29189 17727 29223
rect 19257 29189 19291 29223
rect 19349 29189 19383 29223
rect 19901 29189 19935 29223
rect 20453 29189 20487 29223
rect 20545 29189 20579 29223
rect 2145 29121 2179 29155
rect 3249 29121 3283 29155
rect 5825 29121 5859 29155
rect 6561 29121 6595 29155
rect 7205 29121 7239 29155
rect 8041 29121 8075 29155
rect 10333 29121 10367 29155
rect 10977 29121 11011 29155
rect 11897 29121 11931 29155
rect 12541 29121 12575 29155
rect 17049 29121 17083 29155
rect 21097 29121 21131 29155
rect 22201 29121 22235 29155
rect 23213 29121 23247 29155
rect 30113 29121 30147 29155
rect 13553 29053 13587 29087
rect 15669 29053 15703 29087
rect 17601 29053 17635 29087
rect 22109 29053 22143 29087
rect 38025 29053 38059 29087
rect 38301 29053 38335 29087
rect 7297 28985 7331 29019
rect 11069 28985 11103 29019
rect 11989 28985 12023 29019
rect 15025 28985 15059 29019
rect 16957 28985 16991 29019
rect 18153 28985 18187 29019
rect 18797 28985 18831 29019
rect 22753 28985 22787 29019
rect 23857 28985 23891 29019
rect 30205 28985 30239 29019
rect 3512 28917 3546 28951
rect 2237 28713 2271 28747
rect 4721 28713 4755 28747
rect 14381 28713 14415 28747
rect 18521 28713 18555 28747
rect 19533 28713 19567 28747
rect 23305 28713 23339 28747
rect 4077 28645 4111 28679
rect 5365 28645 5399 28679
rect 6009 28645 6043 28679
rect 7849 28645 7883 28679
rect 17877 28645 17911 28679
rect 22201 28645 22235 28679
rect 38301 28645 38335 28679
rect 2881 28577 2915 28611
rect 12081 28577 12115 28611
rect 14933 28577 14967 28611
rect 15577 28577 15611 28611
rect 16681 28577 16715 28611
rect 20453 28577 20487 28611
rect 21741 28577 21775 28611
rect 2145 28509 2179 28543
rect 2789 28509 2823 28543
rect 3985 28509 4019 28543
rect 4629 28509 4663 28543
rect 5273 28509 5307 28543
rect 5917 28509 5951 28543
rect 6929 28509 6963 28543
rect 7757 28509 7791 28543
rect 8585 28509 8619 28543
rect 9621 28509 9655 28543
rect 12909 28509 12943 28543
rect 13553 28509 13587 28543
rect 18429 28509 18463 28543
rect 19441 28509 19475 28543
rect 20545 28509 20579 28543
rect 21189 28509 21223 28543
rect 7021 28441 7055 28475
rect 11805 28441 11839 28475
rect 15025 28441 15059 28475
rect 16037 28441 16071 28475
rect 16589 28441 16623 28475
rect 17325 28441 17359 28475
rect 17417 28441 17451 28475
rect 21097 28441 21131 28475
rect 22753 28441 22787 28475
rect 1685 28373 1719 28407
rect 8493 28373 8527 28407
rect 9689 28373 9723 28407
rect 10333 28373 10367 28407
rect 13001 28373 13035 28407
rect 13645 28373 13679 28407
rect 4997 28169 5031 28203
rect 7573 28169 7607 28203
rect 22017 28169 22051 28203
rect 23765 28169 23799 28203
rect 2421 28101 2455 28135
rect 6929 28101 6963 28135
rect 11897 28101 11931 28135
rect 13461 28101 13495 28135
rect 13553 28101 13587 28135
rect 15025 28101 15059 28135
rect 17417 28101 17451 28135
rect 17509 28101 17543 28135
rect 18429 28101 18463 28135
rect 18981 28101 19015 28135
rect 1685 28033 1719 28067
rect 2329 28033 2363 28067
rect 2973 28033 3007 28067
rect 3617 28033 3651 28067
rect 4261 28033 4295 28067
rect 5089 28033 5123 28067
rect 5825 28033 5859 28067
rect 6837 28033 6871 28067
rect 7481 28033 7515 28067
rect 10793 28033 10827 28067
rect 12449 28033 12483 28067
rect 16129 28033 16163 28067
rect 19625 28033 19659 28067
rect 20269 28033 20303 28067
rect 20821 28033 20855 28067
rect 20913 28033 20947 28067
rect 22753 28033 22787 28067
rect 3709 27965 3743 27999
rect 8585 27965 8619 27999
rect 10517 27965 10551 27999
rect 11805 27965 11839 27999
rect 15117 27965 15151 27999
rect 16221 27965 16255 27999
rect 18337 27965 18371 27999
rect 21373 27965 21407 27999
rect 1869 27897 1903 27931
rect 3065 27897 3099 27931
rect 13001 27897 13035 27931
rect 14565 27897 14599 27931
rect 16957 27897 16991 27931
rect 20177 27897 20211 27931
rect 23305 27897 23339 27931
rect 4353 27829 4387 27863
rect 5917 27829 5951 27863
rect 9045 27829 9079 27863
rect 19533 27829 19567 27863
rect 2145 27557 2179 27591
rect 4077 27557 4111 27591
rect 4721 27557 4755 27591
rect 6837 27557 6871 27591
rect 9413 27557 9447 27591
rect 13645 27557 13679 27591
rect 16405 27557 16439 27591
rect 22845 27557 22879 27591
rect 2789 27489 2823 27523
rect 8033 27489 8067 27523
rect 10333 27489 10367 27523
rect 11437 27489 11471 27523
rect 14381 27489 14415 27523
rect 17601 27489 17635 27523
rect 20545 27489 20579 27523
rect 20821 27489 20855 27523
rect 2053 27421 2087 27455
rect 2881 27421 2915 27455
rect 3985 27421 4019 27455
rect 4629 27421 4663 27455
rect 9321 27421 9355 27455
rect 12909 27421 12943 27455
rect 13553 27421 13587 27455
rect 16313 27421 16347 27455
rect 19441 27421 19475 27455
rect 23949 27421 23983 27455
rect 3433 27353 3467 27387
rect 8585 27353 8619 27387
rect 10517 27353 10551 27387
rect 10609 27353 10643 27387
rect 11713 27353 11747 27387
rect 11805 27353 11839 27387
rect 14473 27353 14507 27387
rect 15393 27353 15427 27387
rect 16957 27353 16991 27387
rect 17509 27353 17543 27387
rect 18153 27353 18187 27387
rect 18705 27353 18739 27387
rect 18797 27353 18831 27387
rect 20637 27353 20671 27387
rect 22385 27353 22419 27387
rect 5733 27285 5767 27319
rect 6377 27285 6411 27319
rect 7481 27285 7515 27319
rect 12449 27285 12483 27319
rect 13001 27285 13035 27319
rect 19533 27285 19567 27319
rect 21833 27285 21867 27319
rect 23397 27285 23431 27319
rect 2421 27081 2455 27115
rect 3709 27081 3743 27115
rect 6929 27081 6963 27115
rect 8033 27081 8067 27115
rect 11069 27081 11103 27115
rect 3065 27013 3099 27047
rect 9505 27013 9539 27047
rect 9597 27013 9631 27047
rect 12449 27013 12483 27047
rect 13737 27013 13771 27047
rect 13829 27013 13863 27047
rect 14565 27013 14599 27047
rect 15669 27013 15703 27047
rect 15761 27013 15795 27047
rect 17601 27013 17635 27047
rect 18981 27013 19015 27047
rect 20177 27013 20211 27047
rect 21281 27013 21315 27047
rect 22569 27013 22603 27047
rect 23397 27013 23431 27047
rect 1869 26945 1903 26979
rect 2329 26945 2363 26979
rect 2973 26945 3007 26979
rect 3801 26945 3835 26979
rect 7941 26945 7975 26979
rect 10333 26945 10367 26979
rect 10977 26945 11011 26979
rect 16313 26945 16347 26979
rect 21373 26945 21407 26979
rect 22017 26945 22051 26979
rect 38025 26945 38059 26979
rect 9321 26877 9355 26911
rect 11897 26877 11931 26911
rect 12541 26877 12575 26911
rect 14473 26877 14507 26911
rect 17693 26877 17727 26911
rect 18429 26877 18463 26911
rect 19073 26877 19107 26911
rect 20269 26877 20303 26911
rect 22661 26877 22695 26911
rect 23305 26877 23339 26911
rect 23581 26877 23615 26911
rect 7481 26809 7515 26843
rect 13277 26809 13311 26843
rect 15025 26809 15059 26843
rect 17141 26809 17175 26843
rect 19717 26809 19751 26843
rect 1685 26741 1719 26775
rect 4353 26741 4387 26775
rect 4905 26741 4939 26775
rect 5365 26741 5399 26775
rect 5917 26741 5951 26775
rect 10425 26741 10459 26775
rect 38209 26741 38243 26775
rect 1961 26537 1995 26571
rect 2605 26537 2639 26571
rect 3249 26537 3283 26571
rect 7113 26537 7147 26571
rect 8493 26537 8527 26571
rect 12541 26537 12575 26571
rect 16221 26537 16255 26571
rect 18061 26537 18095 26571
rect 22661 26537 22695 26571
rect 23305 26537 23339 26571
rect 29837 26537 29871 26571
rect 15577 26469 15611 26503
rect 16865 26469 16899 26503
rect 18797 26469 18831 26503
rect 20085 26469 20119 26503
rect 4997 26401 5031 26435
rect 7849 26401 7883 26435
rect 10701 26401 10735 26435
rect 11345 26401 11379 26435
rect 14473 26401 14507 26435
rect 17417 26401 17451 26435
rect 19522 26401 19556 26435
rect 21557 26401 21591 26435
rect 1869 26333 1903 26367
rect 2697 26333 2731 26367
rect 3157 26333 3191 26367
rect 6101 26333 6135 26367
rect 7297 26333 7331 26367
rect 7941 26333 7975 26367
rect 8401 26333 8435 26367
rect 11989 26333 12023 26367
rect 16129 26333 16163 26367
rect 18797 26333 18831 26367
rect 20913 26333 20947 26367
rect 22753 26333 22787 26367
rect 23213 26333 23247 26367
rect 24593 26333 24627 26367
rect 29929 26333 29963 26367
rect 4445 26265 4479 26299
rect 5549 26265 5583 26299
rect 9229 26265 9263 26299
rect 9321 26265 9355 26299
rect 10241 26265 10275 26299
rect 11437 26265 11471 26299
rect 13093 26265 13127 26299
rect 13185 26265 13219 26299
rect 13737 26265 13771 26299
rect 15025 26265 15059 26299
rect 15117 26265 15151 26299
rect 17325 26265 17359 26299
rect 19625 26265 19659 26299
rect 21465 26265 21499 26299
rect 23857 26265 23891 26299
rect 6653 26197 6687 26231
rect 1961 25993 1995 26027
rect 2605 25993 2639 26027
rect 6653 25993 6687 26027
rect 7849 25993 7883 26027
rect 11805 25993 11839 26027
rect 17233 25993 17267 26027
rect 17877 25993 17911 26027
rect 18521 25993 18555 26027
rect 20729 25993 20763 26027
rect 21373 25993 21407 26027
rect 9229 25925 9263 25959
rect 10609 25925 10643 25959
rect 11161 25925 11195 25959
rect 12541 25925 12575 25959
rect 13737 25925 13771 25959
rect 14289 25925 14323 25959
rect 14749 25925 14783 25959
rect 15301 25925 15335 25959
rect 15393 25925 15427 25959
rect 19257 25925 19291 25959
rect 22569 25925 22603 25959
rect 23305 25925 23339 25959
rect 1869 25857 1903 25891
rect 2513 25857 2547 25891
rect 5825 25857 5859 25891
rect 7113 25857 7147 25891
rect 7757 25857 7791 25891
rect 8401 25857 8435 25891
rect 11713 25857 11747 25891
rect 16313 25857 16347 25891
rect 17141 25857 17175 25891
rect 17969 25857 18003 25891
rect 18429 25857 18463 25891
rect 20637 25857 20671 25891
rect 21465 25857 21499 25891
rect 23397 25857 23431 25891
rect 23857 25857 23891 25891
rect 3709 25789 3743 25823
rect 9137 25789 9171 25823
rect 10517 25789 10551 25823
rect 12449 25789 12483 25823
rect 13645 25789 13679 25823
rect 19165 25789 19199 25823
rect 20177 25789 20211 25823
rect 22661 25789 22695 25823
rect 4813 25721 4847 25755
rect 5917 25721 5951 25755
rect 9689 25721 9723 25755
rect 13001 25721 13035 25755
rect 22109 25721 22143 25755
rect 4261 25653 4295 25687
rect 5365 25653 5399 25687
rect 7205 25653 7239 25687
rect 8493 25653 8527 25687
rect 16221 25653 16255 25687
rect 2237 25449 2271 25483
rect 2789 25449 2823 25483
rect 4997 25449 5031 25483
rect 5549 25449 5583 25483
rect 7297 25449 7331 25483
rect 9321 25449 9355 25483
rect 21465 25449 21499 25483
rect 29837 25449 29871 25483
rect 6745 25313 6779 25347
rect 7941 25313 7975 25347
rect 10241 25313 10275 25347
rect 11529 25313 11563 25347
rect 13093 25313 13127 25347
rect 15301 25313 15335 25347
rect 15945 25313 15979 25347
rect 16497 25313 16531 25347
rect 16773 25313 16807 25347
rect 18613 25313 18647 25347
rect 7205 25245 7239 25279
rect 9229 25245 9263 25279
rect 14381 25245 14415 25279
rect 19441 25245 19475 25279
rect 21557 25245 21591 25279
rect 22109 25245 22143 25279
rect 29929 25245 29963 25279
rect 1777 25177 1811 25211
rect 10425 25177 10459 25211
rect 10517 25177 10551 25211
rect 11630 25177 11664 25211
rect 12173 25177 12207 25211
rect 13185 25177 13219 25211
rect 13737 25177 13771 25211
rect 15393 25177 15427 25211
rect 16589 25177 16623 25211
rect 17969 25177 18003 25211
rect 18521 25177 18555 25211
rect 20269 25177 20303 25211
rect 20361 25177 20395 25211
rect 20913 25177 20947 25211
rect 23029 25177 23063 25211
rect 23121 25177 23155 25211
rect 24041 25177 24075 25211
rect 3433 25109 3467 25143
rect 4537 25109 4571 25143
rect 6193 25109 6227 25143
rect 8585 25109 8619 25143
rect 14473 25109 14507 25143
rect 19533 25109 19567 25143
rect 38301 25109 38335 25143
rect 4721 24905 4755 24939
rect 9873 24905 9907 24939
rect 18337 24905 18371 24939
rect 22753 24905 22787 24939
rect 23213 24905 23247 24939
rect 10609 24837 10643 24871
rect 11805 24837 11839 24871
rect 11897 24837 11931 24871
rect 13093 24837 13127 24871
rect 14473 24837 14507 24871
rect 19441 24837 19475 24871
rect 20269 24837 20303 24871
rect 1593 24769 1627 24803
rect 2237 24769 2271 24803
rect 2881 24769 2915 24803
rect 3433 24769 3467 24803
rect 5733 24769 5767 24803
rect 6561 24769 6595 24803
rect 7849 24769 7883 24803
rect 7941 24769 7975 24803
rect 8493 24769 8527 24803
rect 9137 24769 9171 24803
rect 9229 24769 9263 24803
rect 9781 24769 9815 24803
rect 13645 24769 13679 24803
rect 16313 24769 16347 24803
rect 17601 24769 17635 24803
rect 18429 24769 18463 24803
rect 21281 24769 21315 24803
rect 21373 24769 21407 24803
rect 29561 24769 29595 24803
rect 5825 24701 5859 24735
rect 10517 24701 10551 24735
rect 11161 24701 11195 24735
rect 13001 24701 13035 24735
rect 14381 24701 14415 24735
rect 15393 24701 15427 24735
rect 17141 24701 17175 24735
rect 17693 24701 17727 24735
rect 19533 24701 19567 24735
rect 20177 24701 20211 24735
rect 22017 24701 22051 24735
rect 38025 24701 38059 24735
rect 38301 24701 38335 24735
rect 1777 24633 1811 24667
rect 6653 24633 6687 24667
rect 8585 24633 8619 24667
rect 12357 24633 12391 24667
rect 18981 24633 19015 24667
rect 20729 24633 20763 24667
rect 23765 24633 23799 24667
rect 4169 24565 4203 24599
rect 5181 24565 5215 24599
rect 7389 24565 7423 24599
rect 16221 24565 16255 24599
rect 29653 24565 29687 24599
rect 1685 24361 1719 24395
rect 3341 24361 3375 24395
rect 4905 24361 4939 24395
rect 7113 24361 7147 24395
rect 8493 24361 8527 24395
rect 23029 24361 23063 24395
rect 33609 24361 33643 24395
rect 2237 24293 2271 24327
rect 5457 24293 5491 24327
rect 9321 24293 9355 24327
rect 15301 24293 15335 24327
rect 10241 24225 10275 24259
rect 10517 24225 10551 24259
rect 12357 24225 12391 24259
rect 17417 24225 17451 24259
rect 20729 24225 20763 24259
rect 21281 24225 21315 24259
rect 21925 24225 21959 24259
rect 22201 24225 22235 24259
rect 7297 24157 7331 24191
rect 7757 24157 7791 24191
rect 8401 24157 8435 24191
rect 9229 24157 9263 24191
rect 11069 24157 11103 24191
rect 19441 24157 19475 24191
rect 19993 24157 20027 24191
rect 20821 24157 20855 24191
rect 33793 24157 33827 24191
rect 34253 24157 34287 24191
rect 37841 24157 37875 24191
rect 6101 24089 6135 24123
rect 10425 24089 10459 24123
rect 11713 24089 11747 24123
rect 12265 24089 12299 24123
rect 13093 24089 13127 24123
rect 13185 24089 13219 24123
rect 13737 24089 13771 24123
rect 14749 24089 14783 24123
rect 14841 24089 14875 24123
rect 16405 24089 16439 24123
rect 16497 24089 16531 24123
rect 18613 24089 18647 24123
rect 20085 24089 20119 24123
rect 22017 24089 22051 24123
rect 2697 24021 2731 24055
rect 4353 24021 4387 24055
rect 6653 24021 6687 24055
rect 7849 24021 7883 24055
rect 11161 24021 11195 24055
rect 17969 24021 18003 24055
rect 18521 24021 18555 24055
rect 38025 24021 38059 24055
rect 2421 23817 2455 23851
rect 2973 23817 3007 23851
rect 3893 23817 3927 23851
rect 5181 23817 5215 23851
rect 5917 23817 5951 23851
rect 7849 23817 7883 23851
rect 11069 23817 11103 23851
rect 22017 23817 22051 23851
rect 26249 23817 26283 23851
rect 27261 23817 27295 23851
rect 30021 23817 30055 23851
rect 10425 23749 10459 23783
rect 12725 23749 12759 23783
rect 13277 23749 13311 23783
rect 13921 23749 13955 23783
rect 15393 23749 15427 23783
rect 16313 23749 16347 23783
rect 17325 23749 17359 23783
rect 17417 23749 17451 23783
rect 18981 23749 19015 23783
rect 19717 23749 19751 23783
rect 21189 23749 21223 23783
rect 1961 23681 1995 23715
rect 7757 23681 7791 23715
rect 9045 23681 9079 23715
rect 9689 23681 9723 23715
rect 10333 23681 10367 23715
rect 10977 23681 11011 23715
rect 11897 23681 11931 23715
rect 19809 23681 19843 23715
rect 26341 23681 26375 23715
rect 30113 23681 30147 23715
rect 30665 23681 30699 23715
rect 38025 23681 38059 23715
rect 7205 23613 7239 23647
rect 8585 23613 8619 23647
rect 9781 23613 9815 23647
rect 12633 23613 12667 23647
rect 13829 23613 13863 23647
rect 15301 23613 15335 23647
rect 19073 23613 19107 23647
rect 6745 23545 6779 23579
rect 14381 23545 14415 23579
rect 17877 23545 17911 23579
rect 18521 23545 18555 23579
rect 1777 23477 1811 23511
rect 4629 23477 4663 23511
rect 9137 23477 9171 23511
rect 11989 23477 12023 23511
rect 20729 23477 20763 23511
rect 38209 23477 38243 23511
rect 1685 23273 1719 23307
rect 2697 23273 2731 23307
rect 3249 23273 3283 23307
rect 7021 23273 7055 23307
rect 8493 23273 8527 23307
rect 13645 23273 13679 23307
rect 16221 23273 16255 23307
rect 18061 23273 18095 23307
rect 9965 23205 9999 23239
rect 13001 23205 13035 23239
rect 15577 23205 15611 23239
rect 18705 23205 18739 23239
rect 9413 23137 9447 23171
rect 10609 23137 10643 23171
rect 11253 23137 11287 23171
rect 14381 23137 14415 23171
rect 17141 23137 17175 23171
rect 21557 23137 21591 23171
rect 7665 23069 7699 23103
rect 8401 23069 8435 23103
rect 13461 23069 13495 23103
rect 15669 23069 15703 23103
rect 16313 23069 16347 23103
rect 18153 23069 18187 23103
rect 18797 23069 18831 23103
rect 19625 23069 19659 23103
rect 20913 23069 20947 23103
rect 29929 23069 29963 23103
rect 30573 23069 30607 23103
rect 2237 23001 2271 23035
rect 4353 23001 4387 23035
rect 6101 23001 6135 23035
rect 9505 23001 9539 23035
rect 10701 23001 10735 23035
rect 11805 23001 11839 23035
rect 11897 23001 11931 23035
rect 12449 23001 12483 23035
rect 14473 23001 14507 23035
rect 15025 23001 15059 23035
rect 17325 23001 17359 23035
rect 17417 23001 17451 23035
rect 19533 23001 19567 23035
rect 21097 23001 21131 23035
rect 4905 22933 4939 22967
rect 5549 22933 5583 22967
rect 7573 22933 7607 22967
rect 20085 22933 20119 22967
rect 30113 22933 30147 22967
rect 2329 22729 2363 22763
rect 3801 22729 3835 22763
rect 5457 22729 5491 22763
rect 8677 22729 8711 22763
rect 9965 22729 9999 22763
rect 13093 22729 13127 22763
rect 18061 22729 18095 22763
rect 4905 22661 4939 22695
rect 7573 22661 7607 22695
rect 11897 22661 11931 22695
rect 14197 22661 14231 22695
rect 14933 22661 14967 22695
rect 15025 22661 15059 22695
rect 16129 22661 16163 22695
rect 18981 22661 19015 22695
rect 19533 22661 19567 22695
rect 20177 22661 20211 22695
rect 20729 22661 20763 22695
rect 1869 22593 1903 22627
rect 2513 22593 2547 22627
rect 8585 22593 8619 22627
rect 9413 22593 9447 22627
rect 9873 22593 9907 22627
rect 13001 22593 13035 22627
rect 16221 22593 16255 22627
rect 17601 22593 17635 22627
rect 18245 22593 18279 22627
rect 2973 22525 3007 22559
rect 8125 22525 8159 22559
rect 10517 22525 10551 22559
rect 10701 22525 10735 22559
rect 11805 22525 11839 22559
rect 12081 22525 12115 22559
rect 14013 22525 14047 22559
rect 14289 22525 14323 22559
rect 16957 22525 16991 22559
rect 18889 22525 18923 22559
rect 20085 22525 20119 22559
rect 1685 22457 1719 22491
rect 9229 22457 9263 22491
rect 15485 22457 15519 22491
rect 6009 22389 6043 22423
rect 6837 22389 6871 22423
rect 11069 22389 11103 22423
rect 17509 22389 17543 22423
rect 38117 22389 38151 22423
rect 2421 22185 2455 22219
rect 8493 22185 8527 22219
rect 6469 22117 6503 22151
rect 11621 22117 11655 22151
rect 12357 22117 12391 22151
rect 1685 22049 1719 22083
rect 9229 22049 9263 22083
rect 13645 22049 13679 22083
rect 17877 22049 17911 22083
rect 18521 22049 18555 22083
rect 20545 22049 20579 22083
rect 21189 22049 21223 22083
rect 5457 21981 5491 22015
rect 5917 21981 5951 22015
rect 7297 21981 7331 22015
rect 8401 21981 8435 22015
rect 9781 21981 9815 22015
rect 9873 21981 9907 22015
rect 10333 21981 10367 22015
rect 12265 21981 12299 22015
rect 14565 21981 14599 22015
rect 17141 21981 17175 22015
rect 21097 21981 21131 22015
rect 21833 21981 21867 22015
rect 38025 21981 38059 22015
rect 7849 21913 7883 21947
rect 10425 21913 10459 21947
rect 11069 21913 11103 21947
rect 11161 21913 11195 21947
rect 13001 21913 13035 21947
rect 13093 21913 13127 21947
rect 15117 21913 15151 21947
rect 15209 21913 15243 21947
rect 15945 21913 15979 21947
rect 17969 21913 18003 21947
rect 3433 21845 3467 21879
rect 4077 21845 4111 21879
rect 4629 21845 4663 21879
rect 5273 21845 5307 21879
rect 16037 21845 16071 21879
rect 17049 21845 17083 21879
rect 19441 21845 19475 21879
rect 19993 21845 20027 21879
rect 37841 21845 37875 21879
rect 2513 21641 2547 21675
rect 3065 21641 3099 21675
rect 3617 21641 3651 21675
rect 4169 21641 4203 21675
rect 4721 21641 4755 21675
rect 6561 21641 6595 21675
rect 9505 21641 9539 21675
rect 18337 21641 18371 21675
rect 19901 21641 19935 21675
rect 5181 21573 5215 21607
rect 8861 21573 8895 21607
rect 10977 21573 11011 21607
rect 12357 21573 12391 21607
rect 14289 21573 14323 21607
rect 14381 21573 14415 21607
rect 15577 21573 15611 21607
rect 17141 21573 17175 21607
rect 1869 21505 1903 21539
rect 8125 21505 8159 21539
rect 8769 21505 8803 21539
rect 9413 21505 9447 21539
rect 17233 21505 17267 21539
rect 18429 21505 18463 21539
rect 19809 21505 19843 21539
rect 20453 21505 20487 21539
rect 38025 21505 38059 21539
rect 7573 21437 7607 21471
rect 10057 21437 10091 21471
rect 11069 21437 11103 21471
rect 12265 21437 12299 21471
rect 14105 21437 14139 21471
rect 15025 21437 15059 21471
rect 15669 21437 15703 21471
rect 8217 21369 8251 21403
rect 12817 21369 12851 21403
rect 16313 21369 16347 21403
rect 18889 21369 18923 21403
rect 1685 21301 1719 21335
rect 17693 21301 17727 21335
rect 38209 21301 38243 21335
rect 2237 21097 2271 21131
rect 2789 21097 2823 21131
rect 4077 21097 4111 21131
rect 4537 21097 4571 21131
rect 8493 21097 8527 21131
rect 9597 21097 9631 21131
rect 11437 21097 11471 21131
rect 10241 21029 10275 21063
rect 18061 21029 18095 21063
rect 3433 20961 3467 20995
rect 12541 20961 12575 20995
rect 13737 20961 13771 20995
rect 14749 20961 14783 20995
rect 15393 20961 15427 20995
rect 16773 20961 16807 20995
rect 9505 20893 9539 20927
rect 12357 20893 12391 20927
rect 16229 20893 16263 20927
rect 16865 20893 16899 20927
rect 17509 20893 17543 20927
rect 18797 20893 18831 20927
rect 19441 20893 19475 20927
rect 10701 20825 10735 20859
rect 10793 20825 10827 20859
rect 13093 20825 13127 20859
rect 13185 20825 13219 20859
rect 15301 20825 15335 20859
rect 11897 20757 11931 20791
rect 16129 20757 16163 20791
rect 17325 20757 17359 20791
rect 18705 20757 18739 20791
rect 3617 20553 3651 20587
rect 9873 20553 9907 20587
rect 11805 20553 11839 20587
rect 13553 20553 13587 20587
rect 15393 20553 15427 20587
rect 16957 20553 16991 20587
rect 17509 20553 17543 20587
rect 18705 20553 18739 20587
rect 10977 20485 11011 20519
rect 12265 20485 12299 20519
rect 12817 20485 12851 20519
rect 14289 20485 14323 20519
rect 16037 20485 16071 20519
rect 9781 20417 9815 20451
rect 13461 20417 13495 20451
rect 15485 20417 15519 20451
rect 15945 20417 15979 20451
rect 17049 20417 17083 20451
rect 37841 20417 37875 20451
rect 10793 20349 10827 20383
rect 11069 20349 11103 20383
rect 12909 20349 12943 20383
rect 14197 20349 14231 20383
rect 14473 20349 14507 20383
rect 9321 20213 9355 20247
rect 18061 20213 18095 20247
rect 38025 20213 38059 20247
rect 9321 20009 9355 20043
rect 9873 20009 9907 20043
rect 14289 20009 14323 20043
rect 16129 20009 16163 20043
rect 16957 20009 16991 20043
rect 21465 20009 21499 20043
rect 12357 19941 12391 19975
rect 11805 19873 11839 19907
rect 13737 19873 13771 19907
rect 15485 19873 15519 19907
rect 17509 19873 17543 19907
rect 22293 19873 22327 19907
rect 7297 19805 7331 19839
rect 9781 19805 9815 19839
rect 10425 19805 10459 19839
rect 11069 19805 11103 19839
rect 16037 19805 16071 19839
rect 22109 19805 22143 19839
rect 38025 19805 38059 19839
rect 10517 19737 10551 19771
rect 11897 19737 11931 19771
rect 13093 19737 13127 19771
rect 13185 19737 13219 19771
rect 14841 19737 14875 19771
rect 15393 19737 15427 19771
rect 18061 19737 18095 19771
rect 7205 19669 7239 19703
rect 11161 19669 11195 19703
rect 38209 19669 38243 19703
rect 10517 19465 10551 19499
rect 11069 19465 11103 19499
rect 11989 19465 12023 19499
rect 13553 19465 13587 19499
rect 16221 19465 16255 19499
rect 14197 19397 14231 19431
rect 14289 19397 14323 19431
rect 15577 19397 15611 19431
rect 1869 19329 1903 19363
rect 11161 19329 11195 19363
rect 12633 19329 12667 19363
rect 13645 19329 13679 19363
rect 15485 19329 15519 19363
rect 16313 19329 16347 19363
rect 9965 19261 9999 19295
rect 12449 19261 12483 19295
rect 14841 19261 14875 19295
rect 16957 19193 16991 19227
rect 17417 19193 17451 19227
rect 1685 19125 1719 19159
rect 4721 18921 4755 18955
rect 10149 18921 10183 18955
rect 10701 18921 10735 18955
rect 12725 18921 12759 18955
rect 13461 18921 13495 18955
rect 14565 18921 14599 18955
rect 15209 18921 15243 18955
rect 15945 18921 15979 18955
rect 16497 18921 16531 18955
rect 12173 18853 12207 18887
rect 4169 18717 4203 18751
rect 12817 18717 12851 18751
rect 13553 18717 13587 18751
rect 14657 18717 14691 18751
rect 15301 18717 15335 18751
rect 3985 18581 4019 18615
rect 11529 18581 11563 18615
rect 2421 18377 2455 18411
rect 13001 18377 13035 18411
rect 13645 18377 13679 18411
rect 14565 18377 14599 18411
rect 15853 18377 15887 18411
rect 12449 18309 12483 18343
rect 15301 18309 15335 18343
rect 1869 18241 1903 18275
rect 4721 18241 4755 18275
rect 13093 18241 13127 18275
rect 13737 18241 13771 18275
rect 14657 18241 14691 18275
rect 11805 18173 11839 18207
rect 1685 18037 1719 18071
rect 4629 18037 4663 18071
rect 13001 17833 13035 17867
rect 15485 17833 15519 17867
rect 14841 17697 14875 17731
rect 30297 17629 30331 17663
rect 13737 17561 13771 17595
rect 14381 17561 14415 17595
rect 14473 17561 14507 17595
rect 30205 17493 30239 17527
rect 13921 17289 13955 17323
rect 14565 17289 14599 17323
rect 15209 17289 15243 17323
rect 14657 17153 14691 17187
rect 25053 17153 25087 17187
rect 25697 17153 25731 17187
rect 25789 16949 25823 16983
rect 21833 16609 21867 16643
rect 21189 16541 21223 16575
rect 21281 16541 21315 16575
rect 1869 16065 1903 16099
rect 38025 16065 38059 16099
rect 1685 15861 1719 15895
rect 38209 15861 38243 15895
rect 38025 14433 38059 14467
rect 38301 14365 38335 14399
rect 38301 14025 38335 14059
rect 1869 13889 1903 13923
rect 1685 13685 1719 13719
rect 13277 13481 13311 13515
rect 20453 13481 20487 13515
rect 13369 13277 13403 13311
rect 19717 13277 19751 13311
rect 19901 13141 19935 13175
rect 16957 12937 16991 12971
rect 1869 12801 1903 12835
rect 16313 12801 16347 12835
rect 38025 12801 38059 12835
rect 37473 12733 37507 12767
rect 1685 12597 1719 12631
rect 16129 12597 16163 12631
rect 38209 12597 38243 12631
rect 15669 12325 15703 12359
rect 15485 12189 15519 12223
rect 16129 12189 16163 12223
rect 37841 12189 37875 12223
rect 38025 12053 38059 12087
rect 24409 11849 24443 11883
rect 24501 11713 24535 11747
rect 24961 11509 24995 11543
rect 37565 11101 37599 11135
rect 38025 11033 38059 11067
rect 38209 11033 38243 11067
rect 13185 10761 13219 10795
rect 2421 10693 2455 10727
rect 1869 10625 1903 10659
rect 13277 10625 13311 10659
rect 1685 10421 1719 10455
rect 13829 10421 13863 10455
rect 9873 10217 9907 10251
rect 12725 10217 12759 10251
rect 9781 10013 9815 10047
rect 13461 10013 13495 10047
rect 13277 9877 13311 9911
rect 20729 9605 20763 9639
rect 21281 9537 21315 9571
rect 21373 9333 21407 9367
rect 38025 8925 38059 8959
rect 1685 8857 1719 8891
rect 1777 8789 1811 8823
rect 38209 8789 38243 8823
rect 1685 8585 1719 8619
rect 1869 7429 1903 7463
rect 38025 7429 38059 7463
rect 1685 7361 1719 7395
rect 37565 7361 37599 7395
rect 38209 7361 38243 7395
rect 1593 6953 1627 6987
rect 7297 6817 7331 6851
rect 6745 6749 6779 6783
rect 23673 6749 23707 6783
rect 6653 6613 6687 6647
rect 23857 6613 23891 6647
rect 24685 6613 24719 6647
rect 32965 6409 32999 6443
rect 32321 6273 32355 6307
rect 32413 6137 32447 6171
rect 38025 5797 38059 5831
rect 37565 5593 37599 5627
rect 38209 5593 38243 5627
rect 1777 5321 1811 5355
rect 1685 5185 1719 5219
rect 1593 4777 1627 4811
rect 1869 3485 1903 3519
rect 38025 3485 38059 3519
rect 2421 3417 2455 3451
rect 1685 3349 1719 3383
rect 37473 3349 37507 3383
rect 38209 3349 38243 3383
rect 5733 3145 5767 3179
rect 35081 3145 35115 3179
rect 34621 3077 34655 3111
rect 1685 3009 1719 3043
rect 2881 3009 2915 3043
rect 8585 3009 8619 3043
rect 13461 3009 13495 3043
rect 19993 3009 20027 3043
rect 20637 3009 20671 3043
rect 33885 3009 33919 3043
rect 38025 3009 38059 3043
rect 13645 2941 13679 2975
rect 1869 2873 1903 2907
rect 20177 2873 20211 2907
rect 34069 2873 34103 2907
rect 2421 2805 2455 2839
rect 8401 2805 8435 2839
rect 29653 2805 29687 2839
rect 37565 2805 37599 2839
rect 38209 2805 38243 2839
rect 11897 2601 11931 2635
rect 18337 2601 18371 2635
rect 32413 2601 32447 2635
rect 33701 2601 33735 2635
rect 36737 2601 36771 2635
rect 37565 2601 37599 2635
rect 2605 2533 2639 2567
rect 15209 2533 15243 2567
rect 21373 2533 21407 2567
rect 23305 2533 23339 2567
rect 4261 2465 4295 2499
rect 30021 2465 30055 2499
rect 1869 2397 1903 2431
rect 3985 2397 4019 2431
rect 5549 2397 5583 2431
rect 6837 2397 6871 2431
rect 8309 2397 8343 2431
rect 9321 2397 9355 2431
rect 9781 2397 9815 2431
rect 10057 2397 10091 2431
rect 13277 2397 13311 2431
rect 16865 2397 16899 2431
rect 20085 2397 20119 2431
rect 22017 2397 22051 2431
rect 25237 2397 25271 2431
rect 27169 2397 27203 2431
rect 28457 2397 28491 2431
rect 29745 2397 29779 2431
rect 35173 2397 35207 2431
rect 35909 2397 35943 2431
rect 37657 2397 37691 2431
rect 38209 2397 38243 2431
rect 2421 2329 2455 2363
rect 7389 2329 7423 2363
rect 11161 2329 11195 2363
rect 11805 2329 11839 2363
rect 14473 2329 14507 2363
rect 15025 2329 15059 2363
rect 17693 2329 17727 2363
rect 18245 2329 18279 2363
rect 22845 2329 22879 2363
rect 23489 2329 23523 2363
rect 32505 2329 32539 2363
rect 33149 2329 33183 2363
rect 33793 2329 33827 2363
rect 36829 2329 36863 2363
rect 1685 2261 1719 2295
rect 3341 2261 3375 2295
rect 5365 2261 5399 2295
rect 6653 2261 6687 2295
rect 8493 2261 8527 2295
rect 13093 2261 13127 2295
rect 17049 2261 17083 2295
rect 20269 2261 20303 2295
rect 22201 2261 22235 2295
rect 25421 2261 25455 2295
rect 27353 2261 27387 2295
rect 28641 2261 28675 2295
rect 31769 2261 31803 2295
rect 34989 2261 35023 2295
rect 36093 2261 36127 2295
<< metal1 >>
rect 4798 37748 4804 37800
rect 4856 37788 4862 37800
rect 16666 37788 16672 37800
rect 4856 37760 16672 37788
rect 4856 37748 4862 37760
rect 16666 37748 16672 37760
rect 16724 37748 16730 37800
rect 10594 37680 10600 37732
rect 10652 37720 10658 37732
rect 22738 37720 22744 37732
rect 10652 37692 22744 37720
rect 10652 37680 10658 37692
rect 22738 37680 22744 37692
rect 22796 37680 22802 37732
rect 14 37612 20 37664
rect 72 37652 78 37664
rect 4890 37652 4896 37664
rect 72 37624 4896 37652
rect 72 37612 78 37624
rect 4890 37612 4896 37624
rect 4948 37612 4954 37664
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 10226 37448 10232 37460
rect 9600 37420 10232 37448
rect 3142 37312 3148 37324
rect 3103 37284 3148 37312
rect 3142 37272 3148 37284
rect 3200 37272 3206 37324
rect 3421 37315 3479 37321
rect 3421 37281 3433 37315
rect 3467 37312 3479 37315
rect 3878 37312 3884 37324
rect 3467 37284 3884 37312
rect 3467 37281 3479 37284
rect 3421 37275 3479 37281
rect 3878 37272 3884 37284
rect 3936 37312 3942 37324
rect 4157 37315 4215 37321
rect 4157 37312 4169 37315
rect 3936 37284 4169 37312
rect 3936 37272 3942 37284
rect 4157 37281 4169 37284
rect 4203 37281 4215 37315
rect 4157 37275 4215 37281
rect 4433 37315 4491 37321
rect 4433 37281 4445 37315
rect 4479 37312 4491 37315
rect 4798 37312 4804 37324
rect 4479 37284 4804 37312
rect 4479 37281 4491 37284
rect 4433 37275 4491 37281
rect 4798 37272 4804 37284
rect 4856 37272 4862 37324
rect 8297 37315 8355 37321
rect 8297 37281 8309 37315
rect 8343 37312 8355 37315
rect 9600 37312 9628 37420
rect 10226 37408 10232 37420
rect 10284 37448 10290 37460
rect 10594 37448 10600 37460
rect 10284 37420 10600 37448
rect 10284 37408 10290 37420
rect 10594 37408 10600 37420
rect 10652 37408 10658 37460
rect 20530 37448 20536 37460
rect 13740 37420 20536 37448
rect 8343 37284 9628 37312
rect 8343 37281 8355 37284
rect 8297 37275 8355 37281
rect 9858 37272 9864 37324
rect 9916 37312 9922 37324
rect 10597 37315 10655 37321
rect 10597 37312 10609 37315
rect 9916 37284 10609 37312
rect 9916 37272 9922 37284
rect 10597 37281 10609 37284
rect 10643 37312 10655 37315
rect 10962 37312 10968 37324
rect 10643 37284 10968 37312
rect 10643 37281 10655 37284
rect 10597 37275 10655 37281
rect 10962 37272 10968 37284
rect 11020 37272 11026 37324
rect 11701 37315 11759 37321
rect 11701 37281 11713 37315
rect 11747 37312 11759 37315
rect 12618 37312 12624 37324
rect 11747 37284 12624 37312
rect 11747 37281 11759 37284
rect 11701 37275 11759 37281
rect 2038 37204 2044 37256
rect 2096 37204 2102 37256
rect 5534 37204 5540 37256
rect 5592 37204 5598 37256
rect 8573 37247 8631 37253
rect 8573 37213 8585 37247
rect 8619 37244 8631 37247
rect 8938 37244 8944 37256
rect 8619 37216 8944 37244
rect 8619 37213 8631 37216
rect 8573 37207 8631 37213
rect 8938 37204 8944 37216
rect 8996 37204 9002 37256
rect 10873 37247 10931 37253
rect 10873 37213 10885 37247
rect 10919 37244 10931 37247
rect 11514 37244 11520 37256
rect 10919 37216 11520 37244
rect 10919 37213 10931 37216
rect 10873 37207 10931 37213
rect 11514 37204 11520 37216
rect 11572 37204 11578 37256
rect 11716 37244 11744 37275
rect 12618 37272 12624 37284
rect 12676 37272 12682 37324
rect 13173 37315 13231 37321
rect 13173 37281 13185 37315
rect 13219 37312 13231 37315
rect 13740 37312 13768 37420
rect 20530 37408 20536 37420
rect 20588 37408 20594 37460
rect 22738 37448 22744 37460
rect 22699 37420 22744 37448
rect 22738 37408 22744 37420
rect 22796 37408 22802 37460
rect 23842 37408 23848 37460
rect 23900 37448 23906 37460
rect 23937 37451 23995 37457
rect 23937 37448 23949 37451
rect 23900 37420 23949 37448
rect 23900 37408 23906 37420
rect 23937 37417 23949 37420
rect 23983 37417 23995 37451
rect 36722 37448 36728 37460
rect 36683 37420 36728 37448
rect 23937 37411 23995 37417
rect 36722 37408 36728 37420
rect 36780 37408 36786 37460
rect 20165 37383 20223 37389
rect 20165 37380 20177 37383
rect 15120 37352 20177 37380
rect 13219 37284 13768 37312
rect 13219 37281 13231 37284
rect 13173 37275 13231 37281
rect 13814 37272 13820 37324
rect 13872 37312 13878 37324
rect 15120 37321 15148 37352
rect 20165 37349 20177 37352
rect 20211 37349 20223 37383
rect 32398 37380 32404 37392
rect 20165 37343 20223 37349
rect 26206 37352 32404 37380
rect 15105 37315 15163 37321
rect 15105 37312 15117 37315
rect 13872 37284 15117 37312
rect 13872 37272 13878 37284
rect 15105 37281 15117 37284
rect 15151 37281 15163 37315
rect 16850 37312 16856 37324
rect 16811 37284 16856 37312
rect 15105 37275 15163 37281
rect 16850 37272 16856 37284
rect 16908 37272 16914 37324
rect 18598 37272 18604 37324
rect 18656 37312 18662 37324
rect 18693 37315 18751 37321
rect 18693 37312 18705 37315
rect 18656 37284 18705 37312
rect 18656 37272 18662 37284
rect 18693 37281 18705 37284
rect 18739 37312 18751 37315
rect 26206 37312 26234 37352
rect 32398 37340 32404 37352
rect 32456 37340 32462 37392
rect 18739 37284 26234 37312
rect 29917 37315 29975 37321
rect 18739 37281 18751 37284
rect 18693 37275 18751 37281
rect 29917 37281 29929 37315
rect 29963 37312 29975 37315
rect 30282 37312 30288 37324
rect 29963 37284 30288 37312
rect 29963 37281 29975 37284
rect 29917 37275 29975 37281
rect 30282 37272 30288 37284
rect 30340 37312 30346 37324
rect 30377 37315 30435 37321
rect 30377 37312 30389 37315
rect 30340 37284 30389 37312
rect 30340 37272 30346 37284
rect 30377 37281 30389 37284
rect 30423 37281 30435 37315
rect 30377 37275 30435 37281
rect 11624 37216 11744 37244
rect 13449 37247 13507 37253
rect 3068 37148 3464 37176
rect 1673 37111 1731 37117
rect 1673 37077 1685 37111
rect 1719 37108 1731 37111
rect 3068 37108 3096 37148
rect 1719 37080 3096 37108
rect 3436 37108 3464 37148
rect 5718 37136 5724 37188
rect 5776 37176 5782 37188
rect 5776 37148 7052 37176
rect 5776 37136 5782 37148
rect 5810 37108 5816 37120
rect 3436 37080 5816 37108
rect 1719 37077 1731 37080
rect 1673 37071 1731 37077
rect 5810 37068 5816 37080
rect 5868 37068 5874 37120
rect 5905 37111 5963 37117
rect 5905 37077 5917 37111
rect 5951 37108 5963 37111
rect 6730 37108 6736 37120
rect 5951 37080 6736 37108
rect 5951 37077 5963 37080
rect 5905 37071 5963 37077
rect 6730 37068 6736 37080
rect 6788 37068 6794 37120
rect 6822 37068 6828 37120
rect 6880 37108 6886 37120
rect 7024 37108 7052 37148
rect 7834 37136 7840 37188
rect 7892 37136 7898 37188
rect 10686 37176 10692 37188
rect 9048 37148 9352 37176
rect 10166 37148 10692 37176
rect 9048 37108 9076 37148
rect 6880 37080 6925 37108
rect 7024 37080 9076 37108
rect 6880 37068 6886 37080
rect 9122 37068 9128 37120
rect 9180 37108 9186 37120
rect 9324 37108 9352 37148
rect 10686 37136 10692 37148
rect 10744 37136 10750 37188
rect 11624 37108 11652 37216
rect 13449 37213 13461 37247
rect 13495 37244 13507 37247
rect 13722 37244 13728 37256
rect 13495 37216 13728 37244
rect 13495 37213 13507 37216
rect 13449 37207 13507 37213
rect 13722 37204 13728 37216
rect 13780 37204 13786 37256
rect 14829 37247 14887 37253
rect 14829 37213 14841 37247
rect 14875 37213 14887 37247
rect 15838 37244 15844 37256
rect 15799 37216 15844 37244
rect 14829 37207 14887 37213
rect 11698 37136 11704 37188
rect 11756 37176 11762 37188
rect 11756 37148 12006 37176
rect 11756 37136 11762 37148
rect 14642 37136 14648 37188
rect 14700 37176 14706 37188
rect 14844 37176 14872 37207
rect 15838 37204 15844 37216
rect 15896 37204 15902 37256
rect 16758 37204 16764 37256
rect 16816 37244 16822 37256
rect 17037 37247 17095 37253
rect 17037 37244 17049 37247
rect 16816 37216 17049 37244
rect 16816 37204 16822 37216
rect 17037 37213 17049 37216
rect 17083 37244 17095 37247
rect 17589 37247 17647 37253
rect 17589 37244 17601 37247
rect 17083 37216 17601 37244
rect 17083 37213 17095 37216
rect 17037 37207 17095 37213
rect 17589 37213 17601 37216
rect 17635 37213 17647 37247
rect 19426 37244 19432 37256
rect 19387 37216 19432 37244
rect 17589 37207 17647 37213
rect 19426 37204 19432 37216
rect 19484 37204 19490 37256
rect 20714 37204 20720 37256
rect 20772 37244 20778 37256
rect 20901 37247 20959 37253
rect 20901 37244 20913 37247
rect 20772 37216 20913 37244
rect 20772 37204 20778 37216
rect 20901 37213 20913 37216
rect 20947 37244 20959 37247
rect 21361 37247 21419 37253
rect 21361 37244 21373 37247
rect 20947 37216 21373 37244
rect 20947 37213 20959 37216
rect 20901 37207 20959 37213
rect 21361 37213 21373 37216
rect 21407 37213 21419 37247
rect 21361 37207 21419 37213
rect 21450 37204 21456 37256
rect 21508 37244 21514 37256
rect 22005 37247 22063 37253
rect 22005 37244 22017 37247
rect 21508 37216 22017 37244
rect 21508 37204 21514 37216
rect 22005 37213 22017 37216
rect 22051 37213 22063 37247
rect 22005 37207 22063 37213
rect 23842 37204 23848 37256
rect 23900 37244 23906 37256
rect 24765 37247 24823 37253
rect 24765 37244 24777 37247
rect 23900 37216 24777 37244
rect 23900 37204 23906 37216
rect 24765 37213 24777 37216
rect 24811 37213 24823 37247
rect 24765 37207 24823 37213
rect 25317 37247 25375 37253
rect 25317 37213 25329 37247
rect 25363 37213 25375 37247
rect 27157 37247 27215 37253
rect 27157 37244 27169 37247
rect 25317 37207 25375 37213
rect 26528 37216 27169 37244
rect 19978 37176 19984 37188
rect 14700 37148 19984 37176
rect 14700 37136 14706 37148
rect 19978 37136 19984 37148
rect 20036 37136 20042 37188
rect 23198 37136 23204 37188
rect 23256 37176 23262 37188
rect 25332 37176 25360 37207
rect 23256 37148 25360 37176
rect 23256 37136 23262 37148
rect 26528 37120 26556 37216
rect 27157 37213 27169 37216
rect 27203 37213 27215 37247
rect 28902 37244 28908 37256
rect 28863 37216 28908 37244
rect 27157 37207 27215 37213
rect 28902 37204 28908 37216
rect 28960 37204 28966 37256
rect 30650 37244 30656 37256
rect 30611 37216 30656 37244
rect 30650 37204 30656 37216
rect 30708 37204 30714 37256
rect 32309 37247 32367 37253
rect 32309 37244 32321 37247
rect 31772 37216 32321 37244
rect 31772 37120 31800 37216
rect 32309 37213 32321 37216
rect 32355 37213 32367 37247
rect 33594 37244 33600 37256
rect 33555 37216 33600 37244
rect 32309 37207 32367 37213
rect 33594 37204 33600 37216
rect 33652 37204 33658 37256
rect 35526 37244 35532 37256
rect 35487 37216 35532 37244
rect 35526 37204 35532 37216
rect 35584 37204 35590 37256
rect 36909 37247 36967 37253
rect 36909 37213 36921 37247
rect 36955 37244 36967 37247
rect 37366 37244 37372 37256
rect 36955 37216 37372 37244
rect 36955 37213 36967 37216
rect 36909 37207 36967 37213
rect 37366 37204 37372 37216
rect 37424 37204 37430 37256
rect 37461 37247 37519 37253
rect 37461 37213 37473 37247
rect 37507 37213 37519 37247
rect 37461 37207 37519 37213
rect 31846 37136 31852 37188
rect 31904 37176 31910 37188
rect 37476 37176 37504 37207
rect 31904 37148 37504 37176
rect 31904 37136 31910 37148
rect 9180 37080 9225 37108
rect 9324 37080 11652 37108
rect 9180 37068 9186 37080
rect 12894 37068 12900 37120
rect 12952 37108 12958 37120
rect 15194 37108 15200 37120
rect 12952 37080 15200 37108
rect 12952 37068 12958 37080
rect 15194 37068 15200 37080
rect 15252 37068 15258 37120
rect 15470 37068 15476 37120
rect 15528 37108 15534 37120
rect 15657 37111 15715 37117
rect 15657 37108 15669 37111
rect 15528 37080 15669 37108
rect 15528 37068 15534 37080
rect 15657 37077 15669 37080
rect 15703 37077 15715 37111
rect 15657 37071 15715 37077
rect 15746 37068 15752 37120
rect 15804 37108 15810 37120
rect 18141 37111 18199 37117
rect 18141 37108 18153 37111
rect 15804 37080 18153 37108
rect 15804 37068 15810 37080
rect 18141 37077 18153 37080
rect 18187 37108 18199 37111
rect 18506 37108 18512 37120
rect 18187 37080 18512 37108
rect 18187 37077 18199 37080
rect 18141 37071 18199 37077
rect 18506 37068 18512 37080
rect 18564 37068 18570 37120
rect 18782 37068 18788 37120
rect 18840 37108 18846 37120
rect 19613 37111 19671 37117
rect 19613 37108 19625 37111
rect 18840 37080 19625 37108
rect 18840 37068 18846 37080
rect 19613 37077 19625 37080
rect 19659 37077 19671 37111
rect 20714 37108 20720 37120
rect 20675 37080 20720 37108
rect 19613 37071 19671 37077
rect 20714 37068 20720 37080
rect 20772 37068 20778 37120
rect 22094 37068 22100 37120
rect 22152 37108 22158 37120
rect 22189 37111 22247 37117
rect 22189 37108 22201 37111
rect 22152 37080 22201 37108
rect 22152 37068 22158 37080
rect 22189 37077 22201 37080
rect 22235 37077 22247 37111
rect 23290 37108 23296 37120
rect 23251 37080 23296 37108
rect 22189 37071 22247 37077
rect 23290 37068 23296 37080
rect 23348 37068 23354 37120
rect 24670 37108 24676 37120
rect 24631 37080 24676 37108
rect 24670 37068 24676 37080
rect 24728 37068 24734 37120
rect 25130 37068 25136 37120
rect 25188 37108 25194 37120
rect 25501 37111 25559 37117
rect 25501 37108 25513 37111
rect 25188 37080 25513 37108
rect 25188 37068 25194 37080
rect 25501 37077 25513 37080
rect 25547 37077 25559 37111
rect 26510 37108 26516 37120
rect 26471 37080 26516 37108
rect 25501 37071 25559 37077
rect 26510 37068 26516 37080
rect 26568 37068 26574 37120
rect 27062 37068 27068 37120
rect 27120 37108 27126 37120
rect 27341 37111 27399 37117
rect 27341 37108 27353 37111
rect 27120 37080 27353 37108
rect 27120 37068 27126 37080
rect 27341 37077 27353 37080
rect 27387 37077 27399 37111
rect 27341 37071 27399 37077
rect 28994 37068 29000 37120
rect 29052 37108 29058 37120
rect 29089 37111 29147 37117
rect 29089 37108 29101 37111
rect 29052 37080 29101 37108
rect 29052 37068 29058 37080
rect 29089 37077 29101 37080
rect 29135 37077 29147 37111
rect 31754 37108 31760 37120
rect 31715 37080 31760 37108
rect 29089 37071 29147 37077
rect 31754 37068 31760 37080
rect 31812 37068 31818 37120
rect 32214 37068 32220 37120
rect 32272 37108 32278 37120
rect 32493 37111 32551 37117
rect 32493 37108 32505 37111
rect 32272 37080 32505 37108
rect 32272 37068 32278 37080
rect 32493 37077 32505 37080
rect 32539 37077 32551 37111
rect 32493 37071 32551 37077
rect 33502 37068 33508 37120
rect 33560 37108 33566 37120
rect 33781 37111 33839 37117
rect 33781 37108 33793 37111
rect 33560 37080 33793 37108
rect 33560 37068 33566 37080
rect 33781 37077 33793 37080
rect 33827 37077 33839 37111
rect 33781 37071 33839 37077
rect 35434 37068 35440 37120
rect 35492 37108 35498 37120
rect 35713 37111 35771 37117
rect 35713 37108 35725 37111
rect 35492 37080 35725 37108
rect 35492 37068 35498 37080
rect 35713 37077 35725 37080
rect 35759 37077 35771 37111
rect 35713 37071 35771 37077
rect 37458 37068 37464 37120
rect 37516 37108 37522 37120
rect 37645 37111 37703 37117
rect 37645 37108 37657 37111
rect 37516 37080 37657 37108
rect 37516 37068 37522 37080
rect 37645 37077 37657 37080
rect 37691 37077 37703 37111
rect 37645 37071 37703 37077
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 7834 36864 7840 36916
rect 7892 36904 7898 36916
rect 12526 36904 12532 36916
rect 7892 36876 12532 36904
rect 7892 36864 7898 36876
rect 12526 36864 12532 36876
rect 12584 36864 12590 36916
rect 12618 36864 12624 36916
rect 12676 36904 12682 36916
rect 15562 36904 15568 36916
rect 12676 36876 15568 36904
rect 12676 36864 12682 36876
rect 15562 36864 15568 36876
rect 15620 36864 15626 36916
rect 16025 36907 16083 36913
rect 16025 36873 16037 36907
rect 16071 36904 16083 36907
rect 21450 36904 21456 36916
rect 16071 36876 21456 36904
rect 16071 36873 16083 36876
rect 16025 36867 16083 36873
rect 21450 36864 21456 36876
rect 21508 36864 21514 36916
rect 30650 36904 30656 36916
rect 22066 36876 30656 36904
rect 1578 36796 1584 36848
rect 1636 36836 1642 36848
rect 2317 36839 2375 36845
rect 2317 36836 2329 36839
rect 1636 36808 2329 36836
rect 1636 36796 1642 36808
rect 2317 36805 2329 36808
rect 2363 36805 2375 36839
rect 3694 36836 3700 36848
rect 3542 36808 3700 36836
rect 2317 36799 2375 36805
rect 3694 36796 3700 36808
rect 3752 36796 3758 36848
rect 5718 36836 5724 36848
rect 5679 36808 5724 36836
rect 5718 36796 5724 36808
rect 5776 36796 5782 36848
rect 8662 36796 8668 36848
rect 8720 36836 8726 36848
rect 9122 36836 9128 36848
rect 8720 36808 9128 36836
rect 8720 36796 8726 36808
rect 9122 36796 9128 36808
rect 9180 36796 9186 36848
rect 9582 36796 9588 36848
rect 9640 36836 9646 36848
rect 9640 36808 9706 36836
rect 9640 36796 9646 36808
rect 10594 36796 10600 36848
rect 10652 36836 10658 36848
rect 10652 36808 11192 36836
rect 10652 36796 10658 36808
rect 1670 36728 1676 36780
rect 1728 36768 1734 36780
rect 2041 36771 2099 36777
rect 2041 36768 2053 36771
rect 1728 36740 2053 36768
rect 1728 36728 1734 36740
rect 2041 36737 2053 36740
rect 2087 36737 2099 36771
rect 6917 36771 6975 36777
rect 6917 36768 6929 36771
rect 2041 36731 2099 36737
rect 1302 36660 1308 36712
rect 1360 36700 1366 36712
rect 4632 36700 4660 36754
rect 6012 36740 6929 36768
rect 1360 36672 4660 36700
rect 1360 36660 1366 36672
rect 5350 36660 5356 36712
rect 5408 36700 5414 36712
rect 6012 36709 6040 36740
rect 5997 36703 6055 36709
rect 5997 36700 6009 36703
rect 5408 36672 6009 36700
rect 5408 36660 5414 36672
rect 5997 36669 6009 36672
rect 6043 36669 6055 36703
rect 5997 36663 6055 36669
rect 3326 36524 3332 36576
rect 3384 36564 3390 36576
rect 3789 36567 3847 36573
rect 3789 36564 3801 36567
rect 3384 36536 3801 36564
rect 3384 36524 3390 36536
rect 3789 36533 3801 36536
rect 3835 36533 3847 36567
rect 3789 36527 3847 36533
rect 4249 36567 4307 36573
rect 4249 36533 4261 36567
rect 4295 36564 4307 36567
rect 4614 36564 4620 36576
rect 4295 36536 4620 36564
rect 4295 36533 4307 36536
rect 4249 36527 4307 36533
rect 4614 36524 4620 36536
rect 4672 36524 4678 36576
rect 6748 36564 6776 36740
rect 6917 36737 6929 36740
rect 6963 36737 6975 36771
rect 8570 36768 8576 36780
rect 8326 36740 8576 36768
rect 6917 36731 6975 36737
rect 8570 36728 8576 36740
rect 8628 36728 8634 36780
rect 11164 36768 11192 36808
rect 11330 36796 11336 36848
rect 11388 36836 11394 36848
rect 11701 36839 11759 36845
rect 11701 36836 11713 36839
rect 11388 36808 11713 36836
rect 11388 36796 11394 36808
rect 11701 36805 11713 36808
rect 11747 36805 11759 36839
rect 11701 36799 11759 36805
rect 11882 36796 11888 36848
rect 11940 36836 11946 36848
rect 13446 36836 13452 36848
rect 11940 36808 12282 36836
rect 13407 36808 13452 36836
rect 11940 36796 11946 36808
rect 13446 36796 13452 36808
rect 13504 36796 13510 36848
rect 17681 36839 17739 36845
rect 17681 36836 17693 36839
rect 14476 36808 17693 36836
rect 8680 36740 9720 36768
rect 11164 36740 11652 36768
rect 6822 36660 6828 36712
rect 6880 36700 6886 36712
rect 8680 36709 8708 36740
rect 7193 36703 7251 36709
rect 7193 36700 7205 36703
rect 6880 36672 7205 36700
rect 6880 36660 6886 36672
rect 7193 36669 7205 36672
rect 7239 36700 7251 36703
rect 8665 36703 8723 36709
rect 7239 36672 8616 36700
rect 7239 36669 7251 36672
rect 7193 36663 7251 36669
rect 8588 36632 8616 36672
rect 8665 36669 8677 36703
rect 8711 36669 8723 36703
rect 8665 36663 8723 36669
rect 9125 36703 9183 36709
rect 9125 36669 9137 36703
rect 9171 36669 9183 36703
rect 9692 36700 9720 36740
rect 9858 36700 9864 36712
rect 9692 36672 9864 36700
rect 9125 36663 9183 36669
rect 9030 36632 9036 36644
rect 8588 36604 9036 36632
rect 9030 36592 9036 36604
rect 9088 36592 9094 36644
rect 8386 36564 8392 36576
rect 6748 36536 8392 36564
rect 8386 36524 8392 36536
rect 8444 36564 8450 36576
rect 8938 36564 8944 36576
rect 8444 36536 8944 36564
rect 8444 36524 8450 36536
rect 8938 36524 8944 36536
rect 8996 36524 9002 36576
rect 9140 36564 9168 36663
rect 9858 36660 9864 36672
rect 9916 36660 9922 36712
rect 10870 36700 10876 36712
rect 10831 36672 10876 36700
rect 10870 36660 10876 36672
rect 10928 36660 10934 36712
rect 11149 36703 11207 36709
rect 11149 36669 11161 36703
rect 11195 36700 11207 36703
rect 11514 36700 11520 36712
rect 11195 36672 11520 36700
rect 11195 36669 11207 36672
rect 11149 36663 11207 36669
rect 11514 36660 11520 36672
rect 11572 36660 11578 36712
rect 11624 36700 11652 36740
rect 13722 36728 13728 36780
rect 13780 36768 13786 36780
rect 14476 36777 14504 36808
rect 17681 36805 17693 36808
rect 17727 36805 17739 36839
rect 17681 36799 17739 36805
rect 17862 36796 17868 36848
rect 17920 36836 17926 36848
rect 22066 36836 22094 36876
rect 30650 36864 30656 36876
rect 30708 36864 30714 36916
rect 38194 36904 38200 36916
rect 38155 36876 38200 36904
rect 38194 36864 38200 36876
rect 38252 36864 38258 36916
rect 17920 36808 22094 36836
rect 17920 36796 17926 36808
rect 27614 36796 27620 36848
rect 27672 36836 27678 36848
rect 35526 36836 35532 36848
rect 27672 36808 35532 36836
rect 27672 36796 27678 36808
rect 35526 36796 35532 36808
rect 35584 36796 35590 36848
rect 14461 36771 14519 36777
rect 13780 36740 13825 36768
rect 13780 36728 13786 36740
rect 14461 36737 14473 36771
rect 14507 36737 14519 36771
rect 14461 36731 14519 36737
rect 14921 36771 14979 36777
rect 14921 36737 14933 36771
rect 14967 36737 14979 36771
rect 14921 36731 14979 36737
rect 14936 36700 14964 36731
rect 15010 36728 15016 36780
rect 15068 36768 15074 36780
rect 15746 36768 15752 36780
rect 15068 36740 15752 36768
rect 15068 36728 15074 36740
rect 15746 36728 15752 36740
rect 15804 36768 15810 36780
rect 15841 36771 15899 36777
rect 15841 36768 15853 36771
rect 15804 36740 15853 36768
rect 15804 36728 15810 36740
rect 15841 36737 15853 36740
rect 15887 36737 15899 36771
rect 15841 36731 15899 36737
rect 17037 36771 17095 36777
rect 17037 36737 17049 36771
rect 17083 36737 17095 36771
rect 17037 36731 17095 36737
rect 11624 36672 14320 36700
rect 12434 36632 12440 36644
rect 11072 36604 12440 36632
rect 11072 36564 11100 36604
rect 12434 36592 12440 36604
rect 12492 36592 12498 36644
rect 14292 36641 14320 36672
rect 14384 36672 14964 36700
rect 14277 36635 14335 36641
rect 14277 36601 14289 36635
rect 14323 36601 14335 36635
rect 14277 36595 14335 36601
rect 9140 36536 11100 36564
rect 11146 36524 11152 36576
rect 11204 36564 11210 36576
rect 14384 36564 14412 36672
rect 15286 36660 15292 36712
rect 15344 36700 15350 36712
rect 17052 36700 17080 36731
rect 17494 36728 17500 36780
rect 17552 36768 17558 36780
rect 17773 36771 17831 36777
rect 17773 36768 17785 36771
rect 17552 36740 17785 36768
rect 17552 36728 17558 36740
rect 17773 36737 17785 36740
rect 17819 36737 17831 36771
rect 17773 36731 17831 36737
rect 18046 36728 18052 36780
rect 18104 36768 18110 36780
rect 18877 36771 18935 36777
rect 18877 36768 18889 36771
rect 18104 36740 18889 36768
rect 18104 36728 18110 36740
rect 18877 36737 18889 36740
rect 18923 36768 18935 36771
rect 19521 36771 19579 36777
rect 19521 36768 19533 36771
rect 18923 36740 19533 36768
rect 18923 36737 18935 36740
rect 18877 36731 18935 36737
rect 19521 36737 19533 36740
rect 19567 36737 19579 36771
rect 19521 36731 19579 36737
rect 19978 36728 19984 36780
rect 20036 36768 20042 36780
rect 23385 36771 23443 36777
rect 23385 36768 23397 36771
rect 20036 36740 23397 36768
rect 20036 36728 20042 36740
rect 23385 36737 23397 36740
rect 23431 36737 23443 36771
rect 25409 36771 25467 36777
rect 25409 36768 25421 36771
rect 23385 36731 23443 36737
rect 23492 36740 25421 36768
rect 20714 36700 20720 36712
rect 15344 36672 20720 36700
rect 15344 36660 15350 36672
rect 20714 36660 20720 36672
rect 20772 36660 20778 36712
rect 20806 36660 20812 36712
rect 20864 36700 20870 36712
rect 23492 36700 23520 36740
rect 25409 36737 25421 36740
rect 25455 36768 25467 36771
rect 26053 36771 26111 36777
rect 26053 36768 26065 36771
rect 25455 36740 26065 36768
rect 25455 36737 25467 36740
rect 25409 36731 25467 36737
rect 26053 36737 26065 36740
rect 26099 36737 26111 36771
rect 26053 36731 26111 36737
rect 31662 36728 31668 36780
rect 31720 36768 31726 36780
rect 32493 36771 32551 36777
rect 32493 36768 32505 36771
rect 31720 36740 32505 36768
rect 31720 36728 31726 36740
rect 32493 36737 32505 36740
rect 32539 36768 32551 36771
rect 33137 36771 33195 36777
rect 33137 36768 33149 36771
rect 32539 36740 33149 36768
rect 32539 36737 32551 36740
rect 32493 36731 32551 36737
rect 33137 36737 33149 36740
rect 33183 36737 33195 36771
rect 34330 36768 34336 36780
rect 34291 36740 34336 36768
rect 33137 36731 33195 36737
rect 34330 36728 34336 36740
rect 34388 36768 34394 36780
rect 34977 36771 35035 36777
rect 34977 36768 34989 36771
rect 34388 36740 34989 36768
rect 34388 36728 34394 36740
rect 34977 36737 34989 36740
rect 35023 36737 35035 36771
rect 38013 36771 38071 36777
rect 38013 36768 38025 36771
rect 34977 36731 35035 36737
rect 35866 36740 38025 36768
rect 31846 36700 31852 36712
rect 20864 36672 23520 36700
rect 24872 36672 31852 36700
rect 20864 36660 20870 36672
rect 21085 36635 21143 36641
rect 21085 36632 21097 36635
rect 19996 36604 21097 36632
rect 19996 36576 20024 36604
rect 21085 36601 21097 36604
rect 21131 36632 21143 36635
rect 22005 36635 22063 36641
rect 22005 36632 22017 36635
rect 21131 36604 22017 36632
rect 21131 36601 21143 36604
rect 21085 36595 21143 36601
rect 22005 36601 22017 36604
rect 22051 36632 22063 36635
rect 22186 36632 22192 36644
rect 22051 36604 22192 36632
rect 22051 36601 22063 36604
rect 22005 36595 22063 36601
rect 22186 36592 22192 36604
rect 22244 36632 22250 36644
rect 22557 36635 22615 36641
rect 22557 36632 22569 36635
rect 22244 36604 22569 36632
rect 22244 36592 22250 36604
rect 22557 36601 22569 36604
rect 22603 36601 22615 36635
rect 22557 36595 22615 36601
rect 23290 36592 23296 36644
rect 23348 36632 23354 36644
rect 24029 36635 24087 36641
rect 24029 36632 24041 36635
rect 23348 36604 24041 36632
rect 23348 36592 23354 36604
rect 24029 36601 24041 36604
rect 24075 36632 24087 36635
rect 24581 36635 24639 36641
rect 24581 36632 24593 36635
rect 24075 36604 24593 36632
rect 24075 36601 24087 36604
rect 24029 36595 24087 36601
rect 24581 36601 24593 36604
rect 24627 36601 24639 36635
rect 24581 36595 24639 36601
rect 11204 36536 14412 36564
rect 11204 36524 11210 36536
rect 15010 36524 15016 36576
rect 15068 36564 15074 36576
rect 16850 36564 16856 36576
rect 15068 36536 15113 36564
rect 16811 36536 16856 36564
rect 15068 36524 15074 36536
rect 16850 36524 16856 36536
rect 16908 36524 16914 36576
rect 18782 36564 18788 36576
rect 18743 36536 18788 36564
rect 18782 36524 18788 36536
rect 18840 36524 18846 36576
rect 19334 36524 19340 36576
rect 19392 36564 19398 36576
rect 19429 36567 19487 36573
rect 19429 36564 19441 36567
rect 19392 36536 19441 36564
rect 19392 36524 19398 36536
rect 19429 36533 19441 36536
rect 19475 36533 19487 36567
rect 19978 36564 19984 36576
rect 19939 36536 19984 36564
rect 19429 36527 19487 36533
rect 19978 36524 19984 36536
rect 20036 36524 20042 36576
rect 20530 36564 20536 36576
rect 20491 36536 20536 36564
rect 20530 36524 20536 36536
rect 20588 36524 20594 36576
rect 23569 36567 23627 36573
rect 23569 36533 23581 36567
rect 23615 36564 23627 36567
rect 24872 36564 24900 36672
rect 31846 36660 31852 36672
rect 31904 36660 31910 36712
rect 32585 36703 32643 36709
rect 32585 36669 32597 36703
rect 32631 36700 32643 36703
rect 35866 36700 35894 36740
rect 38013 36737 38025 36740
rect 38059 36737 38071 36771
rect 38013 36731 38071 36737
rect 32631 36672 35894 36700
rect 32631 36669 32643 36672
rect 32585 36663 32643 36669
rect 25593 36635 25651 36641
rect 25593 36601 25605 36635
rect 25639 36632 25651 36635
rect 28902 36632 28908 36644
rect 25639 36604 28908 36632
rect 25639 36601 25651 36604
rect 25593 36595 25651 36601
rect 28902 36592 28908 36604
rect 28960 36592 28966 36644
rect 34422 36564 34428 36576
rect 23615 36536 24900 36564
rect 34383 36536 34428 36564
rect 23615 36533 23627 36536
rect 23569 36527 23627 36533
rect 34422 36524 34428 36536
rect 34480 36524 34486 36576
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 4420 36363 4478 36369
rect 4420 36329 4432 36363
rect 4466 36360 4478 36363
rect 4614 36360 4620 36372
rect 4466 36332 4620 36360
rect 4466 36329 4478 36332
rect 4420 36323 4478 36329
rect 4614 36320 4620 36332
rect 4672 36360 4678 36372
rect 11146 36360 11152 36372
rect 4672 36332 11152 36360
rect 4672 36320 4678 36332
rect 11146 36320 11152 36332
rect 11204 36320 11210 36372
rect 12158 36360 12164 36372
rect 11348 36332 12164 36360
rect 10318 36252 10324 36304
rect 10376 36292 10382 36304
rect 11348 36292 11376 36332
rect 12158 36320 12164 36332
rect 12216 36320 12222 36372
rect 12250 36320 12256 36372
rect 12308 36360 12314 36372
rect 13173 36363 13231 36369
rect 13173 36360 13185 36363
rect 12308 36332 13185 36360
rect 12308 36320 12314 36332
rect 13173 36329 13185 36332
rect 13219 36329 13231 36363
rect 13173 36323 13231 36329
rect 13262 36320 13268 36372
rect 13320 36360 13326 36372
rect 20533 36363 20591 36369
rect 20533 36360 20545 36363
rect 13320 36332 20545 36360
rect 13320 36320 13326 36332
rect 20533 36329 20545 36332
rect 20579 36329 20591 36363
rect 22186 36360 22192 36372
rect 22147 36332 22192 36360
rect 20533 36323 20591 36329
rect 22186 36320 22192 36332
rect 22244 36360 22250 36372
rect 22741 36363 22799 36369
rect 22741 36360 22753 36363
rect 22244 36332 22753 36360
rect 22244 36320 22250 36332
rect 22741 36329 22753 36332
rect 22787 36360 22799 36363
rect 23290 36360 23296 36372
rect 22787 36332 23296 36360
rect 22787 36329 22799 36332
rect 22741 36323 22799 36329
rect 23290 36320 23296 36332
rect 23348 36360 23354 36372
rect 23845 36363 23903 36369
rect 23845 36360 23857 36363
rect 23348 36332 23857 36360
rect 23348 36320 23354 36332
rect 23845 36329 23857 36332
rect 23891 36360 23903 36363
rect 25133 36363 25191 36369
rect 25133 36360 25145 36363
rect 23891 36332 25145 36360
rect 23891 36329 23903 36332
rect 23845 36323 23903 36329
rect 25133 36329 25145 36332
rect 25179 36329 25191 36363
rect 25133 36323 25191 36329
rect 38197 36363 38255 36369
rect 38197 36329 38209 36363
rect 38243 36360 38255 36363
rect 38654 36360 38660 36372
rect 38243 36332 38660 36360
rect 38243 36329 38255 36332
rect 38197 36323 38255 36329
rect 38654 36320 38660 36332
rect 38712 36320 38718 36372
rect 15746 36292 15752 36304
rect 10376 36264 11376 36292
rect 12544 36264 15752 36292
rect 10376 36252 10382 36264
rect 1670 36224 1676 36236
rect 1583 36196 1676 36224
rect 1670 36184 1676 36196
rect 1728 36224 1734 36236
rect 3878 36224 3884 36236
rect 1728 36196 3884 36224
rect 1728 36184 1734 36196
rect 3878 36184 3884 36196
rect 3936 36224 3942 36236
rect 4157 36227 4215 36233
rect 4157 36224 4169 36227
rect 3936 36196 4169 36224
rect 3936 36184 3942 36196
rect 4157 36193 4169 36196
rect 4203 36193 4215 36227
rect 4157 36187 4215 36193
rect 4798 36184 4804 36236
rect 4856 36224 4862 36236
rect 6365 36227 6423 36233
rect 6365 36224 6377 36227
rect 4856 36196 6377 36224
rect 4856 36184 4862 36196
rect 6365 36193 6377 36196
rect 6411 36193 6423 36227
rect 8110 36224 8116 36236
rect 8071 36196 8116 36224
rect 6365 36187 6423 36193
rect 8110 36184 8116 36196
rect 8168 36184 8174 36236
rect 8570 36184 8576 36236
rect 8628 36224 8634 36236
rect 12250 36224 12256 36236
rect 8628 36196 12256 36224
rect 8628 36184 8634 36196
rect 12250 36184 12256 36196
rect 12308 36184 12314 36236
rect 12342 36184 12348 36236
rect 12400 36224 12406 36236
rect 12544 36224 12572 36264
rect 15746 36252 15752 36264
rect 15804 36252 15810 36304
rect 15930 36252 15936 36304
rect 15988 36292 15994 36304
rect 19150 36292 19156 36304
rect 15988 36264 19156 36292
rect 15988 36252 15994 36264
rect 19150 36252 19156 36264
rect 19208 36252 19214 36304
rect 19242 36252 19248 36304
rect 19300 36292 19306 36304
rect 24762 36292 24768 36304
rect 19300 36264 24768 36292
rect 19300 36252 19306 36264
rect 24762 36252 24768 36264
rect 24820 36252 24826 36304
rect 12400 36196 12572 36224
rect 12621 36227 12679 36233
rect 12400 36184 12406 36196
rect 12621 36193 12633 36227
rect 12667 36224 12679 36227
rect 13722 36224 13728 36236
rect 12667 36196 13728 36224
rect 12667 36193 12679 36196
rect 12621 36187 12679 36193
rect 13722 36184 13728 36196
rect 13780 36224 13786 36236
rect 19429 36227 19487 36233
rect 19429 36224 19441 36227
rect 13780 36196 19441 36224
rect 13780 36184 13786 36196
rect 19429 36193 19441 36196
rect 19475 36224 19487 36227
rect 19978 36224 19984 36236
rect 19475 36196 19984 36224
rect 19475 36193 19487 36196
rect 19429 36187 19487 36193
rect 19978 36184 19984 36196
rect 20036 36224 20042 36236
rect 21085 36227 21143 36233
rect 21085 36224 21097 36227
rect 20036 36196 21097 36224
rect 20036 36184 20042 36196
rect 21085 36193 21097 36196
rect 21131 36193 21143 36227
rect 34330 36224 34336 36236
rect 21085 36187 21143 36193
rect 28966 36196 34336 36224
rect 8386 36116 8392 36168
rect 8444 36156 8450 36168
rect 8444 36128 8489 36156
rect 8444 36116 8450 36128
rect 8846 36116 8852 36168
rect 8904 36156 8910 36168
rect 9861 36159 9919 36165
rect 9861 36156 9873 36159
rect 8904 36128 9873 36156
rect 8904 36116 8910 36128
rect 9861 36125 9873 36128
rect 9907 36125 9919 36159
rect 9861 36119 9919 36125
rect 10137 36159 10195 36165
rect 10137 36125 10149 36159
rect 10183 36156 10195 36159
rect 10318 36156 10324 36168
rect 10183 36128 10324 36156
rect 10183 36125 10195 36128
rect 10137 36119 10195 36125
rect 10318 36116 10324 36128
rect 10376 36116 10382 36168
rect 13357 36159 13415 36165
rect 13357 36125 13369 36159
rect 13403 36125 13415 36159
rect 14642 36156 14648 36168
rect 14603 36128 14648 36156
rect 13357 36119 13415 36125
rect 1949 36091 2007 36097
rect 1949 36088 1961 36091
rect 1780 36060 1961 36088
rect 1780 36032 1808 36060
rect 1949 36057 1961 36060
rect 1995 36057 2007 36091
rect 1949 36051 2007 36057
rect 2498 36048 2504 36100
rect 2556 36048 2562 36100
rect 3510 36048 3516 36100
rect 3568 36088 3574 36100
rect 8754 36088 8760 36100
rect 3568 36060 4922 36088
rect 7682 36060 8760 36088
rect 3568 36048 3574 36060
rect 8754 36048 8760 36060
rect 8812 36048 8818 36100
rect 9674 36048 9680 36100
rect 9732 36088 9738 36100
rect 10597 36091 10655 36097
rect 10597 36088 10609 36091
rect 9732 36060 10609 36088
rect 9732 36048 9738 36060
rect 10597 36057 10609 36060
rect 10643 36057 10655 36091
rect 10597 36051 10655 36057
rect 11330 36048 11336 36100
rect 11388 36048 11394 36100
rect 12342 36088 12348 36100
rect 12176 36060 12348 36088
rect 1762 35980 1768 36032
rect 1820 35980 1826 36032
rect 3421 36023 3479 36029
rect 3421 35989 3433 36023
rect 3467 36020 3479 36023
rect 4706 36020 4712 36032
rect 3467 35992 4712 36020
rect 3467 35989 3479 35992
rect 3421 35983 3479 35989
rect 4706 35980 4712 35992
rect 4764 35980 4770 36032
rect 5905 36023 5963 36029
rect 5905 35989 5917 36023
rect 5951 36020 5963 36023
rect 12176 36020 12204 36060
rect 12342 36048 12348 36060
rect 12400 36048 12406 36100
rect 12434 36048 12440 36100
rect 12492 36088 12498 36100
rect 13262 36088 13268 36100
rect 12492 36060 13268 36088
rect 12492 36048 12498 36060
rect 13262 36048 13268 36060
rect 13320 36048 13326 36100
rect 13372 36088 13400 36119
rect 14642 36116 14648 36128
rect 14700 36116 14706 36168
rect 15286 36156 15292 36168
rect 15247 36128 15292 36156
rect 15286 36116 15292 36128
rect 15344 36116 15350 36168
rect 15746 36156 15752 36168
rect 15707 36128 15752 36156
rect 15746 36116 15752 36128
rect 15804 36116 15810 36168
rect 16022 36116 16028 36168
rect 16080 36156 16086 36168
rect 17957 36159 18015 36165
rect 17957 36156 17969 36159
rect 16080 36128 17969 36156
rect 16080 36116 16086 36128
rect 17957 36125 17969 36128
rect 18003 36125 18015 36159
rect 17957 36119 18015 36125
rect 16850 36088 16856 36100
rect 13372 36060 16856 36088
rect 16850 36048 16856 36060
rect 16908 36048 16914 36100
rect 17972 36088 18000 36119
rect 18874 36116 18880 36168
rect 18932 36156 18938 36168
rect 28966 36156 28994 36196
rect 34330 36184 34336 36196
rect 34388 36184 34394 36236
rect 18932 36128 28994 36156
rect 18932 36116 18938 36128
rect 34422 36116 34428 36168
rect 34480 36156 34486 36168
rect 38013 36159 38071 36165
rect 38013 36156 38025 36159
rect 34480 36128 38025 36156
rect 34480 36116 34486 36128
rect 38013 36125 38025 36128
rect 38059 36125 38071 36159
rect 38013 36119 38071 36125
rect 17972 36060 19196 36088
rect 5951 35992 12204 36020
rect 5951 35989 5963 35992
rect 5905 35983 5963 35989
rect 12250 35980 12256 36032
rect 12308 36020 12314 36032
rect 14458 36020 14464 36032
rect 12308 35992 14464 36020
rect 12308 35980 12314 35992
rect 14458 35980 14464 35992
rect 14516 35980 14522 36032
rect 14553 36023 14611 36029
rect 14553 35989 14565 36023
rect 14599 36020 14611 36023
rect 14734 36020 14740 36032
rect 14599 35992 14740 36020
rect 14599 35989 14611 35992
rect 14553 35983 14611 35989
rect 14734 35980 14740 35992
rect 14792 35980 14798 36032
rect 14918 35980 14924 36032
rect 14976 36020 14982 36032
rect 15197 36023 15255 36029
rect 15197 36020 15209 36023
rect 14976 35992 15209 36020
rect 14976 35980 14982 35992
rect 15197 35989 15209 35992
rect 15243 35989 15255 36023
rect 15197 35983 15255 35989
rect 15378 35980 15384 36032
rect 15436 36020 15442 36032
rect 15841 36023 15899 36029
rect 15841 36020 15853 36023
rect 15436 35992 15853 36020
rect 15436 35980 15442 35992
rect 15841 35989 15853 35992
rect 15887 35989 15899 36023
rect 16390 36020 16396 36032
rect 16351 35992 16396 36020
rect 15841 35983 15899 35989
rect 16390 35980 16396 35992
rect 16448 35980 16454 36032
rect 17497 36023 17555 36029
rect 17497 35989 17509 36023
rect 17543 36020 17555 36023
rect 17770 36020 17776 36032
rect 17543 35992 17776 36020
rect 17543 35989 17555 35992
rect 17497 35983 17555 35989
rect 17770 35980 17776 35992
rect 17828 35980 17834 36032
rect 18506 36020 18512 36032
rect 18467 35992 18512 36020
rect 18506 35980 18512 35992
rect 18564 36020 18570 36032
rect 19058 36020 19064 36032
rect 18564 35992 19064 36020
rect 18564 35980 18570 35992
rect 19058 35980 19064 35992
rect 19116 35980 19122 36032
rect 19168 36020 19196 36060
rect 19334 36048 19340 36100
rect 19392 36088 19398 36100
rect 23106 36088 23112 36100
rect 19392 36060 23112 36088
rect 19392 36048 19398 36060
rect 23106 36048 23112 36060
rect 23164 36048 23170 36100
rect 20806 36020 20812 36032
rect 19168 35992 20812 36020
rect 20806 35980 20812 35992
rect 20864 35980 20870 36032
rect 21634 36020 21640 36032
rect 21595 35992 21640 36020
rect 21634 35980 21640 35992
rect 21692 35980 21698 36032
rect 24578 36020 24584 36032
rect 24539 35992 24584 36020
rect 24578 35980 24584 35992
rect 24636 35980 24642 36032
rect 25682 36020 25688 36032
rect 25643 35992 25688 36020
rect 25682 35980 25688 35992
rect 25740 35980 25746 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 3510 35776 3516 35828
rect 3568 35816 3574 35828
rect 8018 35816 8024 35828
rect 3568 35788 8024 35816
rect 3568 35776 3574 35788
rect 8018 35776 8024 35788
rect 8076 35776 8082 35828
rect 8478 35776 8484 35828
rect 8536 35816 8542 35828
rect 10594 35816 10600 35828
rect 8536 35788 10600 35816
rect 8536 35776 8542 35788
rect 10594 35776 10600 35788
rect 10652 35776 10658 35828
rect 10686 35776 10692 35828
rect 10744 35816 10750 35828
rect 10744 35788 11284 35816
rect 10744 35776 10750 35788
rect 1673 35751 1731 35757
rect 1673 35717 1685 35751
rect 1719 35748 1731 35751
rect 2866 35748 2872 35760
rect 1719 35720 2872 35748
rect 1719 35717 1731 35720
rect 1673 35711 1731 35717
rect 2866 35708 2872 35720
rect 2924 35748 2930 35760
rect 3786 35748 3792 35760
rect 2924 35720 3792 35748
rect 2924 35708 2930 35720
rect 3786 35708 3792 35720
rect 3844 35708 3850 35760
rect 5077 35751 5135 35757
rect 5077 35717 5089 35751
rect 5123 35748 5135 35751
rect 5442 35748 5448 35760
rect 5123 35720 5448 35748
rect 5123 35717 5135 35720
rect 5077 35711 5135 35717
rect 5442 35708 5448 35720
rect 5500 35708 5506 35760
rect 8202 35708 8208 35760
rect 8260 35708 8266 35760
rect 8662 35708 8668 35760
rect 8720 35748 8726 35760
rect 8720 35720 8765 35748
rect 8720 35708 8726 35720
rect 10778 35708 10784 35760
rect 10836 35748 10842 35760
rect 11256 35748 11284 35788
rect 11330 35776 11336 35828
rect 11388 35816 11394 35828
rect 11514 35816 11520 35828
rect 11388 35788 11520 35816
rect 11388 35776 11394 35788
rect 11514 35776 11520 35788
rect 11572 35816 11578 35828
rect 11572 35788 13492 35816
rect 11572 35776 11578 35788
rect 13170 35748 13176 35760
rect 10836 35720 11192 35748
rect 11256 35720 12006 35748
rect 13131 35720 13176 35748
rect 10836 35708 10842 35720
rect 1946 35640 1952 35692
rect 2004 35680 2010 35692
rect 2774 35680 2780 35692
rect 2004 35652 2780 35680
rect 2004 35640 2010 35652
rect 2774 35640 2780 35652
rect 2832 35640 2838 35692
rect 3970 35640 3976 35692
rect 4028 35640 4034 35692
rect 5350 35640 5356 35692
rect 5408 35680 5414 35692
rect 5997 35683 6055 35689
rect 5408 35652 5453 35680
rect 5408 35640 5414 35652
rect 5997 35649 6009 35683
rect 6043 35680 6055 35683
rect 6638 35680 6644 35692
rect 6043 35652 6644 35680
rect 6043 35649 6055 35652
rect 5997 35643 6055 35649
rect 6638 35640 6644 35652
rect 6696 35640 6702 35692
rect 8938 35640 8944 35692
rect 8996 35680 9002 35692
rect 8996 35652 9041 35680
rect 8996 35640 9002 35652
rect 9766 35640 9772 35692
rect 9824 35640 9830 35692
rect 11164 35680 11192 35720
rect 13170 35708 13176 35720
rect 13228 35708 13234 35760
rect 13464 35689 13492 35788
rect 14458 35776 14464 35828
rect 14516 35816 14522 35828
rect 17681 35819 17739 35825
rect 17681 35816 17693 35819
rect 14516 35788 17693 35816
rect 14516 35776 14522 35788
rect 17681 35785 17693 35788
rect 17727 35785 17739 35819
rect 17681 35779 17739 35785
rect 17954 35776 17960 35828
rect 18012 35816 18018 35828
rect 18012 35788 19932 35816
rect 18012 35776 18018 35788
rect 14001 35751 14059 35757
rect 14001 35717 14013 35751
rect 14047 35748 14059 35751
rect 14047 35720 15148 35748
rect 14047 35717 14059 35720
rect 14001 35711 14059 35717
rect 13449 35683 13507 35689
rect 11164 35652 11652 35680
rect 2866 35612 2872 35624
rect 2827 35584 2872 35612
rect 2866 35572 2872 35584
rect 2924 35572 2930 35624
rect 3145 35615 3203 35621
rect 3145 35581 3157 35615
rect 3191 35612 3203 35615
rect 5074 35612 5080 35624
rect 3191 35584 5080 35612
rect 3191 35581 3203 35584
rect 3145 35575 3203 35581
rect 5074 35572 5080 35584
rect 5132 35612 5138 35624
rect 7193 35615 7251 35621
rect 5132 35584 5304 35612
rect 5132 35572 5138 35584
rect 1854 35544 1860 35556
rect 1815 35516 1860 35544
rect 1854 35504 1860 35516
rect 1912 35504 1918 35556
rect 1946 35504 1952 35556
rect 2004 35544 2010 35556
rect 5276 35544 5304 35584
rect 7193 35581 7205 35615
rect 7239 35612 7251 35615
rect 9306 35612 9312 35624
rect 7239 35584 9312 35612
rect 7239 35581 7251 35584
rect 7193 35575 7251 35581
rect 9306 35572 9312 35584
rect 9364 35572 9370 35624
rect 9398 35572 9404 35624
rect 9456 35612 9462 35624
rect 10502 35612 10508 35624
rect 9456 35584 10508 35612
rect 9456 35572 9462 35584
rect 10502 35572 10508 35584
rect 10560 35572 10566 35624
rect 10873 35615 10931 35621
rect 10873 35581 10885 35615
rect 10919 35612 10931 35615
rect 11149 35615 11207 35621
rect 10919 35584 11100 35612
rect 10919 35581 10931 35584
rect 10873 35575 10931 35581
rect 7466 35544 7472 35556
rect 2004 35516 4108 35544
rect 5276 35516 7472 35544
rect 2004 35504 2010 35516
rect 3602 35476 3608 35488
rect 3563 35448 3608 35476
rect 3602 35436 3608 35448
rect 3660 35436 3666 35488
rect 4080 35476 4108 35516
rect 7466 35504 7472 35516
rect 7524 35504 7530 35556
rect 9858 35544 9864 35556
rect 9324 35516 9864 35544
rect 5626 35476 5632 35488
rect 4080 35448 5632 35476
rect 5626 35436 5632 35448
rect 5684 35436 5690 35488
rect 5902 35476 5908 35488
rect 5863 35448 5908 35476
rect 5902 35436 5908 35448
rect 5960 35436 5966 35488
rect 6641 35479 6699 35485
rect 6641 35445 6653 35479
rect 6687 35476 6699 35479
rect 7190 35476 7196 35488
rect 6687 35448 7196 35476
rect 6687 35445 6699 35448
rect 6641 35439 6699 35445
rect 7190 35436 7196 35448
rect 7248 35436 7254 35488
rect 8202 35436 8208 35488
rect 8260 35476 8266 35488
rect 9324 35476 9352 35516
rect 9858 35504 9864 35516
rect 9916 35504 9922 35556
rect 11072 35544 11100 35584
rect 11149 35581 11161 35615
rect 11195 35612 11207 35615
rect 11330 35612 11336 35624
rect 11195 35584 11336 35612
rect 11195 35581 11207 35584
rect 11149 35575 11207 35581
rect 11330 35572 11336 35584
rect 11388 35572 11394 35624
rect 11624 35612 11652 35652
rect 13449 35649 13461 35683
rect 13495 35680 13507 35683
rect 13722 35680 13728 35692
rect 13495 35652 13728 35680
rect 13495 35649 13507 35652
rect 13449 35643 13507 35649
rect 13722 35640 13728 35652
rect 13780 35640 13786 35692
rect 14182 35640 14188 35692
rect 14240 35680 14246 35692
rect 14461 35683 14519 35689
rect 14461 35680 14473 35683
rect 14240 35652 14473 35680
rect 14240 35640 14246 35652
rect 14461 35649 14473 35652
rect 14507 35649 14519 35683
rect 15120 35680 15148 35720
rect 15194 35708 15200 35760
rect 15252 35748 15258 35760
rect 15252 35720 16896 35748
rect 15252 35708 15258 35720
rect 15286 35680 15292 35692
rect 15120 35652 15292 35680
rect 14461 35643 14519 35649
rect 15286 35640 15292 35652
rect 15344 35640 15350 35692
rect 15470 35680 15476 35692
rect 15431 35652 15476 35680
rect 15470 35640 15476 35652
rect 15528 35640 15534 35692
rect 16022 35640 16028 35692
rect 16080 35680 16086 35692
rect 16868 35689 16896 35720
rect 16942 35708 16948 35760
rect 17000 35748 17006 35760
rect 18969 35751 19027 35757
rect 18969 35748 18981 35751
rect 17000 35720 18981 35748
rect 17000 35708 17006 35720
rect 18969 35717 18981 35720
rect 19015 35717 19027 35751
rect 19904 35748 19932 35788
rect 19978 35776 19984 35828
rect 20036 35816 20042 35828
rect 20073 35819 20131 35825
rect 20073 35816 20085 35819
rect 20036 35788 20085 35816
rect 20036 35776 20042 35788
rect 20073 35785 20085 35788
rect 20119 35816 20131 35819
rect 20625 35819 20683 35825
rect 20625 35816 20637 35819
rect 20119 35788 20637 35816
rect 20119 35785 20131 35788
rect 20073 35779 20131 35785
rect 20625 35785 20637 35788
rect 20671 35816 20683 35819
rect 21082 35816 21088 35828
rect 20671 35788 21088 35816
rect 20671 35785 20683 35788
rect 20625 35779 20683 35785
rect 21082 35776 21088 35788
rect 21140 35816 21146 35828
rect 21177 35819 21235 35825
rect 21177 35816 21189 35819
rect 21140 35788 21189 35816
rect 21140 35776 21146 35788
rect 21177 35785 21189 35788
rect 21223 35816 21235 35819
rect 22005 35819 22063 35825
rect 22005 35816 22017 35819
rect 21223 35788 22017 35816
rect 21223 35785 21235 35788
rect 21177 35779 21235 35785
rect 22005 35785 22017 35788
rect 22051 35816 22063 35819
rect 23109 35819 23167 35825
rect 23109 35816 23121 35819
rect 22051 35788 23121 35816
rect 22051 35785 22063 35788
rect 22005 35779 22063 35785
rect 23109 35785 23121 35788
rect 23155 35816 23167 35819
rect 23661 35819 23719 35825
rect 23661 35816 23673 35819
rect 23155 35788 23673 35816
rect 23155 35785 23167 35788
rect 23109 35779 23167 35785
rect 23661 35785 23673 35788
rect 23707 35816 23719 35819
rect 24765 35819 24823 35825
rect 24765 35816 24777 35819
rect 23707 35788 24777 35816
rect 23707 35785 23719 35788
rect 23661 35779 23719 35785
rect 24765 35785 24777 35788
rect 24811 35785 24823 35819
rect 24765 35779 24823 35785
rect 27525 35819 27583 35825
rect 27525 35785 27537 35819
rect 27571 35816 27583 35819
rect 27614 35816 27620 35828
rect 27571 35788 27620 35816
rect 27571 35785 27583 35788
rect 27525 35779 27583 35785
rect 27614 35776 27620 35788
rect 27672 35776 27678 35828
rect 21634 35748 21640 35760
rect 19904 35720 21640 35748
rect 18969 35711 19027 35717
rect 21634 35708 21640 35720
rect 21692 35708 21698 35760
rect 22066 35720 26234 35748
rect 16301 35683 16359 35689
rect 16301 35680 16313 35683
rect 16080 35652 16313 35680
rect 16080 35640 16086 35652
rect 16301 35649 16313 35652
rect 16347 35649 16359 35683
rect 16301 35643 16359 35649
rect 16853 35683 16911 35689
rect 16853 35649 16865 35683
rect 16899 35649 16911 35683
rect 17770 35680 17776 35692
rect 17731 35652 17776 35680
rect 16853 35643 16911 35649
rect 17770 35640 17776 35652
rect 17828 35640 17834 35692
rect 18414 35640 18420 35692
rect 18472 35680 18478 35692
rect 22066 35680 22094 35720
rect 18472 35652 22094 35680
rect 26206 35680 26234 35720
rect 27433 35683 27491 35689
rect 27433 35680 27445 35683
rect 26206 35652 27445 35680
rect 18472 35640 18478 35652
rect 27433 35649 27445 35652
rect 27479 35649 27491 35683
rect 27433 35643 27491 35649
rect 37458 35640 37464 35692
rect 37516 35680 37522 35692
rect 38013 35683 38071 35689
rect 38013 35680 38025 35683
rect 37516 35652 38025 35680
rect 37516 35640 37522 35652
rect 38013 35649 38025 35652
rect 38059 35649 38071 35683
rect 38013 35643 38071 35649
rect 12710 35612 12716 35624
rect 11624 35584 12716 35612
rect 12710 35572 12716 35584
rect 12768 35572 12774 35624
rect 12802 35572 12808 35624
rect 12860 35612 12866 35624
rect 15654 35612 15660 35624
rect 12860 35584 15660 35612
rect 12860 35572 12866 35584
rect 15654 35572 15660 35584
rect 15712 35572 15718 35624
rect 16114 35572 16120 35624
rect 16172 35612 16178 35624
rect 19518 35612 19524 35624
rect 16172 35584 19524 35612
rect 16172 35572 16178 35584
rect 19518 35572 19524 35584
rect 19576 35572 19582 35624
rect 25314 35612 25320 35624
rect 25275 35584 25320 35612
rect 25314 35572 25320 35584
rect 25372 35572 25378 35624
rect 11701 35547 11759 35553
rect 11701 35544 11713 35547
rect 11072 35516 11713 35544
rect 11701 35513 11713 35516
rect 11747 35513 11759 35547
rect 11701 35507 11759 35513
rect 8260 35448 9352 35476
rect 9401 35479 9459 35485
rect 8260 35436 8266 35448
rect 9401 35445 9413 35479
rect 9447 35476 9459 35479
rect 10870 35476 10876 35488
rect 9447 35448 10876 35476
rect 9447 35445 9459 35448
rect 9401 35439 9459 35445
rect 10870 35436 10876 35448
rect 10928 35476 10934 35488
rect 11606 35476 11612 35488
rect 10928 35448 11612 35476
rect 10928 35436 10934 35448
rect 11606 35436 11612 35448
rect 11664 35436 11670 35488
rect 11716 35476 11744 35507
rect 13998 35504 14004 35556
rect 14056 35544 14062 35556
rect 24213 35547 24271 35553
rect 24213 35544 24225 35547
rect 14056 35516 24225 35544
rect 14056 35504 14062 35516
rect 24213 35513 24225 35516
rect 24259 35513 24271 35547
rect 24213 35507 24271 35513
rect 12802 35476 12808 35488
rect 11716 35448 12808 35476
rect 12802 35436 12808 35448
rect 12860 35436 12866 35488
rect 14553 35479 14611 35485
rect 14553 35445 14565 35479
rect 14599 35476 14611 35479
rect 15470 35476 15476 35488
rect 14599 35448 15476 35476
rect 14599 35445 14611 35448
rect 14553 35439 14611 35445
rect 15470 35436 15476 35448
rect 15528 35436 15534 35488
rect 15657 35479 15715 35485
rect 15657 35445 15669 35479
rect 15703 35476 15715 35479
rect 16114 35476 16120 35488
rect 15703 35448 16120 35476
rect 15703 35445 15715 35448
rect 15657 35439 15715 35445
rect 16114 35436 16120 35448
rect 16172 35436 16178 35488
rect 16209 35479 16267 35485
rect 16209 35445 16221 35479
rect 16255 35476 16267 35479
rect 16482 35476 16488 35488
rect 16255 35448 16488 35476
rect 16255 35445 16267 35448
rect 16209 35439 16267 35445
rect 16482 35436 16488 35448
rect 16540 35436 16546 35488
rect 16942 35476 16948 35488
rect 16903 35448 16948 35476
rect 16942 35436 16948 35448
rect 17000 35436 17006 35488
rect 17770 35436 17776 35488
rect 17828 35476 17834 35488
rect 18509 35479 18567 35485
rect 18509 35476 18521 35479
rect 17828 35448 18521 35476
rect 17828 35436 17834 35448
rect 18509 35445 18521 35448
rect 18555 35476 18567 35479
rect 19242 35476 19248 35488
rect 18555 35448 19248 35476
rect 18555 35445 18567 35448
rect 18509 35439 18567 35445
rect 19242 35436 19248 35448
rect 19300 35436 19306 35488
rect 19518 35476 19524 35488
rect 19479 35448 19524 35476
rect 19518 35436 19524 35448
rect 19576 35436 19582 35488
rect 20162 35436 20168 35488
rect 20220 35476 20226 35488
rect 22557 35479 22615 35485
rect 22557 35476 22569 35479
rect 20220 35448 22569 35476
rect 20220 35436 20226 35448
rect 22557 35445 22569 35448
rect 22603 35445 22615 35479
rect 37458 35476 37464 35488
rect 37419 35448 37464 35476
rect 22557 35439 22615 35445
rect 37458 35436 37464 35448
rect 37516 35436 37522 35488
rect 38194 35476 38200 35488
rect 38155 35448 38200 35476
rect 38194 35436 38200 35448
rect 38252 35436 38258 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 3421 35275 3479 35281
rect 3421 35241 3433 35275
rect 3467 35272 3479 35275
rect 3510 35272 3516 35284
rect 3467 35244 3516 35272
rect 3467 35241 3479 35244
rect 3421 35235 3479 35241
rect 3510 35232 3516 35244
rect 3568 35232 3574 35284
rect 10686 35272 10692 35284
rect 4448 35244 10692 35272
rect 1670 35136 1676 35148
rect 1631 35108 1676 35136
rect 1670 35096 1676 35108
rect 1728 35096 1734 35148
rect 4448 35068 4476 35244
rect 10686 35232 10692 35244
rect 10744 35232 10750 35284
rect 12250 35272 12256 35284
rect 10796 35244 12256 35272
rect 7650 35164 7656 35216
rect 7708 35204 7714 35216
rect 9355 35207 9413 35213
rect 9355 35204 9367 35207
rect 7708 35176 9367 35204
rect 7708 35164 7714 35176
rect 9355 35173 9367 35176
rect 9401 35173 9413 35207
rect 9355 35167 9413 35173
rect 5445 35139 5503 35145
rect 5445 35105 5457 35139
rect 5491 35136 5503 35139
rect 10796 35136 10824 35244
rect 12250 35232 12256 35244
rect 12308 35232 12314 35284
rect 15102 35272 15108 35284
rect 13096 35244 15108 35272
rect 13096 35204 13124 35244
rect 15102 35232 15108 35244
rect 15160 35232 15166 35284
rect 15194 35232 15200 35284
rect 15252 35272 15258 35284
rect 18046 35272 18052 35284
rect 15252 35244 15516 35272
rect 18007 35244 18052 35272
rect 15252 35232 15258 35244
rect 12176 35176 13124 35204
rect 5491 35108 10824 35136
rect 10873 35139 10931 35145
rect 5491 35105 5503 35108
rect 5445 35099 5503 35105
rect 10873 35105 10885 35139
rect 10919 35136 10931 35139
rect 11514 35136 11520 35148
rect 10919 35108 11520 35136
rect 10919 35105 10931 35108
rect 10873 35099 10931 35105
rect 11514 35096 11520 35108
rect 11572 35096 11578 35148
rect 11606 35096 11612 35148
rect 11664 35136 11670 35148
rect 12176 35136 12204 35176
rect 13170 35164 13176 35216
rect 13228 35204 13234 35216
rect 15488 35204 15516 35244
rect 18046 35232 18052 35244
rect 18104 35232 18110 35284
rect 18690 35272 18696 35284
rect 18651 35244 18696 35272
rect 18690 35232 18696 35244
rect 18748 35232 18754 35284
rect 21082 35272 21088 35284
rect 21043 35244 21088 35272
rect 21082 35232 21088 35244
rect 21140 35272 21146 35284
rect 22189 35275 22247 35281
rect 22189 35272 22201 35275
rect 21140 35244 22201 35272
rect 21140 35232 21146 35244
rect 22189 35241 22201 35244
rect 22235 35241 22247 35275
rect 22189 35235 22247 35241
rect 21637 35207 21695 35213
rect 21637 35204 21649 35207
rect 13228 35176 15424 35204
rect 15488 35176 21649 35204
rect 13228 35164 13234 35176
rect 11664 35108 12204 35136
rect 11664 35096 11670 35108
rect 12710 35096 12716 35148
rect 12768 35136 12774 35148
rect 12768 35108 14320 35136
rect 12768 35096 12774 35108
rect 4370 35040 4476 35068
rect 5721 35071 5779 35077
rect 5721 35037 5733 35071
rect 5767 35068 5779 35071
rect 6270 35068 6276 35080
rect 5767 35040 6276 35068
rect 5767 35037 5779 35040
rect 5721 35031 5779 35037
rect 1946 35000 1952 35012
rect 1907 34972 1952 35000
rect 1946 34960 1952 34972
rect 2004 34960 2010 35012
rect 4062 35000 4068 35012
rect 3174 34972 4068 35000
rect 4062 34960 4068 34972
rect 4120 34960 4126 35012
rect 5350 34960 5356 35012
rect 5408 35000 5414 35012
rect 5736 35000 5764 35031
rect 6270 35028 6276 35040
rect 6328 35028 6334 35080
rect 8110 35028 8116 35080
rect 8168 35068 8174 35080
rect 9122 35068 9128 35080
rect 8168 35040 8432 35068
rect 9083 35040 9128 35068
rect 8168 35028 8174 35040
rect 5408 34972 5764 35000
rect 5408 34960 5414 34972
rect 5810 34960 5816 35012
rect 5868 35000 5874 35012
rect 6546 35000 6552 35012
rect 5868 34972 6552 35000
rect 5868 34960 5874 34972
rect 6546 34960 6552 34972
rect 6604 34960 6610 35012
rect 8018 35000 8024 35012
rect 7774 34972 8024 35000
rect 8018 34960 8024 34972
rect 8076 34960 8082 35012
rect 8294 35000 8300 35012
rect 8255 34972 8300 35000
rect 8294 34960 8300 34972
rect 8352 34960 8358 35012
rect 8404 35000 8432 35040
rect 9122 35028 9128 35040
rect 9180 35068 9186 35080
rect 10778 35068 10784 35080
rect 9180 35040 10784 35068
rect 9180 35028 9186 35040
rect 10778 35028 10784 35040
rect 10836 35028 10842 35080
rect 13541 35071 13599 35077
rect 13541 35037 13553 35071
rect 13587 35068 13599 35071
rect 13906 35068 13912 35080
rect 13587 35040 13912 35068
rect 13587 35037 13599 35040
rect 13541 35031 13599 35037
rect 13906 35028 13912 35040
rect 13964 35068 13970 35080
rect 14292 35077 14320 35108
rect 15396 35077 15424 35176
rect 21637 35173 21649 35176
rect 21683 35173 21695 35207
rect 21637 35167 21695 35173
rect 19981 35139 20039 35145
rect 19981 35136 19993 35139
rect 15481 35108 19993 35136
rect 14277 35071 14335 35077
rect 13964 35040 14136 35068
rect 13964 35028 13970 35040
rect 10870 35000 10876 35012
rect 8404 34972 10876 35000
rect 10870 34960 10876 34972
rect 10928 34960 10934 35012
rect 11146 35000 11152 35012
rect 11107 34972 11152 35000
rect 11146 34960 11152 34972
rect 11204 34960 11210 35012
rect 11238 34960 11244 35012
rect 11296 35000 11302 35012
rect 11296 34972 11638 35000
rect 11296 34960 11302 34972
rect 12434 34960 12440 35012
rect 12492 35000 12498 35012
rect 12897 35003 12955 35009
rect 12897 35000 12909 35003
rect 12492 34972 12909 35000
rect 12492 34960 12498 34972
rect 12897 34969 12909 34972
rect 12943 35000 12955 35003
rect 13998 35000 14004 35012
rect 12943 34972 14004 35000
rect 12943 34969 12955 34972
rect 12897 34963 12955 34969
rect 13998 34960 14004 34972
rect 14056 34960 14062 35012
rect 14108 35000 14136 35040
rect 14277 35037 14289 35071
rect 14323 35037 14335 35071
rect 14277 35031 14335 35037
rect 15381 35071 15439 35077
rect 15381 35037 15393 35071
rect 15427 35037 15439 35071
rect 15381 35031 15439 35037
rect 15481 35000 15509 35108
rect 19981 35105 19993 35108
rect 20027 35105 20039 35139
rect 19981 35099 20039 35105
rect 20346 35096 20352 35148
rect 20404 35136 20410 35148
rect 20533 35139 20591 35145
rect 20533 35136 20545 35139
rect 20404 35108 20545 35136
rect 20404 35096 20410 35108
rect 20533 35105 20545 35108
rect 20579 35105 20591 35139
rect 20533 35099 20591 35105
rect 16114 35068 16120 35080
rect 16075 35040 16120 35068
rect 16114 35028 16120 35040
rect 16172 35028 16178 35080
rect 16206 35028 16212 35080
rect 16264 35068 16270 35080
rect 16853 35071 16911 35077
rect 16264 35040 16309 35068
rect 16264 35028 16270 35040
rect 16853 35037 16865 35071
rect 16899 35037 16911 35071
rect 16853 35031 16911 35037
rect 16945 35071 17003 35077
rect 16945 35037 16957 35071
rect 16991 35068 17003 35071
rect 18690 35068 18696 35080
rect 16991 35040 18696 35068
rect 16991 35037 17003 35040
rect 16945 35031 17003 35037
rect 14108 34972 15509 35000
rect 15562 34960 15568 35012
rect 15620 35000 15626 35012
rect 16868 35000 16896 35031
rect 18690 35028 18696 35040
rect 18748 35028 18754 35080
rect 18785 35071 18843 35077
rect 18785 35037 18797 35071
rect 18831 35068 18843 35071
rect 19242 35068 19248 35080
rect 18831 35040 19248 35068
rect 18831 35037 18843 35040
rect 18785 35031 18843 35037
rect 19242 35028 19248 35040
rect 19300 35028 19306 35080
rect 15620 34972 16896 35000
rect 15620 34960 15626 34972
rect 17310 34960 17316 35012
rect 17368 35000 17374 35012
rect 17773 35003 17831 35009
rect 17773 35000 17785 35003
rect 17368 34972 17785 35000
rect 17368 34960 17374 34972
rect 17773 34969 17785 34972
rect 17819 35000 17831 35003
rect 17862 35000 17868 35012
rect 17819 34972 17868 35000
rect 17819 34969 17831 34972
rect 17773 34963 17831 34969
rect 17862 34960 17868 34972
rect 17920 34960 17926 35012
rect 17954 34960 17960 35012
rect 18012 35000 18018 35012
rect 22741 35003 22799 35009
rect 22741 35000 22753 35003
rect 18012 34972 22753 35000
rect 18012 34960 18018 34972
rect 22741 34969 22753 34972
rect 22787 34969 22799 35003
rect 22741 34963 22799 34969
rect 23014 34960 23020 35012
rect 23072 35000 23078 35012
rect 24581 35003 24639 35009
rect 24581 35000 24593 35003
rect 23072 34972 24593 35000
rect 23072 34960 23078 34972
rect 24581 34969 24593 34972
rect 24627 34969 24639 35003
rect 24581 34963 24639 34969
rect 3786 34892 3792 34944
rect 3844 34932 3850 34944
rect 3973 34935 4031 34941
rect 3973 34932 3985 34935
rect 3844 34904 3985 34932
rect 3844 34892 3850 34904
rect 3973 34901 3985 34904
rect 4019 34901 4031 34935
rect 3973 34895 4031 34901
rect 5626 34892 5632 34944
rect 5684 34932 5690 34944
rect 12710 34932 12716 34944
rect 5684 34904 12716 34932
rect 5684 34892 5690 34904
rect 12710 34892 12716 34904
rect 12768 34892 12774 34944
rect 13633 34935 13691 34941
rect 13633 34901 13645 34935
rect 13679 34932 13691 34935
rect 14090 34932 14096 34944
rect 13679 34904 14096 34932
rect 13679 34901 13691 34904
rect 13633 34895 13691 34901
rect 14090 34892 14096 34904
rect 14148 34892 14154 34944
rect 14369 34935 14427 34941
rect 14369 34901 14381 34935
rect 14415 34932 14427 34935
rect 15286 34932 15292 34944
rect 14415 34904 15292 34932
rect 14415 34901 14427 34904
rect 14369 34895 14427 34901
rect 15286 34892 15292 34904
rect 15344 34892 15350 34944
rect 15473 34935 15531 34941
rect 15473 34901 15485 34935
rect 15519 34932 15531 34935
rect 16850 34932 16856 34944
rect 15519 34904 16856 34932
rect 15519 34901 15531 34904
rect 15473 34895 15531 34901
rect 16850 34892 16856 34904
rect 16908 34892 16914 34944
rect 17034 34892 17040 34944
rect 17092 34932 17098 34944
rect 19521 34935 19579 34941
rect 19521 34932 19533 34935
rect 17092 34904 19533 34932
rect 17092 34892 17098 34904
rect 19521 34901 19533 34904
rect 19567 34932 19579 34935
rect 20438 34932 20444 34944
rect 19567 34904 20444 34932
rect 19567 34901 19579 34904
rect 19521 34895 19579 34901
rect 20438 34892 20444 34904
rect 20496 34892 20502 34944
rect 21358 34892 21364 34944
rect 21416 34932 21422 34944
rect 23293 34935 23351 34941
rect 23293 34932 23305 34935
rect 21416 34904 23305 34932
rect 21416 34892 21422 34904
rect 23293 34901 23305 34904
rect 23339 34901 23351 34935
rect 23293 34895 23351 34901
rect 23382 34892 23388 34944
rect 23440 34932 23446 34944
rect 23845 34935 23903 34941
rect 23845 34932 23857 34935
rect 23440 34904 23857 34932
rect 23440 34892 23446 34904
rect 23845 34901 23857 34904
rect 23891 34901 23903 34935
rect 23845 34895 23903 34901
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 12710 34728 12716 34740
rect 4632 34700 12716 34728
rect 4632 34660 4660 34700
rect 12710 34688 12716 34700
rect 12768 34688 12774 34740
rect 12802 34688 12808 34740
rect 12860 34728 12866 34740
rect 18230 34728 18236 34740
rect 12860 34700 18236 34728
rect 12860 34688 12866 34700
rect 18230 34688 18236 34700
rect 18288 34688 18294 34740
rect 19150 34728 19156 34740
rect 19111 34700 19156 34728
rect 19150 34688 19156 34700
rect 19208 34688 19214 34740
rect 20349 34731 20407 34737
rect 20349 34697 20361 34731
rect 20395 34728 20407 34731
rect 20809 34731 20867 34737
rect 20809 34728 20821 34731
rect 20395 34700 20821 34728
rect 20395 34697 20407 34700
rect 20349 34691 20407 34697
rect 20809 34697 20821 34700
rect 20855 34728 20867 34731
rect 21082 34728 21088 34740
rect 20855 34700 21088 34728
rect 20855 34697 20867 34700
rect 20809 34691 20867 34697
rect 21082 34688 21088 34700
rect 21140 34728 21146 34740
rect 22557 34731 22615 34737
rect 22557 34728 22569 34731
rect 21140 34700 22569 34728
rect 21140 34688 21146 34700
rect 22557 34697 22569 34700
rect 22603 34728 22615 34731
rect 22922 34728 22928 34740
rect 22603 34700 22928 34728
rect 22603 34697 22615 34700
rect 22557 34691 22615 34697
rect 22922 34688 22928 34700
rect 22980 34728 22986 34740
rect 23382 34728 23388 34740
rect 22980 34700 23388 34728
rect 22980 34688 22986 34700
rect 23382 34688 23388 34700
rect 23440 34728 23446 34740
rect 23661 34731 23719 34737
rect 23661 34728 23673 34731
rect 23440 34700 23673 34728
rect 23440 34688 23446 34700
rect 23661 34697 23673 34700
rect 23707 34728 23719 34731
rect 24213 34731 24271 34737
rect 24213 34728 24225 34731
rect 23707 34700 24225 34728
rect 23707 34697 23719 34700
rect 23661 34691 23719 34697
rect 24213 34697 24225 34700
rect 24259 34697 24271 34731
rect 24213 34691 24271 34697
rect 7282 34660 7288 34672
rect 3266 34632 4660 34660
rect 6196 34632 7288 34660
rect 1670 34552 1676 34604
rect 1728 34592 1734 34604
rect 1765 34595 1823 34601
rect 1765 34592 1777 34595
rect 1728 34564 1777 34592
rect 1728 34552 1734 34564
rect 1765 34561 1777 34564
rect 1811 34561 1823 34595
rect 1765 34555 1823 34561
rect 3878 34552 3884 34604
rect 3936 34592 3942 34604
rect 3973 34595 4031 34601
rect 3973 34592 3985 34595
rect 3936 34564 3985 34592
rect 3936 34552 3942 34564
rect 3973 34561 3985 34564
rect 4019 34561 4031 34595
rect 3973 34555 4031 34561
rect 5350 34552 5356 34604
rect 5408 34552 5414 34604
rect 3513 34527 3571 34533
rect 3513 34493 3525 34527
rect 3559 34524 3571 34527
rect 6196 34524 6224 34632
rect 7282 34620 7288 34632
rect 7340 34620 7346 34672
rect 9122 34660 9128 34672
rect 8312 34632 9128 34660
rect 6270 34552 6276 34604
rect 6328 34592 6334 34604
rect 6733 34595 6791 34601
rect 6733 34592 6745 34595
rect 6328 34564 6745 34592
rect 6328 34552 6334 34564
rect 6733 34561 6745 34564
rect 6779 34561 6791 34595
rect 6733 34555 6791 34561
rect 8110 34552 8116 34604
rect 8168 34552 8174 34604
rect 3559 34496 6224 34524
rect 3559 34493 3571 34496
rect 3513 34487 3571 34493
rect 7098 34484 7104 34536
rect 7156 34524 7162 34536
rect 8312 34524 8340 34632
rect 9122 34620 9128 34632
rect 9180 34620 9186 34672
rect 12250 34660 12256 34672
rect 10442 34632 12256 34660
rect 12250 34620 12256 34632
rect 12308 34620 12314 34672
rect 12434 34620 12440 34672
rect 12492 34620 12498 34672
rect 14093 34663 14151 34669
rect 14093 34629 14105 34663
rect 14139 34660 14151 34663
rect 15010 34660 15016 34672
rect 14139 34632 15016 34660
rect 14139 34629 14151 34632
rect 14093 34623 14151 34629
rect 15010 34620 15016 34632
rect 15068 34620 15074 34672
rect 16209 34663 16267 34669
rect 16209 34629 16221 34663
rect 16255 34660 16267 34663
rect 17586 34660 17592 34672
rect 16255 34632 17592 34660
rect 16255 34629 16267 34632
rect 16209 34623 16267 34629
rect 17586 34620 17592 34632
rect 17644 34620 17650 34672
rect 18046 34660 18052 34672
rect 17880 34632 18052 34660
rect 10502 34552 10508 34604
rect 10560 34592 10566 34604
rect 10965 34595 11023 34601
rect 10965 34592 10977 34595
rect 10560 34564 10977 34592
rect 10560 34552 10566 34564
rect 10965 34561 10977 34564
rect 11011 34561 11023 34595
rect 10965 34555 11023 34561
rect 11514 34552 11520 34604
rect 11572 34592 11578 34604
rect 11701 34595 11759 34601
rect 11701 34592 11713 34595
rect 11572 34564 11713 34592
rect 11572 34552 11578 34564
rect 11701 34561 11713 34564
rect 11747 34561 11759 34595
rect 11701 34555 11759 34561
rect 15102 34552 15108 34604
rect 15160 34592 15166 34604
rect 15473 34595 15531 34601
rect 15473 34592 15485 34595
rect 15160 34564 15485 34592
rect 15160 34552 15166 34564
rect 15473 34561 15485 34564
rect 15519 34561 15531 34595
rect 15473 34555 15531 34561
rect 15654 34552 15660 34604
rect 15712 34592 15718 34604
rect 16117 34595 16175 34601
rect 16117 34592 16129 34595
rect 15712 34564 16129 34592
rect 15712 34552 15718 34564
rect 16117 34561 16129 34564
rect 16163 34561 16175 34595
rect 16117 34555 16175 34561
rect 17313 34595 17371 34601
rect 17313 34561 17325 34595
rect 17359 34592 17371 34595
rect 17880 34592 17908 34632
rect 18046 34620 18052 34632
rect 18104 34620 18110 34672
rect 23106 34660 23112 34672
rect 18156 34632 20852 34660
rect 23067 34632 23112 34660
rect 17359 34564 17908 34592
rect 17359 34561 17371 34564
rect 17313 34555 17371 34561
rect 17954 34552 17960 34604
rect 18012 34592 18018 34604
rect 18156 34592 18184 34632
rect 20824 34604 20852 34632
rect 23106 34620 23112 34632
rect 23164 34620 23170 34672
rect 18012 34564 18184 34592
rect 18012 34552 18018 34564
rect 18230 34552 18236 34604
rect 18288 34592 18294 34604
rect 18417 34595 18475 34601
rect 18417 34592 18429 34595
rect 18288 34564 18429 34592
rect 18288 34552 18294 34564
rect 18417 34561 18429 34564
rect 18463 34561 18475 34595
rect 19242 34592 19248 34604
rect 19203 34564 19248 34592
rect 18417 34555 18475 34561
rect 19242 34552 19248 34564
rect 19300 34592 19306 34604
rect 19705 34595 19763 34601
rect 19705 34592 19717 34595
rect 19300 34564 19717 34592
rect 19300 34552 19306 34564
rect 19705 34561 19717 34564
rect 19751 34592 19763 34595
rect 20714 34592 20720 34604
rect 19751 34564 20720 34592
rect 19751 34561 19763 34564
rect 19705 34555 19763 34561
rect 20714 34552 20720 34564
rect 20772 34552 20778 34604
rect 20806 34552 20812 34604
rect 20864 34552 20870 34604
rect 7156 34496 8340 34524
rect 8481 34527 8539 34533
rect 7156 34484 7162 34496
rect 8481 34493 8493 34527
rect 8527 34524 8539 34527
rect 8570 34524 8576 34536
rect 8527 34496 8576 34524
rect 8527 34493 8539 34496
rect 8481 34487 8539 34493
rect 8570 34484 8576 34496
rect 8628 34484 8634 34536
rect 8938 34524 8944 34536
rect 8899 34496 8944 34524
rect 8938 34484 8944 34496
rect 8996 34484 9002 34536
rect 9582 34484 9588 34536
rect 9640 34524 9646 34536
rect 9766 34524 9772 34536
rect 9640 34496 9772 34524
rect 9640 34484 9646 34496
rect 9766 34484 9772 34496
rect 9824 34484 9830 34536
rect 9858 34484 9864 34536
rect 9916 34524 9922 34536
rect 11977 34527 12035 34533
rect 9916 34496 11008 34524
rect 9916 34484 9922 34496
rect 3786 34456 3792 34468
rect 3436 34428 3792 34456
rect 2028 34391 2086 34397
rect 2028 34357 2040 34391
rect 2074 34388 2086 34391
rect 3436 34388 3464 34428
rect 3786 34416 3792 34428
rect 3844 34416 3850 34468
rect 5721 34459 5779 34465
rect 5721 34425 5733 34459
rect 5767 34456 5779 34459
rect 6454 34456 6460 34468
rect 5767 34428 6460 34456
rect 5767 34425 5779 34428
rect 5721 34419 5779 34425
rect 6454 34416 6460 34428
rect 6512 34416 6518 34468
rect 2074 34360 3464 34388
rect 4236 34391 4294 34397
rect 2074 34357 2086 34360
rect 2028 34351 2086 34357
rect 4236 34357 4248 34391
rect 4282 34388 4294 34391
rect 5626 34388 5632 34400
rect 4282 34360 5632 34388
rect 4282 34357 4294 34360
rect 4236 34351 4294 34357
rect 5626 34348 5632 34360
rect 5684 34348 5690 34400
rect 6178 34348 6184 34400
rect 6236 34388 6242 34400
rect 6990 34391 7048 34397
rect 6990 34388 7002 34391
rect 6236 34360 7002 34388
rect 6236 34348 6242 34360
rect 6990 34357 7002 34360
rect 7036 34357 7048 34391
rect 6990 34351 7048 34357
rect 7374 34348 7380 34400
rect 7432 34388 7438 34400
rect 8386 34388 8392 34400
rect 7432 34360 8392 34388
rect 7432 34348 7438 34360
rect 8386 34348 8392 34360
rect 8444 34348 8450 34400
rect 9204 34391 9262 34397
rect 9204 34357 9216 34391
rect 9250 34388 9262 34391
rect 10686 34388 10692 34400
rect 9250 34360 10692 34388
rect 9250 34357 9262 34360
rect 9204 34351 9262 34357
rect 10686 34348 10692 34360
rect 10744 34348 10750 34400
rect 10980 34388 11008 34496
rect 11977 34493 11989 34527
rect 12023 34524 12035 34527
rect 12066 34524 12072 34536
rect 12023 34496 12072 34524
rect 12023 34493 12035 34496
rect 11977 34487 12035 34493
rect 12066 34484 12072 34496
rect 12124 34484 12130 34536
rect 12342 34484 12348 34536
rect 12400 34524 12406 34536
rect 12400 34496 13032 34524
rect 12400 34484 12406 34496
rect 13004 34456 13032 34496
rect 13170 34484 13176 34536
rect 13228 34524 13234 34536
rect 13449 34527 13507 34533
rect 13449 34524 13461 34527
rect 13228 34496 13461 34524
rect 13228 34484 13234 34496
rect 13449 34493 13461 34496
rect 13495 34493 13507 34527
rect 13449 34487 13507 34493
rect 14001 34527 14059 34533
rect 14001 34493 14013 34527
rect 14047 34524 14059 34527
rect 14274 34524 14280 34536
rect 14047 34496 14280 34524
rect 14047 34493 14059 34496
rect 14001 34487 14059 34493
rect 14274 34484 14280 34496
rect 14332 34484 14338 34536
rect 14458 34524 14464 34536
rect 14419 34496 14464 34524
rect 14458 34484 14464 34496
rect 14516 34484 14522 34536
rect 15565 34527 15623 34533
rect 15565 34493 15577 34527
rect 15611 34524 15623 34527
rect 15746 34524 15752 34536
rect 15611 34496 15752 34524
rect 15611 34493 15623 34496
rect 15565 34487 15623 34493
rect 15746 34484 15752 34496
rect 15804 34484 15810 34536
rect 16574 34484 16580 34536
rect 16632 34524 16638 34536
rect 17037 34527 17095 34533
rect 17037 34524 17049 34527
rect 16632 34496 17049 34524
rect 16632 34484 16638 34496
rect 17037 34493 17049 34496
rect 17083 34493 17095 34527
rect 17037 34487 17095 34493
rect 17126 34484 17132 34536
rect 17184 34524 17190 34536
rect 17865 34527 17923 34533
rect 17865 34524 17877 34527
rect 17184 34496 17877 34524
rect 17184 34484 17190 34496
rect 17865 34493 17877 34496
rect 17911 34493 17923 34527
rect 17865 34487 17923 34493
rect 18509 34527 18567 34533
rect 18509 34493 18521 34527
rect 18555 34524 18567 34527
rect 19978 34524 19984 34536
rect 18555 34496 19984 34524
rect 18555 34493 18567 34496
rect 18509 34487 18567 34493
rect 19978 34484 19984 34496
rect 20036 34484 20042 34536
rect 20070 34484 20076 34536
rect 20128 34524 20134 34536
rect 21361 34527 21419 34533
rect 21361 34524 21373 34527
rect 20128 34496 21373 34524
rect 20128 34484 20134 34496
rect 21361 34493 21373 34496
rect 21407 34493 21419 34527
rect 21361 34487 21419 34493
rect 22005 34459 22063 34465
rect 22005 34456 22017 34459
rect 13004 34428 22017 34456
rect 22005 34425 22017 34428
rect 22051 34425 22063 34459
rect 22005 34419 22063 34425
rect 19058 34388 19064 34400
rect 10980 34360 19064 34388
rect 19058 34348 19064 34360
rect 19116 34348 19122 34400
rect 19150 34348 19156 34400
rect 19208 34388 19214 34400
rect 21910 34388 21916 34400
rect 19208 34360 21916 34388
rect 19208 34348 19214 34360
rect 21910 34348 21916 34360
rect 21968 34348 21974 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 6638 34144 6644 34196
rect 6696 34184 6702 34196
rect 8202 34184 8208 34196
rect 6696 34156 8208 34184
rect 6696 34144 6702 34156
rect 8202 34144 8208 34156
rect 8260 34144 8266 34196
rect 8294 34144 8300 34196
rect 8352 34184 8358 34196
rect 9388 34187 9446 34193
rect 9388 34184 9400 34187
rect 8352 34156 9400 34184
rect 8352 34144 8358 34156
rect 9388 34153 9400 34156
rect 9434 34184 9446 34187
rect 12250 34184 12256 34196
rect 9434 34156 12256 34184
rect 9434 34153 9446 34156
rect 9388 34147 9446 34153
rect 12250 34144 12256 34156
rect 12308 34144 12314 34196
rect 12342 34144 12348 34196
rect 12400 34184 12406 34196
rect 12400 34156 12940 34184
rect 12400 34144 12406 34156
rect 11422 34116 11428 34128
rect 7668 34088 9260 34116
rect 3421 34051 3479 34057
rect 3421 34017 3433 34051
rect 3467 34048 3479 34051
rect 3510 34048 3516 34060
rect 3467 34020 3516 34048
rect 3467 34017 3479 34020
rect 3421 34011 3479 34017
rect 3510 34008 3516 34020
rect 3568 34048 3574 34060
rect 3878 34048 3884 34060
rect 3568 34020 3884 34048
rect 3568 34008 3574 34020
rect 3878 34008 3884 34020
rect 3936 34048 3942 34060
rect 3973 34051 4031 34057
rect 3973 34048 3985 34051
rect 3936 34020 3985 34048
rect 3936 34008 3942 34020
rect 3973 34017 3985 34020
rect 4019 34017 4031 34051
rect 3973 34011 4031 34017
rect 5718 33940 5724 33992
rect 5776 33980 5782 33992
rect 6273 33983 6331 33989
rect 6273 33980 6285 33983
rect 5776 33952 6285 33980
rect 5776 33940 5782 33952
rect 6273 33949 6285 33952
rect 6319 33949 6331 33983
rect 7668 33966 7696 34088
rect 8938 34008 8944 34060
rect 8996 34048 9002 34060
rect 9125 34051 9183 34057
rect 9125 34048 9137 34051
rect 8996 34020 9137 34048
rect 8996 34008 9002 34020
rect 9125 34017 9137 34020
rect 9171 34017 9183 34051
rect 9232 34048 9260 34088
rect 10428 34088 11428 34116
rect 10428 34048 10456 34088
rect 11422 34076 11428 34088
rect 11480 34076 11486 34128
rect 12912 34116 12940 34156
rect 16206 34144 16212 34196
rect 16264 34184 16270 34196
rect 17218 34184 17224 34196
rect 16264 34156 17224 34184
rect 16264 34144 16270 34156
rect 17218 34144 17224 34156
rect 17276 34144 17282 34196
rect 19058 34144 19064 34196
rect 19116 34184 19122 34196
rect 20165 34187 20223 34193
rect 20165 34184 20177 34187
rect 19116 34156 20177 34184
rect 19116 34144 19122 34156
rect 20165 34153 20177 34156
rect 20211 34153 20223 34187
rect 20165 34147 20223 34153
rect 21082 34144 21088 34196
rect 21140 34184 21146 34196
rect 21269 34187 21327 34193
rect 21269 34184 21281 34187
rect 21140 34156 21281 34184
rect 21140 34144 21146 34156
rect 21269 34153 21281 34156
rect 21315 34153 21327 34187
rect 22922 34184 22928 34196
rect 22883 34156 22928 34184
rect 21269 34147 21327 34153
rect 22922 34144 22928 34156
rect 22980 34184 22986 34196
rect 23477 34187 23535 34193
rect 23477 34184 23489 34187
rect 22980 34156 23489 34184
rect 22980 34144 22986 34156
rect 23477 34153 23489 34156
rect 23523 34184 23535 34187
rect 24581 34187 24639 34193
rect 24581 34184 24593 34187
rect 23523 34156 24593 34184
rect 23523 34153 23535 34156
rect 23477 34147 23535 34153
rect 24581 34153 24593 34156
rect 24627 34153 24639 34187
rect 24581 34147 24639 34153
rect 14366 34116 14372 34128
rect 12912 34088 14372 34116
rect 14366 34076 14372 34088
rect 14424 34076 14430 34128
rect 14458 34076 14464 34128
rect 14516 34116 14522 34128
rect 14516 34088 18644 34116
rect 14516 34076 14522 34088
rect 18616 34060 18644 34088
rect 19150 34076 19156 34128
rect 19208 34116 19214 34128
rect 19208 34088 20392 34116
rect 19208 34076 19214 34088
rect 9232 34020 10456 34048
rect 9125 34011 9183 34017
rect 10686 34008 10692 34060
rect 10744 34048 10750 34060
rect 11149 34051 11207 34057
rect 11149 34048 11161 34051
rect 10744 34020 11161 34048
rect 10744 34008 10750 34020
rect 11149 34017 11161 34020
rect 11195 34017 11207 34051
rect 11606 34048 11612 34060
rect 11567 34020 11612 34048
rect 11149 34011 11207 34017
rect 11606 34008 11612 34020
rect 11664 34008 11670 34060
rect 12250 34008 12256 34060
rect 12308 34048 12314 34060
rect 12526 34048 12532 34060
rect 12308 34020 12532 34048
rect 12308 34008 12314 34020
rect 12526 34008 12532 34020
rect 12584 34008 12590 34060
rect 12618 34008 12624 34060
rect 12676 34048 12682 34060
rect 16485 34051 16543 34057
rect 16485 34048 16497 34051
rect 12676 34020 16497 34048
rect 12676 34008 12682 34020
rect 16485 34017 16497 34020
rect 16531 34017 16543 34051
rect 17034 34048 17040 34060
rect 16485 34011 16543 34017
rect 16776 34020 17040 34048
rect 10778 33980 10784 33992
rect 6273 33943 6331 33949
rect 8220 33952 9168 33980
rect 10534 33952 10784 33980
rect 2130 33872 2136 33924
rect 2188 33872 2194 33924
rect 3145 33915 3203 33921
rect 3145 33881 3157 33915
rect 3191 33881 3203 33915
rect 4246 33912 4252 33924
rect 4207 33884 4252 33912
rect 3145 33875 3203 33881
rect 1578 33804 1584 33856
rect 1636 33844 1642 33856
rect 1673 33847 1731 33853
rect 1673 33844 1685 33847
rect 1636 33816 1685 33844
rect 1636 33804 1642 33816
rect 1673 33813 1685 33816
rect 1719 33813 1731 33847
rect 3160 33844 3188 33875
rect 4246 33872 4252 33884
rect 4304 33872 4310 33924
rect 4982 33872 4988 33924
rect 5040 33872 5046 33924
rect 5810 33912 5816 33924
rect 5644 33884 5816 33912
rect 5644 33844 5672 33884
rect 5810 33872 5816 33884
rect 5868 33872 5874 33924
rect 6454 33872 6460 33924
rect 6512 33912 6518 33924
rect 6549 33915 6607 33921
rect 6549 33912 6561 33915
rect 6512 33884 6561 33912
rect 6512 33872 6518 33884
rect 6549 33881 6561 33884
rect 6595 33881 6607 33915
rect 6549 33875 6607 33881
rect 3160 33816 5672 33844
rect 5721 33847 5779 33853
rect 1673 33807 1731 33813
rect 5721 33813 5733 33847
rect 5767 33844 5779 33847
rect 8220 33844 8248 33952
rect 9140 33924 9168 33952
rect 10778 33940 10784 33952
rect 10836 33940 10842 33992
rect 14550 33980 14556 33992
rect 13018 33952 14556 33980
rect 14550 33940 14556 33952
rect 14608 33940 14614 33992
rect 15654 33940 15660 33992
rect 15712 33980 15718 33992
rect 16776 33989 16804 34020
rect 17034 34008 17040 34020
rect 17092 34048 17098 34060
rect 17092 34020 18092 34048
rect 17092 34008 17098 34020
rect 18064 33992 18092 34020
rect 18598 34008 18604 34060
rect 18656 34048 18662 34060
rect 19886 34048 19892 34060
rect 18656 34020 19892 34048
rect 18656 34008 18662 34020
rect 19886 34008 19892 34020
rect 19944 34008 19950 34060
rect 16761 33983 16819 33989
rect 15712 33952 16712 33980
rect 15712 33940 15718 33952
rect 8297 33915 8355 33921
rect 8297 33881 8309 33915
rect 8343 33912 8355 33915
rect 8478 33912 8484 33924
rect 8343 33884 8484 33912
rect 8343 33881 8355 33884
rect 8297 33875 8355 33881
rect 8478 33872 8484 33884
rect 8536 33872 8542 33924
rect 9122 33872 9128 33924
rect 9180 33872 9186 33924
rect 11885 33915 11943 33921
rect 11885 33912 11897 33915
rect 10704 33884 11897 33912
rect 5767 33816 8248 33844
rect 5767 33813 5779 33816
rect 5721 33807 5779 33813
rect 8570 33804 8576 33856
rect 8628 33844 8634 33856
rect 9030 33844 9036 33856
rect 8628 33816 9036 33844
rect 8628 33804 8634 33816
rect 9030 33804 9036 33816
rect 9088 33844 9094 33856
rect 10704 33844 10732 33884
rect 11885 33881 11897 33884
rect 11931 33881 11943 33915
rect 14458 33912 14464 33924
rect 14419 33884 14464 33912
rect 11885 33875 11943 33881
rect 14458 33872 14464 33884
rect 14516 33872 14522 33924
rect 15378 33912 15384 33924
rect 15339 33884 15384 33912
rect 15378 33872 15384 33884
rect 15436 33872 15442 33924
rect 15473 33915 15531 33921
rect 15473 33881 15485 33915
rect 15519 33912 15531 33915
rect 15930 33912 15936 33924
rect 15519 33884 15936 33912
rect 15519 33881 15531 33884
rect 15473 33875 15531 33881
rect 15930 33872 15936 33884
rect 15988 33872 15994 33924
rect 16684 33912 16712 33952
rect 16761 33949 16773 33983
rect 16807 33949 16819 33983
rect 16761 33943 16819 33949
rect 17221 33983 17279 33989
rect 17221 33949 17233 33983
rect 17267 33980 17279 33983
rect 17310 33980 17316 33992
rect 17267 33952 17316 33980
rect 17267 33949 17279 33952
rect 17221 33943 17279 33949
rect 17310 33940 17316 33952
rect 17368 33940 17374 33992
rect 17497 33983 17555 33989
rect 17497 33949 17509 33983
rect 17543 33980 17555 33983
rect 17954 33980 17960 33992
rect 17543 33952 17960 33980
rect 17543 33949 17555 33952
rect 17497 33943 17555 33949
rect 17954 33940 17960 33952
rect 18012 33940 18018 33992
rect 18046 33940 18052 33992
rect 18104 33980 18110 33992
rect 18141 33983 18199 33989
rect 18141 33980 18153 33983
rect 18104 33952 18153 33980
rect 18104 33940 18110 33952
rect 18141 33949 18153 33952
rect 18187 33949 18199 33983
rect 20162 33980 20168 33992
rect 18141 33943 18199 33949
rect 18432 33952 20168 33980
rect 18432 33921 18460 33952
rect 20162 33940 20168 33952
rect 20220 33940 20226 33992
rect 20257 33983 20315 33989
rect 20257 33949 20269 33983
rect 20303 33980 20315 33983
rect 20364 33980 20392 34088
rect 20622 34008 20628 34060
rect 20680 34048 20686 34060
rect 31662 34048 31668 34060
rect 20680 34020 31668 34048
rect 20680 34008 20686 34020
rect 31662 34008 31668 34020
rect 31720 34008 31726 34060
rect 20303 33952 20392 33980
rect 20303 33949 20315 33952
rect 20257 33943 20315 33949
rect 18417 33915 18475 33921
rect 18417 33912 18429 33915
rect 16684 33884 18429 33912
rect 18417 33881 18429 33884
rect 18463 33881 18475 33915
rect 20717 33915 20775 33921
rect 20717 33912 20729 33915
rect 18417 33875 18475 33881
rect 18524 33884 20729 33912
rect 9088 33816 10732 33844
rect 9088 33804 9094 33816
rect 10778 33804 10784 33856
rect 10836 33844 10842 33856
rect 12710 33844 12716 33856
rect 10836 33816 12716 33844
rect 10836 33804 10842 33816
rect 12710 33804 12716 33816
rect 12768 33804 12774 33856
rect 13262 33804 13268 33856
rect 13320 33844 13326 33856
rect 13357 33847 13415 33853
rect 13357 33844 13369 33847
rect 13320 33816 13369 33844
rect 13320 33804 13326 33816
rect 13357 33813 13369 33816
rect 13403 33813 13415 33847
rect 13357 33807 13415 33813
rect 13446 33804 13452 33856
rect 13504 33844 13510 33856
rect 18524 33844 18552 33884
rect 20717 33881 20729 33884
rect 20763 33881 20775 33915
rect 22002 33912 22008 33924
rect 20717 33875 20775 33881
rect 20824 33884 22008 33912
rect 13504 33816 18552 33844
rect 13504 33804 13510 33816
rect 19058 33804 19064 33856
rect 19116 33844 19122 33856
rect 19429 33847 19487 33853
rect 19429 33844 19441 33847
rect 19116 33816 19441 33844
rect 19116 33804 19122 33816
rect 19429 33813 19441 33816
rect 19475 33813 19487 33847
rect 19429 33807 19487 33813
rect 19518 33804 19524 33856
rect 19576 33844 19582 33856
rect 20824 33844 20852 33884
rect 22002 33872 22008 33884
rect 22060 33912 22066 33924
rect 22373 33915 22431 33921
rect 22373 33912 22385 33915
rect 22060 33884 22385 33912
rect 22060 33872 22066 33884
rect 22373 33881 22385 33884
rect 22419 33881 22431 33915
rect 22373 33875 22431 33881
rect 21818 33844 21824 33856
rect 19576 33816 20852 33844
rect 21779 33816 21824 33844
rect 19576 33804 19582 33816
rect 21818 33804 21824 33816
rect 21876 33804 21882 33856
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 1854 33600 1860 33652
rect 1912 33640 1918 33652
rect 11330 33640 11336 33652
rect 1912 33612 11336 33640
rect 1912 33600 1918 33612
rect 11330 33600 11336 33612
rect 11388 33600 11394 33652
rect 15102 33640 15108 33652
rect 11440 33612 15108 33640
rect 2682 33532 2688 33584
rect 2740 33532 2746 33584
rect 5721 33575 5779 33581
rect 5721 33541 5733 33575
rect 5767 33572 5779 33575
rect 5994 33572 6000 33584
rect 5767 33544 6000 33572
rect 5767 33541 5779 33544
rect 5721 33535 5779 33541
rect 5994 33532 6000 33544
rect 6052 33572 6058 33584
rect 6822 33572 6828 33584
rect 6052 33544 6828 33572
rect 6052 33532 6058 33544
rect 6822 33532 6828 33544
rect 6880 33532 6886 33584
rect 8386 33532 8392 33584
rect 8444 33572 8450 33584
rect 8570 33572 8576 33584
rect 8444 33544 8576 33572
rect 8444 33532 8450 33544
rect 8570 33532 8576 33544
rect 8628 33572 8634 33584
rect 9401 33575 9459 33581
rect 9401 33572 9413 33575
rect 8628 33544 9413 33572
rect 8628 33532 8634 33544
rect 9401 33541 9413 33544
rect 9447 33541 9459 33575
rect 11440 33572 11468 33612
rect 15102 33600 15108 33612
rect 15160 33600 15166 33652
rect 15562 33640 15568 33652
rect 15396 33612 15568 33640
rect 11882 33572 11888 33584
rect 10626 33544 11468 33572
rect 11532 33544 11888 33572
rect 9401 33535 9459 33541
rect 3510 33464 3516 33516
rect 3568 33504 3574 33516
rect 3568 33476 3613 33504
rect 3712 33476 4646 33504
rect 3568 33464 3574 33476
rect 1765 33439 1823 33445
rect 1765 33405 1777 33439
rect 1811 33436 1823 33439
rect 1946 33436 1952 33448
rect 1811 33408 1952 33436
rect 1811 33405 1823 33408
rect 1765 33399 1823 33405
rect 1946 33396 1952 33408
rect 2004 33396 2010 33448
rect 3234 33436 3240 33448
rect 3195 33408 3240 33436
rect 3234 33396 3240 33408
rect 3292 33396 3298 33448
rect 2222 33260 2228 33312
rect 2280 33300 2286 33312
rect 3712 33300 3740 33476
rect 3973 33439 4031 33445
rect 3973 33405 3985 33439
rect 4019 33436 4031 33439
rect 4706 33436 4712 33448
rect 4019 33408 4712 33436
rect 4019 33405 4031 33408
rect 3973 33399 4031 33405
rect 4706 33396 4712 33408
rect 4764 33396 4770 33448
rect 5718 33396 5724 33448
rect 5776 33436 5782 33448
rect 5997 33439 6055 33445
rect 5997 33436 6009 33439
rect 5776 33408 6009 33436
rect 5776 33396 5782 33408
rect 5997 33405 6009 33408
rect 6043 33436 6055 33439
rect 6825 33439 6883 33445
rect 6825 33436 6837 33439
rect 6043 33408 6837 33436
rect 6043 33405 6055 33408
rect 5997 33399 6055 33405
rect 6825 33405 6837 33408
rect 6871 33405 6883 33439
rect 6825 33399 6883 33405
rect 7101 33439 7159 33445
rect 7101 33405 7113 33439
rect 7147 33436 7159 33439
rect 7834 33436 7840 33448
rect 7147 33408 7840 33436
rect 7147 33405 7159 33408
rect 7101 33399 7159 33405
rect 7834 33396 7840 33408
rect 7892 33396 7898 33448
rect 8220 33368 8248 33490
rect 8938 33464 8944 33516
rect 8996 33504 9002 33516
rect 9125 33507 9183 33513
rect 9125 33504 9137 33507
rect 8996 33476 9137 33504
rect 8996 33464 9002 33476
rect 9125 33473 9137 33476
rect 9171 33473 9183 33507
rect 9125 33467 9183 33473
rect 10778 33464 10784 33516
rect 10836 33504 10842 33516
rect 11532 33504 11560 33544
rect 11882 33532 11888 33544
rect 11940 33532 11946 33584
rect 15396 33572 15424 33612
rect 15562 33600 15568 33612
rect 15620 33600 15626 33652
rect 16390 33640 16396 33652
rect 15672 33612 16396 33640
rect 15672 33572 15700 33612
rect 16390 33600 16396 33612
rect 16448 33600 16454 33652
rect 17402 33600 17408 33652
rect 17460 33640 17466 33652
rect 20070 33640 20076 33652
rect 17460 33612 20076 33640
rect 17460 33600 17466 33612
rect 20070 33600 20076 33612
rect 20128 33600 20134 33652
rect 20714 33640 20720 33652
rect 20675 33612 20720 33640
rect 20714 33600 20720 33612
rect 20772 33600 20778 33652
rect 21910 33600 21916 33652
rect 21968 33640 21974 33652
rect 22005 33643 22063 33649
rect 22005 33640 22017 33643
rect 21968 33612 22017 33640
rect 21968 33600 21974 33612
rect 22005 33609 22017 33612
rect 22051 33609 22063 33643
rect 22005 33603 22063 33609
rect 22649 33643 22707 33649
rect 22649 33609 22661 33643
rect 22695 33640 22707 33643
rect 22922 33640 22928 33652
rect 22695 33612 22928 33640
rect 22695 33609 22707 33612
rect 22649 33603 22707 33609
rect 22922 33600 22928 33612
rect 22980 33640 22986 33652
rect 23109 33643 23167 33649
rect 23109 33640 23121 33643
rect 22980 33612 23121 33640
rect 22980 33600 22986 33612
rect 23109 33609 23121 33612
rect 23155 33640 23167 33643
rect 24213 33643 24271 33649
rect 24213 33640 24225 33643
rect 23155 33612 24225 33640
rect 23155 33609 23167 33612
rect 23109 33603 23167 33609
rect 24213 33609 24225 33612
rect 24259 33609 24271 33643
rect 24762 33640 24768 33652
rect 24723 33612 24768 33640
rect 24213 33603 24271 33609
rect 24762 33600 24768 33612
rect 24820 33600 24826 33652
rect 13202 33544 15424 33572
rect 15488 33544 15700 33572
rect 15749 33575 15807 33581
rect 10836 33476 11560 33504
rect 10836 33464 10842 33476
rect 11606 33464 11612 33516
rect 11664 33504 11670 33516
rect 11701 33507 11759 33513
rect 11701 33504 11713 33507
rect 11664 33476 11713 33504
rect 11664 33464 11670 33476
rect 11701 33473 11713 33476
rect 11747 33473 11759 33507
rect 13722 33504 13728 33516
rect 13683 33476 13728 33504
rect 11701 33467 11759 33473
rect 13722 33464 13728 33476
rect 13780 33464 13786 33516
rect 13906 33464 13912 33516
rect 13964 33504 13970 33516
rect 14366 33504 14372 33516
rect 13964 33476 14372 33504
rect 13964 33464 13970 33476
rect 14366 33464 14372 33476
rect 14424 33504 14430 33516
rect 14645 33507 14703 33513
rect 14645 33504 14657 33507
rect 14424 33476 14657 33504
rect 14424 33464 14430 33476
rect 14645 33473 14657 33476
rect 14691 33504 14703 33507
rect 15488 33504 15516 33544
rect 15749 33541 15761 33575
rect 15795 33572 15807 33575
rect 16942 33572 16948 33584
rect 15795 33544 16948 33572
rect 15795 33541 15807 33544
rect 15749 33535 15807 33541
rect 16942 33532 16948 33544
rect 17000 33532 17006 33584
rect 18414 33572 18420 33584
rect 17144 33544 18420 33572
rect 14691 33476 15516 33504
rect 16301 33507 16359 33513
rect 14691 33473 14703 33476
rect 14645 33467 14703 33473
rect 16301 33473 16313 33507
rect 16347 33504 16359 33507
rect 17144 33504 17172 33544
rect 18414 33532 18420 33544
rect 18472 33532 18478 33584
rect 18690 33532 18696 33584
rect 18748 33572 18754 33584
rect 18785 33575 18843 33581
rect 18785 33572 18797 33575
rect 18748 33544 18797 33572
rect 18748 33532 18754 33544
rect 18785 33541 18797 33544
rect 18831 33541 18843 33575
rect 18785 33535 18843 33541
rect 19058 33532 19064 33584
rect 19116 33572 19122 33584
rect 19521 33575 19579 33581
rect 19521 33572 19533 33575
rect 19116 33544 19533 33572
rect 19116 33532 19122 33544
rect 19521 33541 19533 33544
rect 19567 33541 19579 33575
rect 19521 33535 19579 33541
rect 19613 33575 19671 33581
rect 19613 33541 19625 33575
rect 19659 33572 19671 33575
rect 19978 33572 19984 33584
rect 19659 33544 19984 33572
rect 19659 33541 19671 33544
rect 19613 33535 19671 33541
rect 19978 33532 19984 33544
rect 20036 33532 20042 33584
rect 24578 33572 24584 33584
rect 21192 33544 24584 33572
rect 17310 33504 17316 33516
rect 16347 33476 17172 33504
rect 17271 33476 17316 33504
rect 16347 33473 16359 33476
rect 16301 33467 16359 33473
rect 17310 33464 17316 33476
rect 17368 33464 17374 33516
rect 9858 33396 9864 33448
rect 9916 33436 9922 33448
rect 11149 33439 11207 33445
rect 11149 33436 11161 33439
rect 9916 33408 11161 33436
rect 9916 33396 9922 33408
rect 11149 33405 11161 33408
rect 11195 33405 11207 33439
rect 11149 33399 11207 33405
rect 11238 33396 11244 33448
rect 11296 33436 11302 33448
rect 11624 33436 11652 33464
rect 12710 33436 12716 33448
rect 11296 33408 11652 33436
rect 11808 33408 12716 33436
rect 11296 33396 11302 33408
rect 11808 33368 11836 33408
rect 12710 33396 12716 33408
rect 12768 33396 12774 33448
rect 15654 33436 15660 33448
rect 15615 33408 15660 33436
rect 15654 33396 15660 33408
rect 15712 33396 15718 33448
rect 17129 33439 17187 33445
rect 17129 33405 17141 33439
rect 17175 33436 17187 33439
rect 17218 33436 17224 33448
rect 17175 33408 17224 33436
rect 17175 33405 17187 33408
rect 17129 33399 17187 33405
rect 17218 33396 17224 33408
rect 17276 33396 17282 33448
rect 18598 33436 18604 33448
rect 18559 33408 18604 33436
rect 18598 33396 18604 33408
rect 18656 33396 18662 33448
rect 18877 33439 18935 33445
rect 18877 33405 18889 33439
rect 18923 33436 18935 33439
rect 19794 33436 19800 33448
rect 18923 33408 19288 33436
rect 19755 33408 19800 33436
rect 18923 33405 18935 33408
rect 18877 33399 18935 33405
rect 8220 33340 9260 33368
rect 2280 33272 3740 33300
rect 2280 33260 2286 33272
rect 8294 33260 8300 33312
rect 8352 33300 8358 33312
rect 8573 33303 8631 33309
rect 8573 33300 8585 33303
rect 8352 33272 8585 33300
rect 8352 33260 8358 33272
rect 8573 33269 8585 33272
rect 8619 33269 8631 33303
rect 9232 33300 9260 33340
rect 11624 33340 11836 33368
rect 11624 33300 11652 33340
rect 14550 33328 14556 33380
rect 14608 33368 14614 33380
rect 19260 33368 19288 33408
rect 19794 33396 19800 33408
rect 19852 33396 19858 33448
rect 19334 33368 19340 33380
rect 14608 33340 17448 33368
rect 19260 33340 19340 33368
rect 14608 33328 14614 33340
rect 9232 33272 11652 33300
rect 8573 33263 8631 33269
rect 11790 33260 11796 33312
rect 11848 33300 11854 33312
rect 11964 33303 12022 33309
rect 11964 33300 11976 33303
rect 11848 33272 11976 33300
rect 11848 33260 11854 33272
rect 11964 33269 11976 33272
rect 12010 33300 12022 33303
rect 13446 33300 13452 33312
rect 12010 33272 13452 33300
rect 12010 33269 12022 33272
rect 11964 33263 12022 33269
rect 13446 33260 13452 33272
rect 13504 33260 13510 33312
rect 14737 33303 14795 33309
rect 14737 33269 14749 33303
rect 14783 33300 14795 33303
rect 15378 33300 15384 33312
rect 14783 33272 15384 33300
rect 14783 33269 14795 33272
rect 14737 33263 14795 33269
rect 15378 33260 15384 33272
rect 15436 33260 15442 33312
rect 17420 33300 17448 33340
rect 19334 33328 19340 33340
rect 19392 33328 19398 33380
rect 19518 33300 19524 33312
rect 17420 33272 19524 33300
rect 19518 33260 19524 33272
rect 19576 33260 19582 33312
rect 19610 33260 19616 33312
rect 19668 33300 19674 33312
rect 21192 33309 21220 33544
rect 24578 33532 24584 33544
rect 24636 33532 24642 33584
rect 37553 33507 37611 33513
rect 37553 33473 37565 33507
rect 37599 33504 37611 33507
rect 38194 33504 38200 33516
rect 37599 33476 38200 33504
rect 37599 33473 37611 33476
rect 37553 33467 37611 33473
rect 38194 33464 38200 33476
rect 38252 33464 38258 33516
rect 23658 33368 23664 33380
rect 23619 33340 23664 33368
rect 23658 33328 23664 33340
rect 23716 33328 23722 33380
rect 34514 33328 34520 33380
rect 34572 33368 34578 33380
rect 38013 33371 38071 33377
rect 38013 33368 38025 33371
rect 34572 33340 38025 33368
rect 34572 33328 34578 33340
rect 38013 33337 38025 33340
rect 38059 33337 38071 33371
rect 38013 33331 38071 33337
rect 21177 33303 21235 33309
rect 21177 33300 21189 33303
rect 19668 33272 21189 33300
rect 19668 33260 19674 33272
rect 21177 33269 21189 33272
rect 21223 33269 21235 33303
rect 21177 33263 21235 33269
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 1673 33099 1731 33105
rect 1673 33065 1685 33099
rect 1719 33096 1731 33099
rect 1762 33096 1768 33108
rect 1719 33068 1768 33096
rect 1719 33065 1731 33068
rect 1673 33059 1731 33065
rect 1762 33056 1768 33068
rect 1820 33096 1826 33108
rect 7558 33096 7564 33108
rect 1820 33068 7564 33096
rect 1820 33056 1826 33068
rect 7558 33056 7564 33068
rect 7616 33056 7622 33108
rect 8662 33056 8668 33108
rect 8720 33096 8726 33108
rect 9490 33096 9496 33108
rect 8720 33068 9496 33096
rect 8720 33056 8726 33068
rect 9490 33056 9496 33068
rect 9548 33056 9554 33108
rect 9677 33099 9735 33105
rect 9677 33065 9689 33099
rect 9723 33096 9735 33099
rect 9723 33068 12296 33096
rect 9723 33065 9735 33068
rect 9677 33059 9735 33065
rect 8389 33031 8447 33037
rect 8389 32997 8401 33031
rect 8435 33028 8447 33031
rect 10778 33028 10784 33040
rect 8435 33000 10784 33028
rect 8435 32997 8447 33000
rect 8389 32991 8447 32997
rect 10778 32988 10784 33000
rect 10836 32988 10842 33040
rect 12268 33028 12296 33068
rect 12342 33056 12348 33108
rect 12400 33096 12406 33108
rect 12400 33068 13676 33096
rect 12400 33056 12406 33068
rect 13262 33028 13268 33040
rect 12268 33000 13268 33028
rect 13262 32988 13268 33000
rect 13320 32988 13326 33040
rect 3421 32963 3479 32969
rect 3421 32929 3433 32963
rect 3467 32960 3479 32963
rect 3510 32960 3516 32972
rect 3467 32932 3516 32960
rect 3467 32929 3479 32932
rect 3421 32923 3479 32929
rect 3510 32920 3516 32932
rect 3568 32920 3574 32972
rect 9306 32920 9312 32972
rect 9364 32960 9370 32972
rect 10873 32963 10931 32969
rect 10873 32960 10885 32963
rect 9364 32932 10885 32960
rect 9364 32920 9370 32932
rect 10873 32929 10885 32932
rect 10919 32960 10931 32963
rect 11238 32960 11244 32972
rect 10919 32932 11244 32960
rect 10919 32929 10931 32932
rect 10873 32923 10931 32929
rect 11238 32920 11244 32932
rect 11296 32920 11302 32972
rect 11514 32920 11520 32972
rect 11572 32960 11578 32972
rect 11572 32932 13584 32960
rect 11572 32920 11578 32932
rect 4062 32892 4068 32904
rect 4023 32864 4068 32892
rect 4062 32852 4068 32864
rect 4120 32852 4126 32904
rect 4801 32895 4859 32901
rect 4801 32861 4813 32895
rect 4847 32892 4859 32895
rect 4890 32892 4896 32904
rect 4847 32864 4896 32892
rect 4847 32861 4859 32864
rect 4801 32855 4859 32861
rect 4890 32852 4896 32864
rect 4948 32852 4954 32904
rect 5718 32852 5724 32904
rect 5776 32892 5782 32904
rect 5813 32895 5871 32901
rect 5813 32892 5825 32895
rect 5776 32864 5825 32892
rect 5776 32852 5782 32864
rect 5813 32861 5825 32864
rect 5859 32861 5871 32895
rect 5813 32855 5871 32861
rect 7190 32852 7196 32904
rect 7248 32852 7254 32904
rect 7374 32852 7380 32904
rect 7432 32892 7438 32904
rect 8297 32895 8355 32901
rect 8297 32892 8309 32895
rect 7432 32864 8309 32892
rect 7432 32852 7438 32864
rect 8297 32861 8309 32864
rect 8343 32892 8355 32895
rect 8662 32892 8668 32904
rect 8343 32864 8668 32892
rect 8343 32861 8355 32864
rect 8297 32855 8355 32861
rect 8662 32852 8668 32864
rect 8720 32852 8726 32904
rect 9582 32892 9588 32904
rect 9543 32864 9588 32892
rect 9582 32852 9588 32864
rect 9640 32852 9646 32904
rect 10229 32895 10287 32901
rect 10229 32892 10241 32895
rect 9692 32864 10241 32892
rect 2590 32784 2596 32836
rect 2648 32784 2654 32836
rect 3145 32827 3203 32833
rect 3145 32793 3157 32827
rect 3191 32793 3203 32827
rect 4246 32824 4252 32836
rect 4207 32796 4252 32824
rect 3145 32787 3203 32793
rect 3160 32756 3188 32787
rect 4246 32784 4252 32796
rect 4304 32784 4310 32836
rect 6086 32824 6092 32836
rect 6047 32796 6092 32824
rect 6086 32784 6092 32796
rect 6144 32784 6150 32836
rect 7837 32827 7895 32833
rect 7837 32793 7849 32827
rect 7883 32824 7895 32827
rect 8110 32824 8116 32836
rect 7883 32796 8116 32824
rect 7883 32793 7895 32796
rect 7837 32787 7895 32793
rect 8110 32784 8116 32796
rect 8168 32784 8174 32836
rect 9490 32784 9496 32836
rect 9548 32824 9554 32836
rect 9692 32824 9720 32864
rect 10229 32861 10241 32864
rect 10275 32861 10287 32895
rect 12802 32892 12808 32904
rect 12282 32864 12808 32892
rect 10229 32855 10287 32861
rect 12802 32852 12808 32864
rect 12860 32852 12866 32904
rect 13556 32901 13584 32932
rect 13541 32895 13599 32901
rect 13541 32861 13553 32895
rect 13587 32861 13599 32895
rect 13648 32892 13676 33068
rect 15102 33056 15108 33108
rect 15160 33096 15166 33108
rect 18049 33099 18107 33105
rect 18049 33096 18061 33099
rect 15160 33068 18061 33096
rect 15160 33056 15166 33068
rect 18049 33065 18061 33068
rect 18095 33065 18107 33099
rect 18049 33059 18107 33065
rect 18506 33056 18512 33108
rect 18564 33096 18570 33108
rect 18693 33099 18751 33105
rect 18693 33096 18705 33099
rect 18564 33068 18705 33096
rect 18564 33056 18570 33068
rect 18693 33065 18705 33068
rect 18739 33065 18751 33099
rect 19518 33096 19524 33108
rect 19479 33068 19524 33096
rect 18693 33059 18751 33065
rect 19518 33056 19524 33068
rect 19576 33056 19582 33108
rect 20162 33096 20168 33108
rect 20123 33068 20168 33096
rect 20162 33056 20168 33068
rect 20220 33056 20226 33108
rect 22005 33099 22063 33105
rect 22005 33065 22017 33099
rect 22051 33096 22063 33099
rect 22557 33099 22615 33105
rect 22557 33096 22569 33099
rect 22051 33068 22569 33096
rect 22051 33065 22063 33068
rect 22005 33059 22063 33065
rect 22557 33065 22569 33068
rect 22603 33096 22615 33099
rect 22922 33096 22928 33108
rect 22603 33068 22928 33096
rect 22603 33065 22615 33068
rect 22557 33059 22615 33065
rect 22922 33056 22928 33068
rect 22980 33096 22986 33108
rect 23569 33099 23627 33105
rect 23569 33096 23581 33099
rect 22980 33068 23581 33096
rect 22980 33056 22986 33068
rect 23569 33065 23581 33068
rect 23615 33096 23627 33099
rect 24581 33099 24639 33105
rect 24581 33096 24593 33099
rect 23615 33068 24593 33096
rect 23615 33065 23627 33068
rect 23569 33059 23627 33065
rect 24581 33065 24593 33068
rect 24627 33065 24639 33099
rect 24581 33059 24639 33065
rect 13906 32988 13912 33040
rect 13964 33028 13970 33040
rect 15197 33031 15255 33037
rect 15197 33028 15209 33031
rect 13964 33000 15209 33028
rect 13964 32988 13970 33000
rect 15197 32997 15209 33000
rect 15243 32997 15255 33031
rect 15930 33028 15936 33040
rect 15843 33000 15936 33028
rect 15197 32991 15255 32997
rect 15930 32988 15936 33000
rect 15988 33028 15994 33040
rect 17678 33028 17684 33040
rect 15988 33000 17684 33028
rect 15988 32988 15994 33000
rect 17678 32988 17684 33000
rect 17736 32988 17742 33040
rect 18138 32988 18144 33040
rect 18196 33028 18202 33040
rect 19150 33028 19156 33040
rect 18196 33000 19156 33028
rect 18196 32988 18202 33000
rect 19150 32988 19156 33000
rect 19208 33028 19214 33040
rect 20898 33028 20904 33040
rect 19208 33000 20904 33028
rect 19208 32988 19214 33000
rect 20898 32988 20904 33000
rect 20956 32988 20962 33040
rect 13722 32920 13728 32972
rect 13780 32960 13786 32972
rect 14826 32960 14832 32972
rect 13780 32932 14832 32960
rect 13780 32920 13786 32932
rect 14826 32920 14832 32932
rect 14884 32920 14890 32972
rect 16206 32920 16212 32972
rect 16264 32960 16270 32972
rect 16482 32960 16488 32972
rect 16264 32932 16488 32960
rect 16264 32920 16270 32932
rect 16482 32920 16488 32932
rect 16540 32920 16546 32972
rect 17310 32920 17316 32972
rect 17368 32960 17374 32972
rect 21818 32960 21824 32972
rect 17368 32932 21824 32960
rect 17368 32920 17374 32932
rect 21818 32920 21824 32932
rect 21876 32920 21882 32972
rect 14461 32895 14519 32901
rect 14461 32892 14473 32895
rect 13648 32864 14473 32892
rect 13541 32855 13599 32861
rect 14461 32861 14473 32864
rect 14507 32861 14519 32895
rect 14461 32855 14519 32861
rect 15194 32852 15200 32904
rect 15252 32892 15258 32904
rect 15289 32895 15347 32901
rect 15289 32892 15301 32895
rect 15252 32864 15301 32892
rect 15252 32852 15258 32864
rect 15289 32861 15301 32864
rect 15335 32861 15347 32895
rect 17034 32892 17040 32904
rect 16995 32864 17040 32892
rect 15289 32855 15347 32861
rect 17034 32852 17040 32864
rect 17092 32852 17098 32904
rect 17218 32852 17224 32904
rect 17276 32892 17282 32904
rect 18138 32892 18144 32904
rect 17276 32864 18144 32892
rect 17276 32852 17282 32864
rect 18138 32852 18144 32864
rect 18196 32852 18202 32904
rect 18230 32852 18236 32904
rect 18288 32892 18294 32904
rect 18785 32895 18843 32901
rect 18785 32892 18797 32895
rect 18288 32864 18797 32892
rect 18288 32852 18294 32864
rect 18785 32861 18797 32864
rect 18831 32892 18843 32895
rect 19242 32892 19248 32904
rect 18831 32864 19248 32892
rect 18831 32861 18843 32864
rect 18785 32855 18843 32861
rect 19242 32852 19248 32864
rect 19300 32852 19306 32904
rect 19613 32895 19671 32901
rect 19613 32861 19625 32895
rect 19659 32892 19671 32895
rect 20257 32895 20315 32901
rect 20257 32892 20269 32895
rect 19659 32864 20269 32892
rect 19659 32861 19671 32864
rect 19613 32855 19671 32861
rect 20257 32861 20269 32864
rect 20303 32861 20315 32895
rect 20257 32855 20315 32861
rect 9548 32796 9720 32824
rect 9548 32784 9554 32796
rect 10042 32784 10048 32836
rect 10100 32824 10106 32836
rect 11149 32827 11207 32833
rect 11149 32824 11161 32827
rect 10100 32796 11161 32824
rect 10100 32784 10106 32796
rect 11149 32793 11161 32796
rect 11195 32793 11207 32827
rect 11149 32787 11207 32793
rect 12434 32784 12440 32836
rect 12492 32824 12498 32836
rect 12897 32827 12955 32833
rect 12897 32824 12909 32827
rect 12492 32796 12909 32824
rect 12492 32784 12498 32796
rect 12897 32793 12909 32796
rect 12943 32824 12955 32827
rect 13078 32824 13084 32836
rect 12943 32796 13084 32824
rect 12943 32793 12955 32796
rect 12897 32787 12955 32793
rect 13078 32784 13084 32796
rect 13136 32784 13142 32836
rect 16393 32827 16451 32833
rect 16393 32793 16405 32827
rect 16439 32824 16451 32827
rect 17126 32824 17132 32836
rect 16439 32796 17132 32824
rect 16439 32793 16451 32796
rect 16393 32787 16451 32793
rect 17126 32784 17132 32796
rect 17184 32784 17190 32836
rect 17310 32824 17316 32836
rect 17271 32796 17316 32824
rect 17310 32784 17316 32796
rect 17368 32784 17374 32836
rect 18046 32784 18052 32836
rect 18104 32824 18110 32836
rect 19150 32824 19156 32836
rect 18104 32796 19156 32824
rect 18104 32784 18110 32796
rect 19150 32784 19156 32796
rect 19208 32824 19214 32836
rect 19628 32824 19656 32855
rect 20714 32852 20720 32904
rect 20772 32892 20778 32904
rect 20901 32895 20959 32901
rect 20901 32892 20913 32895
rect 20772 32864 20913 32892
rect 20772 32852 20778 32864
rect 20901 32861 20913 32864
rect 20947 32892 20959 32895
rect 20990 32892 20996 32904
rect 20947 32864 20996 32892
rect 20947 32861 20959 32864
rect 20901 32855 20959 32861
rect 20990 32852 20996 32864
rect 21048 32892 21054 32904
rect 21361 32895 21419 32901
rect 21361 32892 21373 32895
rect 21048 32864 21373 32892
rect 21048 32852 21054 32864
rect 21361 32861 21373 32864
rect 21407 32861 21419 32895
rect 21361 32855 21419 32861
rect 19208 32796 19656 32824
rect 20809 32827 20867 32833
rect 19208 32784 19214 32796
rect 20809 32793 20821 32827
rect 20855 32824 20867 32827
rect 21082 32824 21088 32836
rect 20855 32796 21088 32824
rect 20855 32793 20867 32796
rect 20809 32787 20867 32793
rect 21082 32784 21088 32796
rect 21140 32784 21146 32836
rect 4706 32756 4712 32768
rect 3160 32728 4712 32756
rect 4706 32716 4712 32728
rect 4764 32716 4770 32768
rect 4893 32759 4951 32765
rect 4893 32725 4905 32759
rect 4939 32756 4951 32759
rect 9950 32756 9956 32768
rect 4939 32728 9956 32756
rect 4939 32725 4951 32728
rect 4893 32719 4951 32725
rect 9950 32716 9956 32728
rect 10008 32716 10014 32768
rect 10321 32759 10379 32765
rect 10321 32725 10333 32759
rect 10367 32756 10379 32759
rect 11790 32756 11796 32768
rect 10367 32728 11796 32756
rect 10367 32725 10379 32728
rect 10321 32719 10379 32725
rect 11790 32716 11796 32728
rect 11848 32716 11854 32768
rect 11882 32716 11888 32768
rect 11940 32756 11946 32768
rect 13446 32756 13452 32768
rect 11940 32728 13452 32756
rect 11940 32716 11946 32728
rect 13446 32716 13452 32728
rect 13504 32716 13510 32768
rect 13630 32756 13636 32768
rect 13591 32728 13636 32756
rect 13630 32716 13636 32728
rect 13688 32716 13694 32768
rect 14553 32759 14611 32765
rect 14553 32725 14565 32759
rect 14599 32756 14611 32759
rect 14826 32756 14832 32768
rect 14599 32728 14832 32756
rect 14599 32725 14611 32728
rect 14553 32719 14611 32725
rect 14826 32716 14832 32728
rect 14884 32716 14890 32768
rect 17494 32716 17500 32768
rect 17552 32756 17558 32768
rect 19794 32756 19800 32768
rect 17552 32728 19800 32756
rect 17552 32716 17558 32728
rect 19794 32716 19800 32728
rect 19852 32716 19858 32768
rect 23109 32759 23167 32765
rect 23109 32725 23121 32759
rect 23155 32756 23167 32759
rect 23290 32756 23296 32768
rect 23155 32728 23296 32756
rect 23155 32725 23167 32728
rect 23109 32719 23167 32725
rect 23290 32716 23296 32728
rect 23348 32716 23354 32768
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 7282 32512 7288 32564
rect 7340 32552 7346 32564
rect 9490 32552 9496 32564
rect 7340 32524 9496 32552
rect 7340 32512 7346 32524
rect 9490 32512 9496 32524
rect 9548 32512 9554 32564
rect 9582 32512 9588 32564
rect 9640 32552 9646 32564
rect 11146 32552 11152 32564
rect 9640 32524 11152 32552
rect 9640 32512 9646 32524
rect 11146 32512 11152 32524
rect 11204 32512 11210 32564
rect 13630 32512 13636 32564
rect 13688 32552 13694 32564
rect 21085 32555 21143 32561
rect 13688 32524 17908 32552
rect 13688 32512 13694 32524
rect 2682 32444 2688 32496
rect 2740 32444 2746 32496
rect 5902 32484 5908 32496
rect 5474 32456 5908 32484
rect 5902 32444 5908 32456
rect 5960 32444 5966 32496
rect 5994 32444 6000 32496
rect 6052 32484 6058 32496
rect 6052 32456 6097 32484
rect 6052 32444 6058 32456
rect 6546 32444 6552 32496
rect 6604 32484 6610 32496
rect 6604 32456 6684 32484
rect 6604 32444 6610 32456
rect 3510 32376 3516 32428
rect 3568 32416 3574 32428
rect 3786 32416 3792 32428
rect 3568 32388 3792 32416
rect 3568 32376 3574 32388
rect 3786 32376 3792 32388
rect 3844 32416 3850 32428
rect 3973 32419 4031 32425
rect 3973 32416 3985 32419
rect 3844 32388 3985 32416
rect 3844 32376 3850 32388
rect 3973 32385 3985 32388
rect 4019 32385 4031 32419
rect 3973 32379 4031 32385
rect 3237 32351 3295 32357
rect 3237 32317 3249 32351
rect 3283 32348 3295 32351
rect 4249 32351 4307 32357
rect 3283 32320 4108 32348
rect 3283 32317 3295 32320
rect 3237 32311 3295 32317
rect 1762 32212 1768 32224
rect 1723 32184 1768 32212
rect 1762 32172 1768 32184
rect 1820 32172 1826 32224
rect 4080 32212 4108 32320
rect 4249 32317 4261 32351
rect 4295 32348 4307 32351
rect 4798 32348 4804 32360
rect 4295 32320 4804 32348
rect 4295 32317 4307 32320
rect 4249 32311 4307 32317
rect 4798 32308 4804 32320
rect 4856 32308 4862 32360
rect 6546 32348 6552 32360
rect 6507 32320 6552 32348
rect 6546 32308 6552 32320
rect 6604 32308 6610 32360
rect 6656 32348 6684 32456
rect 7006 32444 7012 32496
rect 7064 32484 7070 32496
rect 8297 32487 8355 32493
rect 7064 32456 7130 32484
rect 7064 32444 7070 32456
rect 8297 32453 8309 32487
rect 8343 32484 8355 32487
rect 9674 32484 9680 32496
rect 8343 32456 9680 32484
rect 8343 32453 8355 32456
rect 8297 32447 8355 32453
rect 9674 32444 9680 32456
rect 9732 32444 9738 32496
rect 11514 32484 11520 32496
rect 10810 32456 11520 32484
rect 11514 32444 11520 32456
rect 11572 32444 11578 32496
rect 12618 32444 12624 32496
rect 12676 32444 12682 32496
rect 13170 32484 13176 32496
rect 13131 32456 13176 32484
rect 13170 32444 13176 32456
rect 13228 32444 13234 32496
rect 14090 32484 14096 32496
rect 14051 32456 14096 32484
rect 14090 32444 14096 32456
rect 14148 32444 14154 32496
rect 15470 32484 15476 32496
rect 15431 32456 15476 32484
rect 15470 32444 15476 32456
rect 15528 32444 15534 32496
rect 17880 32493 17908 32524
rect 21085 32521 21097 32555
rect 21131 32552 21143 32555
rect 21634 32552 21640 32564
rect 21131 32524 21640 32552
rect 21131 32521 21143 32524
rect 21085 32515 21143 32521
rect 21634 32512 21640 32524
rect 21692 32512 21698 32564
rect 22649 32555 22707 32561
rect 22649 32521 22661 32555
rect 22695 32552 22707 32555
rect 22922 32552 22928 32564
rect 22695 32524 22928 32552
rect 22695 32521 22707 32524
rect 22649 32515 22707 32521
rect 22922 32512 22928 32524
rect 22980 32552 22986 32564
rect 23109 32555 23167 32561
rect 23109 32552 23121 32555
rect 22980 32524 23121 32552
rect 22980 32512 22986 32524
rect 23109 32521 23121 32524
rect 23155 32552 23167 32555
rect 23661 32555 23719 32561
rect 23661 32552 23673 32555
rect 23155 32524 23673 32552
rect 23155 32521 23167 32524
rect 23109 32515 23167 32521
rect 23661 32521 23673 32524
rect 23707 32521 23719 32555
rect 23661 32515 23719 32521
rect 17865 32487 17923 32493
rect 17865 32453 17877 32487
rect 17911 32453 17923 32487
rect 18414 32484 18420 32496
rect 18375 32456 18420 32484
rect 17865 32447 17923 32453
rect 18414 32444 18420 32456
rect 18472 32444 18478 32496
rect 19242 32444 19248 32496
rect 19300 32484 19306 32496
rect 20714 32484 20720 32496
rect 19300 32456 20720 32484
rect 19300 32444 19306 32456
rect 20714 32444 20720 32456
rect 20772 32444 20778 32496
rect 8573 32419 8631 32425
rect 8573 32385 8585 32419
rect 8619 32416 8631 32419
rect 9306 32416 9312 32428
rect 8619 32388 9312 32416
rect 8619 32385 8631 32388
rect 8573 32379 8631 32385
rect 9306 32376 9312 32388
rect 9364 32376 9370 32428
rect 14642 32376 14648 32428
rect 14700 32416 14706 32428
rect 17037 32419 17095 32425
rect 17037 32416 17049 32419
rect 14700 32388 14745 32416
rect 16960 32388 17049 32416
rect 14700 32376 14706 32388
rect 6656 32320 8524 32348
rect 8496 32280 8524 32320
rect 9122 32308 9128 32360
rect 9180 32348 9186 32360
rect 9582 32348 9588 32360
rect 9180 32320 9588 32348
rect 9180 32308 9186 32320
rect 9582 32308 9588 32320
rect 9640 32308 9646 32360
rect 11238 32308 11244 32360
rect 11296 32348 11302 32360
rect 13449 32351 13507 32357
rect 13449 32348 13461 32351
rect 11296 32320 13461 32348
rect 11296 32308 11302 32320
rect 13449 32317 13461 32320
rect 13495 32348 13507 32351
rect 13722 32348 13728 32360
rect 13495 32320 13728 32348
rect 13495 32317 13507 32320
rect 13449 32311 13507 32317
rect 13722 32308 13728 32320
rect 13780 32308 13786 32360
rect 14001 32351 14059 32357
rect 14001 32317 14013 32351
rect 14047 32317 14059 32351
rect 14001 32311 14059 32317
rect 15381 32351 15439 32357
rect 15381 32317 15393 32351
rect 15427 32348 15439 32351
rect 15470 32348 15476 32360
rect 15427 32320 15476 32348
rect 15427 32317 15439 32320
rect 15381 32311 15439 32317
rect 9306 32280 9312 32292
rect 8496 32252 9312 32280
rect 9306 32240 9312 32252
rect 9364 32240 9370 32292
rect 11057 32283 11115 32289
rect 11057 32249 11069 32283
rect 11103 32280 11115 32283
rect 11882 32280 11888 32292
rect 11103 32252 11888 32280
rect 11103 32249 11115 32252
rect 11057 32243 11115 32249
rect 11882 32240 11888 32252
rect 11940 32240 11946 32292
rect 13538 32240 13544 32292
rect 13596 32280 13602 32292
rect 14016 32280 14044 32311
rect 15470 32308 15476 32320
rect 15528 32308 15534 32360
rect 16666 32308 16672 32360
rect 16724 32348 16730 32360
rect 16960 32348 16988 32388
rect 17037 32385 17049 32388
rect 17083 32385 17095 32419
rect 17037 32379 17095 32385
rect 17402 32376 17408 32428
rect 17460 32376 17466 32428
rect 19150 32376 19156 32428
rect 19208 32416 19214 32428
rect 19889 32419 19947 32425
rect 19889 32416 19901 32419
rect 19208 32388 19901 32416
rect 19208 32376 19214 32388
rect 19889 32385 19901 32388
rect 19935 32416 19947 32419
rect 20349 32419 20407 32425
rect 20349 32416 20361 32419
rect 19935 32388 20361 32416
rect 19935 32385 19947 32388
rect 19889 32379 19947 32385
rect 20349 32385 20361 32388
rect 20395 32385 20407 32419
rect 20349 32379 20407 32385
rect 20898 32376 20904 32428
rect 20956 32416 20962 32428
rect 20993 32419 21051 32425
rect 20993 32416 21005 32419
rect 20956 32388 21005 32416
rect 20956 32376 20962 32388
rect 20993 32385 21005 32388
rect 21039 32385 21051 32419
rect 20993 32379 21051 32385
rect 37553 32419 37611 32425
rect 37553 32385 37565 32419
rect 37599 32416 37611 32419
rect 38194 32416 38200 32428
rect 37599 32388 38200 32416
rect 37599 32385 37611 32388
rect 37553 32379 37611 32385
rect 38194 32376 38200 32388
rect 38252 32376 38258 32428
rect 16724 32320 16988 32348
rect 16724 32308 16730 32320
rect 13596 32252 14044 32280
rect 15933 32283 15991 32289
rect 13596 32240 13602 32252
rect 15933 32249 15945 32283
rect 15979 32280 15991 32283
rect 16298 32280 16304 32292
rect 15979 32252 16304 32280
rect 15979 32249 15991 32252
rect 15933 32243 15991 32249
rect 16298 32240 16304 32252
rect 16356 32280 16362 32292
rect 17420 32280 17448 32376
rect 17773 32351 17831 32357
rect 17773 32317 17785 32351
rect 17819 32348 17831 32351
rect 19245 32351 19303 32357
rect 17819 32320 19196 32348
rect 17819 32317 17831 32320
rect 17773 32311 17831 32317
rect 16356 32252 17448 32280
rect 19168 32280 19196 32320
rect 19245 32317 19257 32351
rect 19291 32348 19303 32351
rect 20070 32348 20076 32360
rect 19291 32320 20076 32348
rect 19291 32317 19303 32320
rect 19245 32311 19303 32317
rect 20070 32308 20076 32320
rect 20128 32308 20134 32360
rect 22097 32283 22155 32289
rect 22097 32280 22109 32283
rect 19168 32252 22109 32280
rect 16356 32240 16362 32252
rect 22097 32249 22109 32252
rect 22143 32280 22155 32283
rect 23566 32280 23572 32292
rect 22143 32252 23572 32280
rect 22143 32249 22155 32252
rect 22097 32243 22155 32249
rect 23566 32240 23572 32252
rect 23624 32240 23630 32292
rect 38010 32280 38016 32292
rect 37971 32252 38016 32280
rect 38010 32240 38016 32252
rect 38068 32240 38074 32292
rect 7282 32212 7288 32224
rect 4080 32184 7288 32212
rect 7282 32172 7288 32184
rect 7340 32172 7346 32224
rect 8662 32172 8668 32224
rect 8720 32212 8726 32224
rect 10962 32212 10968 32224
rect 8720 32184 10968 32212
rect 8720 32172 8726 32184
rect 10962 32172 10968 32184
rect 11020 32172 11026 32224
rect 11146 32172 11152 32224
rect 11204 32212 11210 32224
rect 11701 32215 11759 32221
rect 11701 32212 11713 32215
rect 11204 32184 11713 32212
rect 11204 32172 11210 32184
rect 11701 32181 11713 32184
rect 11747 32181 11759 32215
rect 11701 32175 11759 32181
rect 12618 32172 12624 32224
rect 12676 32212 12682 32224
rect 12986 32212 12992 32224
rect 12676 32184 12992 32212
rect 12676 32172 12682 32184
rect 12986 32172 12992 32184
rect 13044 32212 13050 32224
rect 16942 32212 16948 32224
rect 13044 32184 16948 32212
rect 13044 32172 13050 32184
rect 16942 32172 16948 32184
rect 17000 32172 17006 32224
rect 17129 32215 17187 32221
rect 17129 32181 17141 32215
rect 17175 32212 17187 32215
rect 17310 32212 17316 32224
rect 17175 32184 17316 32212
rect 17175 32181 17187 32184
rect 17129 32175 17187 32181
rect 17310 32172 17316 32184
rect 17368 32172 17374 32224
rect 17402 32172 17408 32224
rect 17460 32212 17466 32224
rect 19797 32215 19855 32221
rect 19797 32212 19809 32215
rect 17460 32184 19809 32212
rect 17460 32172 17466 32184
rect 19797 32181 19809 32184
rect 19843 32181 19855 32215
rect 19797 32175 19855 32181
rect 20162 32172 20168 32224
rect 20220 32212 20226 32224
rect 20441 32215 20499 32221
rect 20441 32212 20453 32215
rect 20220 32184 20453 32212
rect 20220 32172 20226 32184
rect 20441 32181 20453 32184
rect 20487 32181 20499 32215
rect 20441 32175 20499 32181
rect 22462 32172 22468 32224
rect 22520 32212 22526 32224
rect 24213 32215 24271 32221
rect 24213 32212 24225 32215
rect 22520 32184 24225 32212
rect 22520 32172 22526 32184
rect 24213 32181 24225 32184
rect 24259 32181 24271 32215
rect 24213 32175 24271 32181
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 7558 31968 7564 32020
rect 7616 32008 7622 32020
rect 7616 31980 13492 32008
rect 7616 31968 7622 31980
rect 6730 31940 6736 31952
rect 5644 31912 6736 31940
rect 2593 31875 2651 31881
rect 2593 31841 2605 31875
rect 2639 31872 2651 31875
rect 3050 31872 3056 31884
rect 2639 31844 3056 31872
rect 2639 31841 2651 31844
rect 2593 31835 2651 31841
rect 3050 31832 3056 31844
rect 3108 31832 3114 31884
rect 3602 31832 3608 31884
rect 3660 31872 3666 31884
rect 3973 31875 4031 31881
rect 3973 31872 3985 31875
rect 3660 31844 3985 31872
rect 3660 31832 3666 31844
rect 3973 31841 3985 31844
rect 4019 31841 4031 31875
rect 3973 31835 4031 31841
rect 4890 31832 4896 31884
rect 4948 31872 4954 31884
rect 5074 31872 5080 31884
rect 4948 31844 5080 31872
rect 4948 31832 4954 31844
rect 5074 31832 5080 31844
rect 5132 31832 5138 31884
rect 5445 31875 5503 31881
rect 5445 31841 5457 31875
rect 5491 31872 5503 31875
rect 5644 31872 5672 31912
rect 6730 31900 6736 31912
rect 6788 31900 6794 31952
rect 9490 31940 9496 31952
rect 9451 31912 9496 31940
rect 9490 31900 9496 31912
rect 9548 31900 9554 31952
rect 11422 31900 11428 31952
rect 11480 31940 11486 31952
rect 12989 31943 13047 31949
rect 12989 31940 13001 31943
rect 11480 31912 13001 31940
rect 11480 31900 11486 31912
rect 12989 31909 13001 31912
rect 13035 31909 13047 31943
rect 12989 31903 13047 31909
rect 5491 31844 5672 31872
rect 5736 31844 8524 31872
rect 5491 31841 5503 31844
rect 5445 31835 5503 31841
rect 5736 31816 5764 31844
rect 2774 31764 2780 31816
rect 2832 31804 2838 31816
rect 2869 31807 2927 31813
rect 2869 31804 2881 31807
rect 2832 31776 2881 31804
rect 2832 31764 2838 31776
rect 2869 31773 2881 31776
rect 2915 31804 2927 31807
rect 3142 31804 3148 31816
rect 2915 31776 3148 31804
rect 2915 31773 2927 31776
rect 2869 31767 2927 31773
rect 3142 31764 3148 31776
rect 3200 31764 3206 31816
rect 3418 31804 3424 31816
rect 3379 31776 3424 31804
rect 3418 31764 3424 31776
rect 3476 31764 3482 31816
rect 5718 31764 5724 31816
rect 5776 31804 5782 31816
rect 8496 31813 8524 31844
rect 9674 31832 9680 31884
rect 9732 31872 9738 31884
rect 10962 31872 10968 31884
rect 9732 31844 10968 31872
rect 9732 31832 9738 31844
rect 10962 31832 10968 31844
rect 11020 31832 11026 31884
rect 11238 31872 11244 31884
rect 11199 31844 11244 31872
rect 11238 31832 11244 31844
rect 11296 31832 11302 31884
rect 11790 31832 11796 31884
rect 11848 31872 11854 31884
rect 13354 31872 13360 31884
rect 11848 31844 13360 31872
rect 11848 31832 11854 31844
rect 13354 31832 13360 31844
rect 13412 31832 13418 31884
rect 8481 31807 8539 31813
rect 5776 31776 5821 31804
rect 5776 31764 5782 31776
rect 8481 31773 8493 31807
rect 8527 31804 8539 31807
rect 8662 31804 8668 31816
rect 8527 31776 8668 31804
rect 8527 31773 8539 31776
rect 8481 31767 8539 31773
rect 8662 31764 8668 31776
rect 8720 31764 8726 31816
rect 8772 31776 9674 31804
rect 4890 31696 4896 31748
rect 4948 31696 4954 31748
rect 5442 31696 5448 31748
rect 5500 31736 5506 31748
rect 5902 31736 5908 31748
rect 5500 31708 5908 31736
rect 5500 31696 5506 31708
rect 5902 31696 5908 31708
rect 5960 31696 5966 31748
rect 6362 31696 6368 31748
rect 6420 31736 6426 31748
rect 6457 31739 6515 31745
rect 6457 31736 6469 31739
rect 6420 31708 6469 31736
rect 6420 31696 6426 31708
rect 6457 31705 6469 31708
rect 6503 31705 6515 31739
rect 6457 31699 6515 31705
rect 6914 31696 6920 31748
rect 6972 31736 6978 31748
rect 6972 31708 7038 31736
rect 6972 31696 6978 31708
rect 8110 31696 8116 31748
rect 8168 31736 8174 31748
rect 8205 31739 8263 31745
rect 8205 31736 8217 31739
rect 8168 31708 8217 31736
rect 8168 31696 8174 31708
rect 8205 31705 8217 31708
rect 8251 31736 8263 31739
rect 8772 31736 8800 31776
rect 8251 31708 8800 31736
rect 8251 31705 8263 31708
rect 8205 31699 8263 31705
rect 4798 31628 4804 31680
rect 4856 31668 4862 31680
rect 7926 31668 7932 31680
rect 4856 31640 7932 31668
rect 4856 31628 4862 31640
rect 7926 31628 7932 31640
rect 7984 31628 7990 31680
rect 9646 31668 9674 31776
rect 9858 31764 9864 31816
rect 9916 31764 9922 31816
rect 11330 31764 11336 31816
rect 11388 31804 11394 31816
rect 12253 31807 12311 31813
rect 12253 31804 12265 31807
rect 11388 31776 12265 31804
rect 11388 31764 11394 31776
rect 12253 31773 12265 31776
rect 12299 31773 12311 31807
rect 13078 31804 13084 31816
rect 13039 31776 13084 31804
rect 12253 31767 12311 31773
rect 13078 31764 13084 31776
rect 13136 31764 13142 31816
rect 13464 31804 13492 31980
rect 13630 31968 13636 32020
rect 13688 32008 13694 32020
rect 16853 32011 16911 32017
rect 16853 32008 16865 32011
rect 13688 31980 16865 32008
rect 13688 31968 13694 31980
rect 16853 31977 16865 31980
rect 16899 31977 16911 32011
rect 16853 31971 16911 31977
rect 16942 31968 16948 32020
rect 17000 32008 17006 32020
rect 22465 32011 22523 32017
rect 17000 31980 22094 32008
rect 17000 31968 17006 31980
rect 15286 31900 15292 31952
rect 15344 31940 15350 31952
rect 15841 31943 15899 31949
rect 15344 31912 15792 31940
rect 15344 31900 15350 31912
rect 13633 31875 13691 31881
rect 13633 31841 13645 31875
rect 13679 31872 13691 31875
rect 15470 31872 15476 31884
rect 13679 31844 15476 31872
rect 13679 31841 13691 31844
rect 13633 31835 13691 31841
rect 15470 31832 15476 31844
rect 15528 31832 15534 31884
rect 15764 31872 15792 31912
rect 15841 31909 15853 31943
rect 15887 31940 15899 31943
rect 16298 31940 16304 31952
rect 15887 31912 16304 31940
rect 15887 31909 15899 31912
rect 15841 31903 15899 31909
rect 16298 31900 16304 31912
rect 16356 31900 16362 31952
rect 16390 31900 16396 31952
rect 16448 31940 16454 31952
rect 20714 31940 20720 31952
rect 16448 31912 20208 31940
rect 20675 31912 20720 31940
rect 16448 31900 16454 31912
rect 15764 31844 15976 31872
rect 13541 31817 13599 31823
rect 13541 31804 13553 31817
rect 13464 31783 13553 31804
rect 13587 31783 13599 31817
rect 13464 31777 13599 31783
rect 13464 31776 13584 31777
rect 14090 31764 14096 31816
rect 14148 31804 14154 31816
rect 14737 31807 14795 31813
rect 14737 31804 14749 31807
rect 14148 31776 14749 31804
rect 14148 31764 14154 31776
rect 14737 31773 14749 31776
rect 14783 31804 14795 31807
rect 15102 31804 15108 31816
rect 14783 31776 15108 31804
rect 14783 31773 14795 31776
rect 14737 31767 14795 31773
rect 15102 31764 15108 31776
rect 15160 31764 15166 31816
rect 10965 31739 11023 31745
rect 10965 31705 10977 31739
rect 11011 31736 11023 31739
rect 12158 31736 12164 31748
rect 11011 31708 12164 31736
rect 11011 31705 11023 31708
rect 10965 31699 11023 31705
rect 12158 31696 12164 31708
rect 12216 31696 12222 31748
rect 13170 31696 13176 31748
rect 13228 31736 13234 31748
rect 13538 31736 13544 31748
rect 13228 31708 13544 31736
rect 13228 31696 13234 31708
rect 13538 31696 13544 31708
rect 13596 31696 13602 31748
rect 14642 31736 14648 31748
rect 14603 31708 14648 31736
rect 14642 31696 14648 31708
rect 14700 31696 14706 31748
rect 15286 31736 15292 31748
rect 15248 31708 15292 31736
rect 15286 31696 15292 31708
rect 15344 31696 15350 31748
rect 15381 31739 15439 31745
rect 15381 31705 15393 31739
rect 15427 31736 15439 31739
rect 15948 31736 15976 31844
rect 16114 31832 16120 31884
rect 16172 31872 16178 31884
rect 17497 31875 17555 31881
rect 17497 31872 17509 31875
rect 16172 31844 17509 31872
rect 16172 31832 16178 31844
rect 17497 31841 17509 31844
rect 17543 31841 17555 31875
rect 17497 31835 17555 31841
rect 17678 31832 17684 31884
rect 17736 31872 17742 31884
rect 19429 31875 19487 31881
rect 19429 31872 19441 31875
rect 17736 31844 19441 31872
rect 17736 31832 17742 31844
rect 19429 31841 19441 31844
rect 19475 31841 19487 31875
rect 20070 31872 20076 31884
rect 20031 31844 20076 31872
rect 19429 31835 19487 31841
rect 20070 31832 20076 31844
rect 20128 31832 20134 31884
rect 20180 31872 20208 31912
rect 20714 31900 20720 31912
rect 20772 31900 20778 31952
rect 22066 31940 22094 31980
rect 22465 31977 22477 32011
rect 22511 32008 22523 32011
rect 22922 32008 22928 32020
rect 22511 31980 22928 32008
rect 22511 31977 22523 31980
rect 22465 31971 22523 31977
rect 22922 31968 22928 31980
rect 22980 31968 22986 32020
rect 23477 31943 23535 31949
rect 23477 31940 23489 31943
rect 22066 31912 23489 31940
rect 23477 31909 23489 31912
rect 23523 31909 23535 31943
rect 23477 31903 23535 31909
rect 22925 31875 22983 31881
rect 22925 31872 22937 31875
rect 20180 31844 22937 31872
rect 22925 31841 22937 31844
rect 22971 31841 22983 31875
rect 22925 31835 22983 31841
rect 16666 31764 16672 31816
rect 16724 31804 16730 31816
rect 16945 31807 17003 31813
rect 16945 31804 16957 31807
rect 16724 31776 16957 31804
rect 16724 31764 16730 31776
rect 16945 31773 16957 31776
rect 16991 31804 17003 31807
rect 17218 31804 17224 31816
rect 16991 31776 17224 31804
rect 16991 31773 17003 31776
rect 16945 31767 17003 31773
rect 17218 31764 17224 31776
rect 17276 31764 17282 31816
rect 20809 31807 20867 31813
rect 20809 31773 20821 31807
rect 20855 31804 20867 31807
rect 20990 31804 20996 31816
rect 20855 31776 20996 31804
rect 20855 31773 20867 31776
rect 20809 31767 20867 31773
rect 20990 31764 20996 31776
rect 21048 31804 21054 31816
rect 21266 31804 21272 31816
rect 21048 31776 21272 31804
rect 21048 31764 21054 31776
rect 21266 31764 21272 31776
rect 21324 31804 21330 31816
rect 21821 31807 21879 31813
rect 21821 31804 21833 31807
rect 21324 31776 21833 31804
rect 21324 31764 21330 31776
rect 21821 31773 21833 31776
rect 21867 31773 21879 31807
rect 21821 31767 21879 31773
rect 17586 31736 17592 31748
rect 15427 31708 15976 31736
rect 17547 31708 17592 31736
rect 15427 31705 15439 31708
rect 15381 31699 15439 31705
rect 17586 31696 17592 31708
rect 17644 31696 17650 31748
rect 17862 31696 17868 31748
rect 17920 31736 17926 31748
rect 18509 31739 18567 31745
rect 18509 31736 18521 31739
rect 17920 31708 18521 31736
rect 17920 31696 17926 31708
rect 18509 31705 18521 31708
rect 18555 31736 18567 31739
rect 18874 31736 18880 31748
rect 18555 31708 18880 31736
rect 18555 31705 18567 31708
rect 18509 31699 18567 31705
rect 18874 31696 18880 31708
rect 18932 31696 18938 31748
rect 19978 31736 19984 31748
rect 19939 31708 19984 31736
rect 19978 31696 19984 31708
rect 20036 31696 20042 31748
rect 11793 31671 11851 31677
rect 11793 31668 11805 31671
rect 9646 31640 11805 31668
rect 11793 31637 11805 31640
rect 11839 31668 11851 31671
rect 12250 31668 12256 31680
rect 11839 31640 12256 31668
rect 11839 31637 11851 31640
rect 11793 31631 11851 31637
rect 12250 31628 12256 31640
rect 12308 31628 12314 31680
rect 12345 31671 12403 31677
rect 12345 31637 12357 31671
rect 12391 31668 12403 31671
rect 13446 31668 13452 31680
rect 12391 31640 13452 31668
rect 12391 31637 12403 31640
rect 12345 31631 12403 31637
rect 13446 31628 13452 31640
rect 13504 31628 13510 31680
rect 13556 31668 13584 31696
rect 14918 31668 14924 31680
rect 13556 31640 14924 31668
rect 14918 31628 14924 31640
rect 14976 31628 14982 31680
rect 15562 31628 15568 31680
rect 15620 31668 15626 31680
rect 20990 31668 20996 31680
rect 15620 31640 20996 31668
rect 15620 31628 15626 31640
rect 20990 31628 20996 31640
rect 21048 31628 21054 31680
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 1670 31464 1676 31476
rect 1631 31436 1676 31464
rect 1670 31424 1676 31436
rect 1728 31424 1734 31476
rect 3421 31467 3479 31473
rect 3421 31433 3433 31467
rect 3467 31464 3479 31467
rect 7098 31464 7104 31476
rect 3467 31436 7104 31464
rect 3467 31433 3479 31436
rect 3421 31427 3479 31433
rect 7098 31424 7104 31436
rect 7156 31424 7162 31476
rect 9122 31424 9128 31476
rect 9180 31464 9186 31476
rect 10134 31464 10140 31476
rect 9180 31436 10140 31464
rect 9180 31424 9186 31436
rect 10134 31424 10140 31436
rect 10192 31424 10198 31476
rect 12158 31424 12164 31476
rect 12216 31464 12222 31476
rect 16574 31464 16580 31476
rect 12216 31436 16580 31464
rect 12216 31424 12222 31436
rect 16574 31424 16580 31436
rect 16632 31424 16638 31476
rect 16850 31424 16856 31476
rect 16908 31424 16914 31476
rect 16942 31424 16948 31476
rect 17000 31464 17006 31476
rect 18230 31464 18236 31476
rect 17000 31436 18236 31464
rect 17000 31424 17006 31436
rect 18230 31424 18236 31436
rect 18288 31464 18294 31476
rect 18598 31464 18604 31476
rect 18288 31436 18604 31464
rect 18288 31424 18294 31436
rect 18598 31424 18604 31436
rect 18656 31424 18662 31476
rect 18708 31436 19656 31464
rect 4706 31356 4712 31408
rect 4764 31356 4770 31408
rect 5810 31356 5816 31408
rect 5868 31356 5874 31408
rect 7006 31356 7012 31408
rect 7064 31396 7070 31408
rect 8389 31399 8447 31405
rect 7064 31368 7222 31396
rect 7064 31356 7070 31368
rect 8389 31365 8401 31399
rect 8435 31396 8447 31399
rect 9490 31396 9496 31408
rect 8435 31368 9496 31396
rect 8435 31365 8447 31368
rect 8389 31359 8447 31365
rect 9490 31356 9496 31368
rect 9548 31356 9554 31408
rect 10410 31356 10416 31408
rect 10468 31356 10474 31408
rect 10594 31356 10600 31408
rect 10652 31396 10658 31408
rect 10652 31368 11744 31396
rect 10652 31356 10658 31368
rect 1857 31331 1915 31337
rect 1857 31297 1869 31331
rect 1903 31297 1915 31331
rect 1857 31291 1915 31297
rect 1872 31260 1900 31291
rect 2314 31288 2320 31340
rect 2372 31328 2378 31340
rect 2409 31331 2467 31337
rect 2409 31328 2421 31331
rect 2372 31300 2421 31328
rect 2372 31288 2378 31300
rect 2409 31297 2421 31300
rect 2455 31297 2467 31331
rect 2409 31291 2467 31297
rect 3329 31331 3387 31337
rect 3329 31297 3341 31331
rect 3375 31328 3387 31331
rect 3418 31328 3424 31340
rect 3375 31300 3424 31328
rect 3375 31297 3387 31300
rect 3329 31291 3387 31297
rect 3418 31288 3424 31300
rect 3476 31288 3482 31340
rect 3786 31288 3792 31340
rect 3844 31328 3850 31340
rect 3973 31331 4031 31337
rect 3973 31328 3985 31331
rect 3844 31300 3985 31328
rect 3844 31288 3850 31300
rect 3973 31297 3985 31300
rect 4019 31297 4031 31331
rect 5828 31328 5856 31356
rect 5828 31300 7236 31328
rect 3973 31291 4031 31297
rect 2774 31260 2780 31272
rect 1872 31232 2780 31260
rect 2774 31220 2780 31232
rect 2832 31220 2838 31272
rect 4249 31263 4307 31269
rect 4249 31229 4261 31263
rect 4295 31260 4307 31263
rect 5258 31260 5264 31272
rect 4295 31232 5264 31260
rect 4295 31229 4307 31232
rect 4249 31223 4307 31229
rect 5258 31220 5264 31232
rect 5316 31220 5322 31272
rect 5534 31220 5540 31272
rect 5592 31260 5598 31272
rect 5810 31260 5816 31272
rect 5592 31232 5816 31260
rect 5592 31220 5598 31232
rect 5810 31220 5816 31232
rect 5868 31220 5874 31272
rect 6641 31263 6699 31269
rect 6641 31229 6653 31263
rect 6687 31260 6699 31263
rect 6730 31260 6736 31272
rect 6687 31232 6736 31260
rect 6687 31229 6699 31232
rect 6641 31223 6699 31229
rect 6730 31220 6736 31232
rect 6788 31220 6794 31272
rect 7208 31260 7236 31300
rect 8662 31288 8668 31340
rect 8720 31328 8726 31340
rect 11149 31331 11207 31337
rect 8720 31300 8765 31328
rect 8720 31288 8726 31300
rect 11149 31297 11161 31331
rect 11195 31328 11207 31331
rect 11238 31328 11244 31340
rect 11195 31300 11244 31328
rect 11195 31297 11207 31300
rect 11149 31291 11207 31297
rect 11238 31288 11244 31300
rect 11296 31288 11302 31340
rect 11716 31337 11744 31368
rect 13170 31356 13176 31408
rect 13228 31396 13234 31408
rect 13449 31399 13507 31405
rect 13449 31396 13461 31399
rect 13228 31368 13461 31396
rect 13228 31356 13234 31368
rect 13449 31365 13461 31368
rect 13495 31365 13507 31399
rect 13449 31359 13507 31365
rect 13538 31356 13544 31408
rect 13596 31396 13602 31408
rect 14553 31399 14611 31405
rect 14553 31396 14565 31399
rect 13596 31368 14565 31396
rect 13596 31356 13602 31368
rect 14553 31365 14565 31368
rect 14599 31365 14611 31399
rect 14553 31359 14611 31365
rect 14918 31356 14924 31408
rect 14976 31396 14982 31408
rect 16868 31396 16896 31424
rect 17037 31399 17095 31405
rect 17037 31396 17049 31399
rect 14976 31368 15792 31396
rect 16868 31368 17049 31396
rect 14976 31356 14982 31368
rect 11701 31331 11759 31337
rect 11701 31297 11713 31331
rect 11747 31297 11759 31331
rect 11701 31291 11759 31297
rect 12084 31300 12374 31328
rect 9125 31263 9183 31269
rect 9125 31260 9137 31263
rect 7208 31232 9137 31260
rect 9125 31229 9137 31232
rect 9171 31260 9183 31263
rect 10778 31260 10784 31272
rect 9171 31232 10784 31260
rect 9171 31229 9183 31232
rect 9125 31223 9183 31229
rect 10778 31220 10784 31232
rect 10836 31220 10842 31272
rect 10873 31263 10931 31269
rect 10873 31229 10885 31263
rect 10919 31260 10931 31263
rect 11974 31260 11980 31272
rect 10919 31232 11980 31260
rect 10919 31229 10931 31232
rect 10873 31223 10931 31229
rect 11974 31220 11980 31232
rect 12032 31220 12038 31272
rect 2593 31195 2651 31201
rect 2593 31161 2605 31195
rect 2639 31192 2651 31195
rect 2639 31164 2774 31192
rect 2639 31161 2651 31164
rect 2593 31155 2651 31161
rect 2746 31124 2774 31164
rect 5276 31164 7420 31192
rect 5276 31124 5304 31164
rect 2746 31096 5304 31124
rect 5721 31127 5779 31133
rect 5721 31093 5733 31127
rect 5767 31124 5779 31127
rect 6086 31124 6092 31136
rect 5767 31096 6092 31124
rect 5767 31093 5779 31096
rect 5721 31087 5779 31093
rect 6086 31084 6092 31096
rect 6144 31124 6150 31136
rect 6270 31124 6276 31136
rect 6144 31096 6276 31124
rect 6144 31084 6150 31096
rect 6270 31084 6276 31096
rect 6328 31084 6334 31136
rect 7392 31124 7420 31164
rect 11238 31152 11244 31204
rect 11296 31192 11302 31204
rect 12084 31192 12112 31300
rect 13722 31288 13728 31340
rect 13780 31328 13786 31340
rect 15105 31331 15163 31337
rect 13780 31300 13825 31328
rect 13780 31288 13786 31300
rect 15105 31297 15117 31331
rect 15151 31328 15163 31331
rect 15562 31328 15568 31340
rect 15151 31300 15568 31328
rect 15151 31297 15163 31300
rect 15105 31291 15163 31297
rect 15562 31288 15568 31300
rect 15620 31288 15626 31340
rect 15764 31337 15792 31368
rect 17037 31365 17049 31368
rect 17083 31365 17095 31399
rect 17037 31359 17095 31365
rect 15749 31331 15807 31337
rect 15749 31297 15761 31331
rect 15795 31297 15807 31331
rect 15749 31291 15807 31297
rect 15838 31288 15844 31340
rect 15896 31328 15902 31340
rect 16298 31328 16304 31340
rect 15896 31300 16304 31328
rect 15896 31288 15902 31300
rect 16298 31288 16304 31300
rect 16356 31288 16362 31340
rect 17954 31288 17960 31340
rect 18012 31328 18018 31340
rect 18601 31331 18659 31337
rect 18601 31328 18613 31331
rect 18012 31300 18613 31328
rect 18012 31288 18018 31300
rect 18601 31297 18613 31300
rect 18647 31297 18659 31331
rect 18601 31291 18659 31297
rect 11296 31164 12112 31192
rect 12360 31232 14228 31260
rect 11296 31152 11302 31164
rect 12360 31124 12388 31232
rect 14200 31192 14228 31232
rect 14274 31220 14280 31272
rect 14332 31260 14338 31272
rect 14461 31263 14519 31269
rect 14461 31260 14473 31263
rect 14332 31232 14473 31260
rect 14332 31220 14338 31232
rect 14461 31229 14473 31232
rect 14507 31229 14519 31263
rect 16022 31260 16028 31272
rect 14461 31223 14519 31229
rect 14844 31232 16028 31260
rect 14844 31192 14872 31232
rect 16022 31220 16028 31232
rect 16080 31220 16086 31272
rect 16945 31263 17003 31269
rect 16945 31229 16957 31263
rect 16991 31229 17003 31263
rect 17862 31260 17868 31272
rect 17823 31232 17868 31260
rect 16945 31223 17003 31229
rect 16960 31192 16988 31223
rect 17862 31220 17868 31232
rect 17920 31220 17926 31272
rect 18708 31260 18736 31436
rect 19628 31405 19656 31436
rect 19978 31424 19984 31476
rect 20036 31464 20042 31476
rect 20349 31467 20407 31473
rect 20349 31464 20361 31467
rect 20036 31436 20361 31464
rect 20036 31424 20042 31436
rect 20349 31433 20361 31436
rect 20395 31433 20407 31467
rect 20990 31464 20996 31476
rect 20951 31436 20996 31464
rect 20349 31427 20407 31433
rect 20990 31424 20996 31436
rect 21048 31424 21054 31476
rect 21266 31424 21272 31476
rect 21324 31464 21330 31476
rect 22097 31467 22155 31473
rect 22097 31464 22109 31467
rect 21324 31436 22109 31464
rect 21324 31424 21330 31436
rect 22097 31433 22109 31436
rect 22143 31433 22155 31467
rect 22097 31427 22155 31433
rect 22922 31424 22928 31476
rect 22980 31464 22986 31476
rect 23109 31467 23167 31473
rect 23109 31464 23121 31467
rect 22980 31436 23121 31464
rect 22980 31424 22986 31436
rect 23109 31433 23121 31436
rect 23155 31433 23167 31467
rect 23109 31427 23167 31433
rect 19613 31399 19671 31405
rect 19613 31365 19625 31399
rect 19659 31365 19671 31399
rect 19613 31359 19671 31365
rect 19705 31399 19763 31405
rect 19705 31365 19717 31399
rect 19751 31396 19763 31399
rect 20622 31396 20628 31408
rect 19751 31368 20628 31396
rect 19751 31365 19763 31368
rect 19705 31359 19763 31365
rect 20622 31356 20628 31368
rect 20680 31356 20686 31408
rect 20441 31331 20499 31337
rect 20441 31297 20453 31331
rect 20487 31328 20499 31331
rect 20530 31328 20536 31340
rect 20487 31300 20536 31328
rect 20487 31297 20499 31300
rect 20441 31291 20499 31297
rect 20530 31288 20536 31300
rect 20588 31288 20594 31340
rect 20898 31328 20904 31340
rect 20859 31300 20904 31328
rect 20898 31288 20904 31300
rect 20956 31288 20962 31340
rect 17972 31232 18736 31260
rect 17770 31192 17776 31204
rect 14200 31164 14872 31192
rect 15120 31164 15976 31192
rect 16960 31164 17776 31192
rect 7392 31096 12388 31124
rect 13354 31084 13360 31136
rect 13412 31124 13418 31136
rect 15120 31124 15148 31164
rect 13412 31096 15148 31124
rect 13412 31084 13418 31096
rect 15746 31084 15752 31136
rect 15804 31124 15810 31136
rect 15841 31127 15899 31133
rect 15841 31124 15853 31127
rect 15804 31096 15853 31124
rect 15804 31084 15810 31096
rect 15841 31093 15853 31096
rect 15887 31093 15899 31127
rect 15948 31124 15976 31164
rect 17770 31152 17776 31164
rect 17828 31152 17834 31204
rect 17972 31124 18000 31232
rect 18874 31220 18880 31272
rect 18932 31260 18938 31272
rect 22094 31260 22100 31272
rect 18932 31232 22100 31260
rect 18932 31220 18938 31232
rect 22094 31220 22100 31232
rect 22152 31260 22158 31272
rect 22462 31260 22468 31272
rect 22152 31232 22468 31260
rect 22152 31220 22158 31232
rect 22462 31220 22468 31232
rect 22520 31220 22526 31272
rect 18414 31152 18420 31204
rect 18472 31192 18478 31204
rect 19153 31195 19211 31201
rect 19153 31192 19165 31195
rect 18472 31164 19165 31192
rect 18472 31152 18478 31164
rect 19153 31161 19165 31164
rect 19199 31161 19211 31195
rect 22557 31195 22615 31201
rect 22557 31192 22569 31195
rect 19153 31155 19211 31161
rect 22066 31164 22569 31192
rect 18506 31124 18512 31136
rect 15948 31096 18000 31124
rect 18467 31096 18512 31124
rect 15841 31087 15899 31093
rect 18506 31084 18512 31096
rect 18564 31084 18570 31136
rect 18598 31084 18604 31136
rect 18656 31124 18662 31136
rect 22066 31124 22094 31164
rect 22557 31161 22569 31164
rect 22603 31161 22615 31195
rect 22557 31155 22615 31161
rect 18656 31096 22094 31124
rect 18656 31084 18662 31096
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 3329 30923 3387 30929
rect 3329 30889 3341 30923
rect 3375 30920 3387 30923
rect 6914 30920 6920 30932
rect 3375 30892 6920 30920
rect 3375 30889 3387 30892
rect 3329 30883 3387 30889
rect 6914 30880 6920 30892
rect 6972 30880 6978 30932
rect 7926 30880 7932 30932
rect 7984 30920 7990 30932
rect 11514 30920 11520 30932
rect 7984 30892 11520 30920
rect 7984 30880 7990 30892
rect 11514 30880 11520 30892
rect 11572 30880 11578 30932
rect 11974 30880 11980 30932
rect 12032 30920 12038 30932
rect 12032 30892 12664 30920
rect 12032 30880 12038 30892
rect 6362 30812 6368 30864
rect 6420 30852 6426 30864
rect 6420 30824 7033 30852
rect 6420 30812 6426 30824
rect 3973 30787 4031 30793
rect 3973 30753 3985 30787
rect 4019 30784 4031 30787
rect 4246 30784 4252 30796
rect 4019 30756 4252 30784
rect 4019 30753 4031 30756
rect 3973 30747 4031 30753
rect 4246 30744 4252 30756
rect 4304 30744 4310 30796
rect 5442 30784 5448 30796
rect 5355 30756 5448 30784
rect 5442 30744 5448 30756
rect 5500 30784 5506 30796
rect 6549 30787 6607 30793
rect 6549 30784 6561 30787
rect 5500 30756 6561 30784
rect 5500 30744 5506 30756
rect 6549 30753 6561 30756
rect 6595 30753 6607 30787
rect 7005 30784 7033 30824
rect 9306 30812 9312 30864
rect 9364 30852 9370 30864
rect 10594 30852 10600 30864
rect 9364 30824 10600 30852
rect 9364 30812 9370 30824
rect 10594 30812 10600 30824
rect 10652 30852 10658 30864
rect 10870 30852 10876 30864
rect 10652 30824 10876 30852
rect 10652 30812 10658 30824
rect 10870 30812 10876 30824
rect 10928 30812 10934 30864
rect 8297 30787 8355 30793
rect 8297 30784 8309 30787
rect 7005 30756 8309 30784
rect 6549 30747 6607 30753
rect 8297 30753 8309 30756
rect 8343 30753 8355 30787
rect 11606 30784 11612 30796
rect 8297 30747 8355 30753
rect 8772 30756 11612 30784
rect 1857 30719 1915 30725
rect 1857 30685 1869 30719
rect 1903 30716 1915 30719
rect 1946 30716 1952 30728
rect 1903 30688 1952 30716
rect 1903 30685 1915 30688
rect 1857 30679 1915 30685
rect 1946 30676 1952 30688
rect 2004 30676 2010 30728
rect 2317 30719 2375 30725
rect 2317 30685 2329 30719
rect 2363 30685 2375 30719
rect 2317 30679 2375 30685
rect 2332 30648 2360 30679
rect 2866 30676 2872 30728
rect 2924 30716 2930 30728
rect 3237 30719 3295 30725
rect 3237 30716 3249 30719
rect 2924 30688 3249 30716
rect 2924 30676 2930 30688
rect 3237 30685 3249 30688
rect 3283 30716 3295 30719
rect 4062 30716 4068 30728
rect 3283 30688 4068 30716
rect 3283 30685 3295 30688
rect 3237 30679 3295 30685
rect 4062 30676 4068 30688
rect 4120 30676 4126 30728
rect 5718 30676 5724 30728
rect 5776 30716 5782 30728
rect 8573 30719 8631 30725
rect 5776 30688 5869 30716
rect 5776 30676 5782 30688
rect 8573 30685 8585 30719
rect 8619 30716 8631 30719
rect 8662 30716 8668 30728
rect 8619 30688 8668 30716
rect 8619 30685 8631 30688
rect 8573 30679 8631 30685
rect 8662 30676 8668 30688
rect 8720 30676 8726 30728
rect 1872 30620 2360 30648
rect 1872 30592 1900 30620
rect 4798 30608 4804 30660
rect 4856 30608 4862 30660
rect 5534 30608 5540 30660
rect 5592 30648 5598 30660
rect 5736 30648 5764 30676
rect 5592 30620 5764 30648
rect 5592 30608 5598 30620
rect 6914 30608 6920 30660
rect 6972 30648 6978 30660
rect 6972 30620 7130 30648
rect 6972 30608 6978 30620
rect 1670 30580 1676 30592
rect 1631 30552 1676 30580
rect 1670 30540 1676 30552
rect 1728 30540 1734 30592
rect 1854 30540 1860 30592
rect 1912 30540 1918 30592
rect 2406 30580 2412 30592
rect 2367 30552 2412 30580
rect 2406 30540 2412 30552
rect 2464 30540 2470 30592
rect 3234 30540 3240 30592
rect 3292 30580 3298 30592
rect 8772 30580 8800 30756
rect 11606 30744 11612 30756
rect 11664 30744 11670 30796
rect 11977 30787 12035 30793
rect 11977 30753 11989 30787
rect 12023 30784 12035 30787
rect 12342 30784 12348 30796
rect 12023 30756 12348 30784
rect 12023 30753 12035 30756
rect 11977 30747 12035 30753
rect 12342 30744 12348 30756
rect 12400 30744 12406 30796
rect 12636 30784 12664 30892
rect 12710 30880 12716 30932
rect 12768 30920 12774 30932
rect 13633 30923 13691 30929
rect 13633 30920 13645 30923
rect 12768 30892 13645 30920
rect 12768 30880 12774 30892
rect 13633 30889 13645 30892
rect 13679 30889 13691 30923
rect 13633 30883 13691 30889
rect 15654 30880 15660 30932
rect 15712 30920 15718 30932
rect 16022 30920 16028 30932
rect 15712 30892 16028 30920
rect 15712 30880 15718 30892
rect 16022 30880 16028 30892
rect 16080 30880 16086 30932
rect 18414 30880 18420 30932
rect 18472 30920 18478 30932
rect 23014 30920 23020 30932
rect 18472 30892 21956 30920
rect 22975 30892 23020 30920
rect 18472 30880 18478 30892
rect 12802 30812 12808 30864
rect 12860 30852 12866 30864
rect 13722 30852 13728 30864
rect 12860 30824 13728 30852
rect 12860 30812 12866 30824
rect 13722 30812 13728 30824
rect 13780 30812 13786 30864
rect 14550 30812 14556 30864
rect 14608 30852 14614 30864
rect 14737 30855 14795 30861
rect 14737 30852 14749 30855
rect 14608 30824 14749 30852
rect 14608 30812 14614 30824
rect 14737 30821 14749 30824
rect 14783 30821 14795 30855
rect 14737 30815 14795 30821
rect 15562 30812 15568 30864
rect 15620 30852 15626 30864
rect 15933 30855 15991 30861
rect 15933 30852 15945 30855
rect 15620 30824 15945 30852
rect 15620 30812 15626 30824
rect 15933 30821 15945 30824
rect 15979 30852 15991 30855
rect 17773 30855 17831 30861
rect 17773 30852 17785 30855
rect 15979 30824 17785 30852
rect 15979 30821 15991 30824
rect 15933 30815 15991 30821
rect 17773 30821 17785 30824
rect 17819 30852 17831 30855
rect 17819 30824 21404 30852
rect 17819 30821 17831 30824
rect 17773 30815 17831 30821
rect 13446 30784 13452 30796
rect 12636 30756 13452 30784
rect 13446 30744 13452 30756
rect 13504 30744 13510 30796
rect 14660 30756 20300 30784
rect 9582 30716 9588 30728
rect 9543 30688 9588 30716
rect 9582 30676 9588 30688
rect 9640 30676 9646 30728
rect 10226 30716 10232 30728
rect 10187 30688 10232 30716
rect 10226 30676 10232 30688
rect 10284 30716 10290 30728
rect 10594 30716 10600 30728
rect 10284 30688 10600 30716
rect 10284 30676 10290 30688
rect 10594 30676 10600 30688
rect 10652 30676 10658 30728
rect 12253 30719 12311 30725
rect 12253 30685 12265 30719
rect 12299 30716 12311 30719
rect 12802 30716 12808 30728
rect 12299 30688 12808 30716
rect 12299 30685 12311 30688
rect 12253 30679 12311 30685
rect 12802 30676 12808 30688
rect 12860 30676 12866 30728
rect 13078 30676 13084 30728
rect 13136 30716 13142 30728
rect 14660 30725 14688 30756
rect 13725 30719 13783 30725
rect 13725 30716 13737 30719
rect 13136 30688 13737 30716
rect 13136 30676 13142 30688
rect 13725 30685 13737 30688
rect 13771 30685 13783 30719
rect 13725 30679 13783 30685
rect 14645 30719 14703 30725
rect 14645 30685 14657 30719
rect 14691 30685 14703 30719
rect 16666 30716 16672 30728
rect 16627 30688 16672 30716
rect 14645 30679 14703 30685
rect 10502 30608 10508 30660
rect 10560 30648 10566 30660
rect 10560 30620 10810 30648
rect 11624 30620 12664 30648
rect 10560 30608 10566 30620
rect 11624 30592 11652 30620
rect 9674 30580 9680 30592
rect 3292 30552 8800 30580
rect 9635 30552 9680 30580
rect 3292 30540 3298 30552
rect 9674 30540 9680 30552
rect 9732 30540 9738 30592
rect 11606 30540 11612 30592
rect 11664 30540 11670 30592
rect 12636 30580 12664 30620
rect 12710 30608 12716 30660
rect 12768 30648 12774 30660
rect 12989 30651 13047 30657
rect 12989 30648 13001 30651
rect 12768 30620 13001 30648
rect 12768 30608 12774 30620
rect 12989 30617 13001 30620
rect 13035 30617 13047 30651
rect 12989 30611 13047 30617
rect 14660 30580 14688 30679
rect 16666 30676 16672 30688
rect 16724 30676 16730 30728
rect 18414 30676 18420 30728
rect 18472 30716 18478 30728
rect 18509 30719 18567 30725
rect 18509 30716 18521 30719
rect 18472 30688 18521 30716
rect 18472 30676 18478 30688
rect 18509 30685 18521 30688
rect 18555 30685 18567 30719
rect 18509 30679 18567 30685
rect 15381 30651 15439 30657
rect 15381 30617 15393 30651
rect 15427 30617 15439 30651
rect 15381 30611 15439 30617
rect 12636 30552 14688 30580
rect 15396 30580 15424 30611
rect 15470 30608 15476 30660
rect 15528 30648 15534 30660
rect 15528 30620 15573 30648
rect 15528 30608 15534 30620
rect 17034 30608 17040 30660
rect 17092 30648 17098 30660
rect 17221 30651 17279 30657
rect 17221 30648 17233 30651
rect 17092 30620 17233 30648
rect 17092 30608 17098 30620
rect 17221 30617 17233 30620
rect 17267 30617 17279 30651
rect 17221 30611 17279 30617
rect 17310 30608 17316 30660
rect 17368 30648 17374 30660
rect 17368 30620 17413 30648
rect 17368 30608 17374 30620
rect 18782 30608 18788 30660
rect 18840 30648 18846 30660
rect 19521 30651 19579 30657
rect 19521 30648 19533 30651
rect 18840 30620 19533 30648
rect 18840 30608 18846 30620
rect 19521 30617 19533 30620
rect 19567 30617 19579 30651
rect 19521 30611 19579 30617
rect 19613 30651 19671 30657
rect 19613 30617 19625 30651
rect 19659 30648 19671 30651
rect 19978 30648 19984 30660
rect 19659 30620 19984 30648
rect 19659 30617 19671 30620
rect 19613 30611 19671 30617
rect 19978 30608 19984 30620
rect 20036 30608 20042 30660
rect 20165 30651 20223 30657
rect 20165 30617 20177 30651
rect 20211 30617 20223 30651
rect 20272 30648 20300 30756
rect 20530 30744 20536 30796
rect 20588 30784 20594 30796
rect 21269 30787 21327 30793
rect 21269 30784 21281 30787
rect 20588 30756 21281 30784
rect 20588 30744 20594 30756
rect 21269 30753 21281 30756
rect 21315 30753 21327 30787
rect 21269 30747 21327 30753
rect 20809 30719 20867 30725
rect 20809 30685 20821 30719
rect 20855 30716 20867 30719
rect 20898 30716 20904 30728
rect 20855 30688 20904 30716
rect 20855 30685 20867 30688
rect 20809 30679 20867 30685
rect 20898 30676 20904 30688
rect 20956 30676 20962 30728
rect 21376 30716 21404 30824
rect 21928 30793 21956 30892
rect 23014 30880 23020 30892
rect 23072 30880 23078 30932
rect 21913 30787 21971 30793
rect 21913 30753 21925 30787
rect 21959 30784 21971 30787
rect 25682 30784 25688 30796
rect 21959 30756 25688 30784
rect 21959 30753 21971 30756
rect 21913 30747 21971 30753
rect 25682 30744 25688 30756
rect 25740 30744 25746 30796
rect 24118 30716 24124 30728
rect 21376 30688 24124 30716
rect 24118 30676 24124 30688
rect 24176 30676 24182 30728
rect 23014 30648 23020 30660
rect 20272 30620 23020 30648
rect 20165 30611 20223 30617
rect 15654 30580 15660 30592
rect 15396 30552 15660 30580
rect 15654 30540 15660 30552
rect 15712 30540 15718 30592
rect 16574 30580 16580 30592
rect 16535 30552 16580 30580
rect 16574 30540 16580 30552
rect 16632 30540 16638 30592
rect 18414 30580 18420 30592
rect 18375 30552 18420 30580
rect 18414 30540 18420 30552
rect 18472 30540 18478 30592
rect 19334 30540 19340 30592
rect 19392 30580 19398 30592
rect 20180 30580 20208 30611
rect 23014 30608 23020 30620
rect 23072 30608 23078 30660
rect 20714 30580 20720 30592
rect 19392 30552 20208 30580
rect 20675 30552 20720 30580
rect 19392 30540 19398 30552
rect 20714 30540 20720 30552
rect 20772 30540 20778 30592
rect 22094 30540 22100 30592
rect 22152 30580 22158 30592
rect 22373 30583 22431 30589
rect 22373 30580 22385 30583
rect 22152 30552 22385 30580
rect 22152 30540 22158 30552
rect 22373 30549 22385 30552
rect 22419 30549 22431 30583
rect 22373 30543 22431 30549
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 4246 30336 4252 30388
rect 4304 30376 4310 30388
rect 5902 30376 5908 30388
rect 4304 30348 5908 30376
rect 4304 30336 4310 30348
rect 5902 30336 5908 30348
rect 5960 30376 5966 30388
rect 6362 30376 6368 30388
rect 5960 30348 6368 30376
rect 5960 30336 5966 30348
rect 6362 30336 6368 30348
rect 6420 30336 6426 30388
rect 9674 30336 9680 30388
rect 9732 30376 9738 30388
rect 13998 30376 14004 30388
rect 9732 30348 14004 30376
rect 9732 30336 9738 30348
rect 13998 30336 14004 30348
rect 14056 30336 14062 30388
rect 14274 30336 14280 30388
rect 14332 30376 14338 30388
rect 15930 30376 15936 30388
rect 14332 30348 15936 30376
rect 14332 30336 14338 30348
rect 15930 30336 15936 30348
rect 15988 30336 15994 30388
rect 16209 30379 16267 30385
rect 16209 30345 16221 30379
rect 16255 30376 16267 30379
rect 16850 30376 16856 30388
rect 16255 30348 16856 30376
rect 16255 30345 16267 30348
rect 16209 30339 16267 30345
rect 16850 30336 16856 30348
rect 16908 30376 16914 30388
rect 18782 30376 18788 30388
rect 16908 30348 18788 30376
rect 16908 30336 16914 30348
rect 18782 30336 18788 30348
rect 18840 30336 18846 30388
rect 19058 30336 19064 30388
rect 19116 30376 19122 30388
rect 20714 30376 20720 30388
rect 19116 30348 20720 30376
rect 19116 30336 19122 30348
rect 20714 30336 20720 30348
rect 20772 30336 20778 30388
rect 3418 30268 3424 30320
rect 3476 30308 3482 30320
rect 3602 30308 3608 30320
rect 3476 30280 3608 30308
rect 3476 30268 3482 30280
rect 3602 30268 3608 30280
rect 3660 30268 3666 30320
rect 6822 30308 6828 30320
rect 5290 30280 6828 30308
rect 6822 30268 6828 30280
rect 6880 30268 6886 30320
rect 8662 30268 8668 30320
rect 8720 30308 8726 30320
rect 10413 30311 10471 30317
rect 8720 30280 9076 30308
rect 8720 30268 8726 30280
rect 2406 30200 2412 30252
rect 2464 30200 2470 30252
rect 3786 30200 3792 30252
rect 3844 30240 3850 30252
rect 3844 30212 3889 30240
rect 3844 30200 3850 30212
rect 5994 30200 6000 30252
rect 6052 30240 6058 30252
rect 6052 30212 6097 30240
rect 6052 30200 6058 30212
rect 6730 30200 6736 30252
rect 6788 30240 6794 30252
rect 6788 30212 7682 30240
rect 6788 30200 6794 30212
rect 3418 30132 3424 30184
rect 3476 30172 3482 30184
rect 3513 30175 3571 30181
rect 3513 30172 3525 30175
rect 3476 30144 3525 30172
rect 3476 30132 3482 30144
rect 3513 30141 3525 30144
rect 3559 30141 3571 30175
rect 5258 30172 5264 30184
rect 3513 30135 3571 30141
rect 3712 30144 5264 30172
rect 2041 30039 2099 30045
rect 2041 30005 2053 30039
rect 2087 30036 2099 30039
rect 3712 30036 3740 30144
rect 5258 30132 5264 30144
rect 5316 30132 5322 30184
rect 5721 30175 5779 30181
rect 5721 30141 5733 30175
rect 5767 30172 5779 30175
rect 7009 30175 7067 30181
rect 5767 30144 6224 30172
rect 5767 30141 5779 30144
rect 5721 30135 5779 30141
rect 6196 30104 6224 30144
rect 7009 30141 7021 30175
rect 7055 30172 7067 30175
rect 7098 30172 7104 30184
rect 7055 30144 7104 30172
rect 7055 30141 7067 30144
rect 7009 30135 7067 30141
rect 7098 30132 7104 30144
rect 7156 30172 7162 30184
rect 7282 30172 7288 30184
rect 7156 30144 7288 30172
rect 7156 30132 7162 30144
rect 7282 30132 7288 30144
rect 7340 30132 7346 30184
rect 7742 30132 7748 30184
rect 7800 30172 7806 30184
rect 8294 30172 8300 30184
rect 7800 30144 8300 30172
rect 7800 30132 7806 30144
rect 8294 30132 8300 30144
rect 8352 30132 8358 30184
rect 9048 30181 9076 30280
rect 10413 30277 10425 30311
rect 10459 30308 10471 30311
rect 11882 30308 11888 30320
rect 10459 30280 11888 30308
rect 10459 30277 10471 30280
rect 10413 30271 10471 30277
rect 11882 30268 11888 30280
rect 11940 30268 11946 30320
rect 11974 30268 11980 30320
rect 12032 30308 12038 30320
rect 15473 30311 15531 30317
rect 15473 30308 15485 30311
rect 12032 30280 12077 30308
rect 13924 30280 15485 30308
rect 12032 30268 12038 30280
rect 9861 30243 9919 30249
rect 9861 30209 9873 30243
rect 9907 30240 9919 30243
rect 10042 30240 10048 30252
rect 9907 30212 10048 30240
rect 9907 30209 9919 30212
rect 9861 30203 9919 30209
rect 10042 30200 10048 30212
rect 10100 30200 10106 30252
rect 10318 30240 10324 30252
rect 10279 30212 10324 30240
rect 10318 30200 10324 30212
rect 10376 30200 10382 30252
rect 10962 30240 10968 30252
rect 10923 30212 10968 30240
rect 10962 30200 10968 30212
rect 11020 30200 11026 30252
rect 11054 30200 11060 30252
rect 11112 30240 11118 30252
rect 11606 30240 11612 30252
rect 11112 30212 11612 30240
rect 11112 30200 11118 30212
rect 11606 30200 11612 30212
rect 11664 30200 11670 30252
rect 13078 30200 13084 30252
rect 13136 30200 13142 30252
rect 8757 30175 8815 30181
rect 8757 30141 8769 30175
rect 8803 30172 8815 30175
rect 9033 30175 9091 30181
rect 8803 30144 8984 30172
rect 8803 30141 8815 30144
rect 8757 30135 8815 30141
rect 7760 30104 7788 30132
rect 6196 30076 7788 30104
rect 8956 30104 8984 30144
rect 9033 30141 9045 30175
rect 9079 30172 9091 30175
rect 11330 30172 11336 30184
rect 9079 30144 11336 30172
rect 9079 30141 9091 30144
rect 9033 30135 9091 30141
rect 11330 30132 11336 30144
rect 11388 30172 11394 30184
rect 11698 30172 11704 30184
rect 11388 30144 11704 30172
rect 11388 30132 11394 30144
rect 11698 30132 11704 30144
rect 11756 30132 11762 30184
rect 12066 30132 12072 30184
rect 12124 30172 12130 30184
rect 13924 30172 13952 30280
rect 15473 30277 15485 30280
rect 15519 30277 15531 30311
rect 15473 30271 15531 30277
rect 15838 30268 15844 30320
rect 15896 30308 15902 30320
rect 17037 30311 17095 30317
rect 17037 30308 17049 30311
rect 15896 30280 17049 30308
rect 15896 30268 15902 30280
rect 17037 30277 17049 30280
rect 17083 30277 17095 30311
rect 17037 30271 17095 30277
rect 17770 30268 17776 30320
rect 17828 30308 17834 30320
rect 19334 30308 19340 30320
rect 17828 30280 19340 30308
rect 17828 30268 17834 30280
rect 19334 30268 19340 30280
rect 19392 30268 19398 30320
rect 19518 30308 19524 30320
rect 19479 30280 19524 30308
rect 19518 30268 19524 30280
rect 19576 30268 19582 30320
rect 19794 30268 19800 30320
rect 19852 30308 19858 30320
rect 20349 30311 20407 30317
rect 20349 30308 20361 30311
rect 19852 30280 20361 30308
rect 19852 30268 19858 30280
rect 20349 30277 20361 30280
rect 20395 30277 20407 30311
rect 20349 30271 20407 30277
rect 21453 30311 21511 30317
rect 21453 30277 21465 30311
rect 21499 30308 21511 30311
rect 22094 30308 22100 30320
rect 21499 30280 22100 30308
rect 21499 30277 21511 30280
rect 21453 30271 21511 30277
rect 22094 30268 22100 30280
rect 22152 30268 22158 30320
rect 14274 30200 14280 30252
rect 14332 30240 14338 30252
rect 14461 30243 14519 30249
rect 14461 30240 14473 30243
rect 14332 30212 14473 30240
rect 14332 30200 14338 30212
rect 14461 30209 14473 30212
rect 14507 30240 14519 30243
rect 14918 30240 14924 30252
rect 14507 30212 14924 30240
rect 14507 30209 14519 30212
rect 14461 30203 14519 30209
rect 14918 30200 14924 30212
rect 14976 30200 14982 30252
rect 16301 30243 16359 30249
rect 16301 30209 16313 30243
rect 16347 30240 16359 30243
rect 16666 30240 16672 30252
rect 16347 30212 16672 30240
rect 16347 30209 16359 30212
rect 16301 30203 16359 30209
rect 16666 30200 16672 30212
rect 16724 30200 16730 30252
rect 20901 30243 20959 30249
rect 19812 30212 20024 30240
rect 12124 30144 13952 30172
rect 12124 30132 12130 30144
rect 14550 30132 14556 30184
rect 14608 30172 14614 30184
rect 15562 30172 15568 30184
rect 14608 30144 15424 30172
rect 15523 30144 15568 30172
rect 14608 30132 14614 30144
rect 9306 30104 9312 30116
rect 8956 30076 9312 30104
rect 9306 30064 9312 30076
rect 9364 30064 9370 30116
rect 9769 30107 9827 30113
rect 9769 30073 9781 30107
rect 9815 30104 9827 30107
rect 13446 30104 13452 30116
rect 9815 30076 11192 30104
rect 13407 30076 13452 30104
rect 9815 30073 9827 30076
rect 9769 30067 9827 30073
rect 2087 30008 3740 30036
rect 4249 30039 4307 30045
rect 2087 30005 2099 30008
rect 2041 29999 2099 30005
rect 4249 30005 4261 30039
rect 4295 30036 4307 30039
rect 4614 30036 4620 30048
rect 4295 30008 4620 30036
rect 4295 30005 4307 30008
rect 4249 29999 4307 30005
rect 4614 29996 4620 30008
rect 4672 29996 4678 30048
rect 5534 29996 5540 30048
rect 5592 30036 5598 30048
rect 5994 30036 6000 30048
rect 5592 30008 6000 30036
rect 5592 29996 5598 30008
rect 5994 29996 6000 30008
rect 6052 29996 6058 30048
rect 6270 29996 6276 30048
rect 6328 30036 6334 30048
rect 10318 30036 10324 30048
rect 6328 30008 10324 30036
rect 6328 29996 6334 30008
rect 10318 29996 10324 30008
rect 10376 29996 10382 30048
rect 11054 30036 11060 30048
rect 11015 30008 11060 30036
rect 11054 29996 11060 30008
rect 11112 29996 11118 30048
rect 11164 30036 11192 30076
rect 13446 30064 13452 30076
rect 13504 30064 13510 30116
rect 14642 30064 14648 30116
rect 14700 30104 14706 30116
rect 15013 30107 15071 30113
rect 15013 30104 15025 30107
rect 14700 30076 15025 30104
rect 14700 30064 14706 30076
rect 15013 30073 15025 30076
rect 15059 30073 15071 30107
rect 15396 30104 15424 30144
rect 15562 30132 15568 30144
rect 15620 30132 15626 30184
rect 16758 30132 16764 30184
rect 16816 30172 16822 30184
rect 16945 30175 17003 30181
rect 16945 30172 16957 30175
rect 16816 30144 16957 30172
rect 16816 30132 16822 30144
rect 16945 30141 16957 30144
rect 16991 30141 17003 30175
rect 17862 30172 17868 30184
rect 17823 30144 17868 30172
rect 16945 30135 17003 30141
rect 17862 30132 17868 30144
rect 17920 30132 17926 30184
rect 18046 30132 18052 30184
rect 18104 30172 18110 30184
rect 18969 30175 19027 30181
rect 18969 30172 18981 30175
rect 18104 30144 18981 30172
rect 18104 30132 18110 30144
rect 18969 30141 18981 30144
rect 19015 30141 19027 30175
rect 18969 30135 19027 30141
rect 19150 30132 19156 30184
rect 19208 30172 19214 30184
rect 19613 30175 19671 30181
rect 19613 30172 19625 30175
rect 19208 30144 19625 30172
rect 19208 30132 19214 30144
rect 19613 30141 19625 30144
rect 19659 30172 19671 30175
rect 19812 30172 19840 30212
rect 19659 30144 19840 30172
rect 19659 30141 19671 30144
rect 19613 30135 19671 30141
rect 19794 30104 19800 30116
rect 15396 30076 19800 30104
rect 15013 30067 15071 30073
rect 19794 30064 19800 30076
rect 19852 30064 19858 30116
rect 19996 30104 20024 30212
rect 20901 30209 20913 30243
rect 20947 30240 20959 30243
rect 21542 30240 21548 30252
rect 20947 30212 21548 30240
rect 20947 30209 20959 30212
rect 20901 30203 20959 30209
rect 21542 30200 21548 30212
rect 21600 30200 21606 30252
rect 20070 30132 20076 30184
rect 20128 30172 20134 30184
rect 20257 30175 20315 30181
rect 20257 30172 20269 30175
rect 20128 30144 20269 30172
rect 20128 30132 20134 30144
rect 20257 30141 20269 30144
rect 20303 30141 20315 30175
rect 22005 30175 22063 30181
rect 22005 30172 22017 30175
rect 20257 30135 20315 30141
rect 20824 30144 22017 30172
rect 20714 30104 20720 30116
rect 19996 30076 20720 30104
rect 20714 30064 20720 30076
rect 20772 30064 20778 30116
rect 13170 30036 13176 30048
rect 11164 30008 13176 30036
rect 13170 29996 13176 30008
rect 13228 29996 13234 30048
rect 13722 29996 13728 30048
rect 13780 30036 13786 30048
rect 14369 30039 14427 30045
rect 14369 30036 14381 30039
rect 13780 30008 14381 30036
rect 13780 29996 13786 30008
rect 14369 30005 14381 30008
rect 14415 30005 14427 30039
rect 14369 29999 14427 30005
rect 14826 29996 14832 30048
rect 14884 30036 14890 30048
rect 17126 30036 17132 30048
rect 14884 30008 17132 30036
rect 14884 29996 14890 30008
rect 17126 29996 17132 30008
rect 17184 29996 17190 30048
rect 18322 29996 18328 30048
rect 18380 30036 18386 30048
rect 18417 30039 18475 30045
rect 18417 30036 18429 30039
rect 18380 30008 18429 30036
rect 18380 29996 18386 30008
rect 18417 30005 18429 30008
rect 18463 30005 18475 30039
rect 18417 29999 18475 30005
rect 19886 29996 19892 30048
rect 19944 30036 19950 30048
rect 20824 30036 20852 30144
rect 22005 30141 22017 30144
rect 22051 30141 22063 30175
rect 22005 30135 22063 30141
rect 37826 30132 37832 30184
rect 37884 30172 37890 30184
rect 38013 30175 38071 30181
rect 38013 30172 38025 30175
rect 37884 30144 38025 30172
rect 37884 30132 37890 30144
rect 38013 30141 38025 30144
rect 38059 30141 38071 30175
rect 38286 30172 38292 30184
rect 38247 30144 38292 30172
rect 38013 30135 38071 30141
rect 38286 30132 38292 30144
rect 38344 30132 38350 30184
rect 20898 30064 20904 30116
rect 20956 30104 20962 30116
rect 20956 30076 22692 30104
rect 20956 30064 20962 30076
rect 22664 30045 22692 30076
rect 19944 30008 20852 30036
rect 22649 30039 22707 30045
rect 19944 29996 19950 30008
rect 22649 30005 22661 30039
rect 22695 30036 22707 30039
rect 22922 30036 22928 30048
rect 22695 30008 22928 30036
rect 22695 30005 22707 30008
rect 22649 29999 22707 30005
rect 22922 29996 22928 30008
rect 22980 29996 22986 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 1762 29792 1768 29844
rect 1820 29792 1826 29844
rect 6638 29792 6644 29844
rect 6696 29832 6702 29844
rect 6733 29835 6791 29841
rect 6733 29832 6745 29835
rect 6696 29804 6745 29832
rect 6696 29792 6702 29804
rect 6733 29801 6745 29804
rect 6779 29801 6791 29835
rect 6733 29795 6791 29801
rect 6822 29792 6828 29844
rect 6880 29832 6886 29844
rect 11330 29832 11336 29844
rect 6880 29804 11336 29832
rect 6880 29792 6886 29804
rect 11330 29792 11336 29804
rect 11388 29792 11394 29844
rect 13078 29792 13084 29844
rect 13136 29832 13142 29844
rect 18506 29832 18512 29844
rect 13136 29804 18512 29832
rect 13136 29792 13142 29804
rect 18506 29792 18512 29804
rect 18564 29792 18570 29844
rect 19518 29792 19524 29844
rect 19576 29832 19582 29844
rect 21085 29835 21143 29841
rect 21085 29832 21097 29835
rect 19576 29804 21097 29832
rect 19576 29792 19582 29804
rect 21085 29801 21097 29804
rect 21131 29801 21143 29835
rect 38286 29832 38292 29844
rect 38247 29804 38292 29832
rect 21085 29795 21143 29801
rect 38286 29792 38292 29804
rect 38344 29792 38350 29844
rect 1780 29696 1808 29792
rect 7377 29767 7435 29773
rect 7377 29764 7389 29767
rect 7300 29736 7389 29764
rect 1949 29699 2007 29705
rect 1949 29696 1961 29699
rect 1780 29668 1961 29696
rect 1949 29665 1961 29668
rect 1995 29696 2007 29699
rect 2406 29696 2412 29708
rect 1995 29668 2412 29696
rect 1995 29665 2007 29668
rect 1949 29659 2007 29665
rect 2406 29656 2412 29668
rect 2464 29656 2470 29708
rect 3421 29699 3479 29705
rect 3421 29665 3433 29699
rect 3467 29696 3479 29699
rect 3602 29696 3608 29708
rect 3467 29668 3608 29696
rect 3467 29665 3479 29668
rect 3421 29659 3479 29665
rect 3602 29656 3608 29668
rect 3660 29656 3666 29708
rect 3786 29656 3792 29708
rect 3844 29696 3850 29708
rect 3973 29699 4031 29705
rect 3973 29696 3985 29699
rect 3844 29668 3985 29696
rect 3844 29656 3850 29668
rect 3973 29665 3985 29668
rect 4019 29696 4031 29699
rect 5534 29696 5540 29708
rect 4019 29668 5540 29696
rect 4019 29665 4031 29668
rect 3973 29659 4031 29665
rect 5534 29656 5540 29668
rect 5592 29656 5598 29708
rect 5718 29656 5724 29708
rect 5776 29656 5782 29708
rect 6730 29656 6736 29708
rect 6788 29696 6794 29708
rect 7300 29696 7328 29736
rect 7377 29733 7389 29736
rect 7423 29733 7435 29767
rect 7377 29727 7435 29733
rect 8021 29767 8079 29773
rect 8021 29733 8033 29767
rect 8067 29764 8079 29767
rect 9858 29764 9864 29776
rect 8067 29736 9864 29764
rect 8067 29733 8079 29736
rect 8021 29727 8079 29733
rect 9858 29724 9864 29736
rect 9916 29724 9922 29776
rect 12618 29724 12624 29776
rect 12676 29764 12682 29776
rect 13446 29764 13452 29776
rect 12676 29736 13452 29764
rect 12676 29724 12682 29736
rect 13446 29724 13452 29736
rect 13504 29724 13510 29776
rect 15470 29764 15476 29776
rect 13740 29736 15476 29764
rect 6788 29668 7328 29696
rect 6788 29656 6794 29668
rect 8294 29656 8300 29708
rect 8352 29696 8358 29708
rect 10410 29696 10416 29708
rect 8352 29668 10416 29696
rect 8352 29656 8358 29668
rect 10410 29656 10416 29668
rect 10468 29656 10474 29708
rect 11238 29696 11244 29708
rect 10520 29668 11244 29696
rect 1673 29631 1731 29637
rect 1673 29597 1685 29631
rect 1719 29597 1731 29631
rect 1673 29591 1731 29597
rect 1688 29504 1716 29591
rect 3050 29588 3056 29640
rect 3108 29588 3114 29640
rect 5736 29628 5764 29656
rect 6270 29628 6276 29640
rect 5736 29600 6276 29628
rect 6270 29588 6276 29600
rect 6328 29628 6334 29640
rect 6641 29631 6699 29637
rect 7929 29631 7987 29637
rect 6641 29628 6653 29631
rect 6328 29600 6653 29628
rect 6328 29588 6334 29600
rect 6641 29597 6653 29600
rect 6687 29597 6699 29631
rect 6641 29591 6699 29597
rect 7277 29625 7335 29631
rect 7277 29591 7289 29625
rect 7323 29591 7335 29625
rect 7929 29597 7941 29631
rect 7975 29597 7987 29631
rect 9306 29628 9312 29640
rect 9267 29600 9312 29628
rect 7929 29591 7987 29597
rect 7277 29585 7335 29591
rect 4249 29563 4307 29569
rect 4249 29529 4261 29563
rect 4295 29529 4307 29563
rect 6822 29560 6828 29572
rect 5474 29532 6828 29560
rect 4249 29523 4307 29529
rect 1670 29492 1676 29504
rect 1583 29464 1676 29492
rect 1670 29452 1676 29464
rect 1728 29492 1734 29504
rect 3234 29492 3240 29504
rect 1728 29464 3240 29492
rect 1728 29452 1734 29464
rect 3234 29452 3240 29464
rect 3292 29492 3298 29504
rect 3786 29492 3792 29504
rect 3292 29464 3792 29492
rect 3292 29452 3298 29464
rect 3786 29452 3792 29464
rect 3844 29452 3850 29504
rect 4264 29492 4292 29523
rect 6822 29520 6828 29532
rect 6880 29520 6886 29572
rect 4614 29492 4620 29504
rect 4264 29464 4620 29492
rect 4614 29452 4620 29464
rect 4672 29492 4678 29504
rect 4890 29492 4896 29504
rect 4672 29464 4896 29492
rect 4672 29452 4678 29464
rect 4890 29452 4896 29464
rect 4948 29452 4954 29504
rect 5626 29452 5632 29504
rect 5684 29492 5690 29504
rect 5721 29495 5779 29501
rect 5721 29492 5733 29495
rect 5684 29464 5733 29492
rect 5684 29452 5690 29464
rect 5721 29461 5733 29464
rect 5767 29492 5779 29495
rect 5810 29492 5816 29504
rect 5767 29464 5816 29492
rect 5767 29461 5779 29464
rect 5721 29455 5779 29461
rect 5810 29452 5816 29464
rect 5868 29452 5874 29504
rect 5994 29452 6000 29504
rect 6052 29492 6058 29504
rect 6914 29492 6920 29504
rect 6052 29464 6920 29492
rect 6052 29452 6058 29464
rect 6914 29452 6920 29464
rect 6972 29452 6978 29504
rect 7300 29492 7328 29585
rect 7944 29560 7972 29591
rect 9306 29588 9312 29600
rect 9364 29588 9370 29640
rect 9582 29588 9588 29640
rect 9640 29628 9646 29640
rect 10520 29628 10548 29668
rect 11238 29656 11244 29668
rect 11296 29656 11302 29708
rect 11698 29656 11704 29708
rect 11756 29696 11762 29708
rect 11977 29699 12035 29705
rect 11977 29696 11989 29699
rect 11756 29668 11989 29696
rect 11756 29656 11762 29668
rect 11977 29665 11989 29668
rect 12023 29665 12035 29699
rect 13262 29696 13268 29708
rect 13223 29668 13268 29696
rect 11977 29659 12035 29665
rect 13262 29656 13268 29668
rect 13320 29656 13326 29708
rect 9640 29600 10548 29628
rect 9640 29588 9646 29600
rect 9122 29560 9128 29572
rect 7944 29532 9128 29560
rect 8036 29504 8064 29532
rect 9122 29520 9128 29532
rect 9180 29520 9186 29572
rect 9490 29520 9496 29572
rect 9548 29560 9554 29572
rect 9674 29560 9680 29572
rect 9548 29532 9680 29560
rect 9548 29520 9554 29532
rect 9674 29520 9680 29532
rect 9732 29560 9738 29572
rect 9953 29563 10011 29569
rect 9953 29560 9965 29563
rect 9732 29532 9965 29560
rect 9732 29520 9738 29532
rect 9953 29529 9965 29532
rect 9999 29560 10011 29563
rect 10134 29560 10140 29572
rect 9999 29532 10140 29560
rect 9999 29529 10011 29532
rect 9953 29523 10011 29529
rect 10134 29520 10140 29532
rect 10192 29520 10198 29572
rect 10226 29520 10232 29572
rect 10284 29560 10290 29572
rect 10284 29532 10534 29560
rect 10284 29520 10290 29532
rect 11606 29520 11612 29572
rect 11664 29560 11670 29572
rect 11701 29563 11759 29569
rect 11701 29560 11713 29563
rect 11664 29532 11713 29560
rect 11664 29520 11670 29532
rect 11701 29529 11713 29532
rect 11747 29529 11759 29563
rect 11701 29523 11759 29529
rect 11790 29520 11796 29572
rect 11848 29560 11854 29572
rect 12621 29563 12679 29569
rect 12621 29560 12633 29563
rect 11848 29532 12633 29560
rect 11848 29520 11854 29532
rect 12621 29529 12633 29532
rect 12667 29529 12679 29563
rect 13170 29560 13176 29572
rect 13131 29532 13176 29560
rect 12621 29523 12679 29529
rect 13170 29520 13176 29532
rect 13228 29520 13234 29572
rect 7926 29492 7932 29504
rect 7300 29464 7932 29492
rect 7926 29452 7932 29464
rect 7984 29452 7990 29504
rect 8018 29452 8024 29504
rect 8076 29452 8082 29504
rect 8478 29452 8484 29504
rect 8536 29492 8542 29504
rect 8754 29492 8760 29504
rect 8536 29464 8760 29492
rect 8536 29452 8542 29464
rect 8754 29452 8760 29464
rect 8812 29452 8818 29504
rect 9401 29495 9459 29501
rect 9401 29461 9413 29495
rect 9447 29492 9459 29495
rect 13740 29492 13768 29736
rect 15470 29724 15476 29736
rect 15528 29724 15534 29776
rect 16206 29724 16212 29776
rect 16264 29724 16270 29776
rect 16666 29724 16672 29776
rect 16724 29764 16730 29776
rect 20898 29764 20904 29776
rect 16724 29736 20904 29764
rect 16724 29724 16730 29736
rect 20898 29724 20904 29736
rect 20956 29724 20962 29776
rect 13814 29656 13820 29708
rect 13872 29696 13878 29708
rect 14642 29696 14648 29708
rect 13872 29668 14648 29696
rect 13872 29656 13878 29668
rect 14642 29656 14648 29668
rect 14700 29656 14706 29708
rect 14921 29699 14979 29705
rect 14921 29665 14933 29699
rect 14967 29696 14979 29699
rect 16224 29696 16252 29724
rect 14967 29668 16252 29696
rect 14967 29665 14979 29668
rect 14921 29659 14979 29665
rect 18046 29656 18052 29708
rect 18104 29696 18110 29708
rect 18141 29699 18199 29705
rect 18141 29696 18153 29699
rect 18104 29668 18153 29696
rect 18104 29656 18110 29668
rect 18141 29665 18153 29668
rect 18187 29665 18199 29699
rect 18782 29696 18788 29708
rect 18743 29668 18788 29696
rect 18141 29659 18199 29665
rect 18782 29656 18788 29668
rect 18840 29656 18846 29708
rect 18966 29656 18972 29708
rect 19024 29696 19030 29708
rect 20070 29696 20076 29708
rect 19024 29668 20076 29696
rect 19024 29656 19030 29668
rect 20070 29656 20076 29668
rect 20128 29656 20134 29708
rect 20165 29699 20223 29705
rect 20165 29665 20177 29699
rect 20211 29696 20223 29699
rect 20438 29696 20444 29708
rect 20211 29668 20444 29696
rect 20211 29665 20223 29668
rect 20165 29659 20223 29665
rect 20438 29656 20444 29668
rect 20496 29656 20502 29708
rect 22094 29696 22100 29708
rect 21192 29668 22100 29696
rect 13906 29588 13912 29640
rect 13964 29588 13970 29640
rect 21192 29637 21220 29668
rect 22094 29656 22100 29668
rect 22152 29656 22158 29708
rect 21177 29631 21235 29637
rect 21177 29597 21189 29631
rect 21223 29597 21235 29631
rect 21177 29591 21235 29597
rect 21821 29631 21879 29637
rect 21821 29597 21833 29631
rect 21867 29628 21879 29631
rect 21910 29628 21916 29640
rect 21867 29600 21916 29628
rect 21867 29597 21879 29600
rect 21821 29591 21879 29597
rect 21910 29588 21916 29600
rect 21968 29628 21974 29640
rect 21968 29600 22094 29628
rect 21968 29588 21974 29600
rect 13924 29560 13952 29588
rect 14829 29563 14887 29569
rect 14829 29560 14841 29563
rect 13924 29532 14841 29560
rect 14829 29529 14841 29532
rect 14875 29529 14887 29563
rect 14829 29523 14887 29529
rect 14918 29520 14924 29572
rect 14976 29560 14982 29572
rect 15657 29563 15715 29569
rect 15657 29560 15669 29563
rect 14976 29532 15669 29560
rect 14976 29520 14982 29532
rect 15657 29529 15669 29532
rect 15703 29529 15715 29563
rect 15657 29523 15715 29529
rect 15749 29563 15807 29569
rect 15749 29529 15761 29563
rect 15795 29529 15807 29563
rect 15749 29523 15807 29529
rect 9447 29464 13768 29492
rect 9447 29461 9459 29464
rect 9401 29455 9459 29461
rect 13906 29452 13912 29504
rect 13964 29492 13970 29504
rect 14458 29492 14464 29504
rect 13964 29464 14464 29492
rect 13964 29452 13970 29464
rect 14458 29452 14464 29464
rect 14516 29452 14522 29504
rect 15764 29492 15792 29523
rect 15930 29520 15936 29572
rect 15988 29560 15994 29572
rect 16301 29563 16359 29569
rect 16301 29560 16313 29563
rect 15988 29532 16313 29560
rect 15988 29520 15994 29532
rect 16301 29529 16313 29532
rect 16347 29560 16359 29563
rect 16390 29560 16396 29572
rect 16347 29532 16396 29560
rect 16347 29529 16359 29532
rect 16301 29523 16359 29529
rect 16390 29520 16396 29532
rect 16448 29520 16454 29572
rect 17034 29560 17040 29572
rect 16995 29532 17040 29560
rect 17034 29520 17040 29532
rect 17092 29520 17098 29572
rect 17126 29520 17132 29572
rect 17184 29560 17190 29572
rect 17681 29563 17739 29569
rect 17184 29532 17229 29560
rect 17184 29520 17190 29532
rect 17681 29529 17693 29563
rect 17727 29560 17739 29563
rect 17770 29560 17776 29572
rect 17727 29532 17776 29560
rect 17727 29529 17739 29532
rect 17681 29523 17739 29529
rect 17770 29520 17776 29532
rect 17828 29520 17834 29572
rect 18690 29560 18696 29572
rect 18651 29532 18696 29560
rect 18690 29520 18696 29532
rect 18748 29520 18754 29572
rect 20070 29520 20076 29572
rect 20128 29560 20134 29572
rect 20254 29560 20260 29572
rect 20128 29532 20260 29560
rect 20128 29520 20134 29532
rect 20254 29520 20260 29532
rect 20312 29520 20318 29572
rect 20349 29563 20407 29569
rect 20349 29529 20361 29563
rect 20395 29529 20407 29563
rect 20349 29523 20407 29529
rect 16574 29492 16580 29504
rect 15764 29464 16580 29492
rect 16574 29452 16580 29464
rect 16632 29452 16638 29504
rect 16666 29452 16672 29504
rect 16724 29492 16730 29504
rect 19058 29492 19064 29504
rect 16724 29464 19064 29492
rect 16724 29452 16730 29464
rect 19058 29452 19064 29464
rect 19116 29492 19122 29504
rect 19886 29492 19892 29504
rect 19116 29464 19892 29492
rect 19116 29452 19122 29464
rect 19886 29452 19892 29464
rect 19944 29452 19950 29504
rect 20364 29492 20392 29523
rect 20438 29520 20444 29572
rect 20496 29560 20502 29572
rect 20496 29532 20541 29560
rect 20496 29520 20502 29532
rect 20990 29492 20996 29504
rect 20364 29464 20996 29492
rect 20990 29452 20996 29464
rect 21048 29452 21054 29504
rect 21726 29492 21732 29504
rect 21687 29464 21732 29492
rect 21726 29452 21732 29464
rect 21784 29452 21790 29504
rect 22066 29492 22094 29600
rect 22373 29495 22431 29501
rect 22373 29492 22385 29495
rect 22066 29464 22385 29492
rect 22373 29461 22385 29464
rect 22419 29492 22431 29495
rect 38010 29492 38016 29504
rect 22419 29464 38016 29492
rect 22419 29461 22431 29464
rect 22373 29455 22431 29461
rect 38010 29452 38016 29464
rect 38068 29452 38074 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 1670 29288 1676 29300
rect 1631 29260 1676 29288
rect 1670 29248 1676 29260
rect 1728 29248 1734 29300
rect 2225 29291 2283 29297
rect 2225 29257 2237 29291
rect 2271 29288 2283 29291
rect 4798 29288 4804 29300
rect 2271 29260 4804 29288
rect 2271 29257 2283 29260
rect 2225 29251 2283 29257
rect 4798 29248 4804 29260
rect 4856 29248 4862 29300
rect 4985 29291 5043 29297
rect 4985 29257 4997 29291
rect 5031 29288 5043 29291
rect 5626 29288 5632 29300
rect 5031 29260 5632 29288
rect 5031 29257 5043 29260
rect 4985 29251 5043 29257
rect 5626 29248 5632 29260
rect 5684 29248 5690 29300
rect 5905 29291 5963 29297
rect 5905 29257 5917 29291
rect 5951 29288 5963 29291
rect 5994 29288 6000 29300
rect 5951 29260 6000 29288
rect 5951 29257 5963 29260
rect 5905 29251 5963 29257
rect 5994 29248 6000 29260
rect 6052 29248 6058 29300
rect 7929 29291 7987 29297
rect 7929 29288 7941 29291
rect 6472 29260 7941 29288
rect 5350 29180 5356 29232
rect 5408 29220 5414 29232
rect 6472 29220 6500 29260
rect 7929 29257 7941 29260
rect 7975 29257 7987 29291
rect 7929 29251 7987 29257
rect 8573 29291 8631 29297
rect 8573 29257 8585 29291
rect 8619 29288 8631 29291
rect 8754 29288 8760 29300
rect 8619 29260 8760 29288
rect 8619 29257 8631 29260
rect 8573 29251 8631 29257
rect 8754 29248 8760 29260
rect 8812 29248 8818 29300
rect 10410 29288 10416 29300
rect 10060 29260 10416 29288
rect 6638 29220 6644 29232
rect 5408 29192 6500 29220
rect 6599 29192 6644 29220
rect 5408 29180 5414 29192
rect 6638 29180 6644 29192
rect 6696 29180 6702 29232
rect 8662 29180 8668 29232
rect 8720 29220 8726 29232
rect 8720 29192 8878 29220
rect 8720 29180 8726 29192
rect 9766 29180 9772 29232
rect 9824 29220 9830 29232
rect 10060 29229 10088 29260
rect 10410 29248 10416 29260
rect 10468 29248 10474 29300
rect 11054 29248 11060 29300
rect 11112 29288 11118 29300
rect 19150 29288 19156 29300
rect 11112 29260 13860 29288
rect 11112 29248 11118 29260
rect 10045 29223 10103 29229
rect 10045 29220 10057 29223
rect 9824 29192 10057 29220
rect 9824 29180 9830 29192
rect 10045 29189 10057 29192
rect 10091 29189 10103 29223
rect 10045 29183 10103 29189
rect 10336 29192 11100 29220
rect 1854 29112 1860 29164
rect 1912 29152 1918 29164
rect 2133 29155 2191 29161
rect 2133 29152 2145 29155
rect 1912 29124 2145 29152
rect 1912 29112 1918 29124
rect 2133 29121 2145 29124
rect 2179 29152 2191 29155
rect 2406 29152 2412 29164
rect 2179 29124 2412 29152
rect 2179 29121 2191 29124
rect 2133 29115 2191 29121
rect 2406 29112 2412 29124
rect 2464 29112 2470 29164
rect 3234 29152 3240 29164
rect 3195 29124 3240 29152
rect 3234 29112 3240 29124
rect 3292 29112 3298 29164
rect 4614 29112 4620 29164
rect 4672 29112 4678 29164
rect 5813 29155 5871 29161
rect 5813 29121 5825 29155
rect 5859 29121 5871 29155
rect 5813 29115 5871 29121
rect 6549 29155 6607 29161
rect 6549 29121 6561 29155
rect 6595 29152 6607 29155
rect 6730 29152 6736 29164
rect 6595 29124 6736 29152
rect 6595 29121 6607 29124
rect 6549 29115 6607 29121
rect 2774 29044 2780 29096
rect 2832 29084 2838 29096
rect 4522 29084 4528 29096
rect 2832 29056 4528 29084
rect 2832 29044 2838 29056
rect 4522 29044 4528 29056
rect 4580 29044 4586 29096
rect 5828 29084 5856 29115
rect 6730 29112 6736 29124
rect 6788 29112 6794 29164
rect 7193 29155 7251 29161
rect 7193 29121 7205 29155
rect 7239 29152 7251 29155
rect 7374 29152 7380 29164
rect 7239 29124 7380 29152
rect 7239 29121 7251 29124
rect 7193 29115 7251 29121
rect 7374 29112 7380 29124
rect 7432 29112 7438 29164
rect 8029 29155 8087 29161
rect 8029 29121 8041 29155
rect 8075 29152 8087 29155
rect 8202 29152 8208 29164
rect 8075 29124 8208 29152
rect 8075 29121 8087 29124
rect 8029 29115 8087 29121
rect 8202 29112 8208 29124
rect 8260 29112 8266 29164
rect 10336 29161 10364 29192
rect 10321 29155 10379 29161
rect 10321 29121 10333 29155
rect 10367 29121 10379 29155
rect 10321 29115 10379 29121
rect 10965 29155 11023 29161
rect 10965 29121 10977 29155
rect 11011 29121 11023 29155
rect 10965 29115 11023 29121
rect 6638 29084 6644 29096
rect 5828 29056 6644 29084
rect 6638 29044 6644 29056
rect 6696 29044 6702 29096
rect 10502 29084 10508 29096
rect 7952 29072 9904 29084
rect 10060 29072 10508 29084
rect 7952 29056 10508 29072
rect 6270 28976 6276 29028
rect 6328 29016 6334 29028
rect 7285 29019 7343 29025
rect 6328 28988 7236 29016
rect 6328 28976 6334 28988
rect 3500 28951 3558 28957
rect 3500 28917 3512 28951
rect 3546 28948 3558 28951
rect 3602 28948 3608 28960
rect 3546 28920 3608 28948
rect 3546 28917 3558 28920
rect 3500 28911 3558 28917
rect 3602 28908 3608 28920
rect 3660 28908 3666 28960
rect 4522 28908 4528 28960
rect 4580 28948 4586 28960
rect 4798 28948 4804 28960
rect 4580 28920 4804 28948
rect 4580 28908 4586 28920
rect 4798 28908 4804 28920
rect 4856 28908 4862 28960
rect 7208 28948 7236 28988
rect 7285 28985 7297 29019
rect 7331 29016 7343 29019
rect 7952 29016 7980 29056
rect 9876 29044 10088 29056
rect 10502 29044 10508 29056
rect 10560 29044 10566 29096
rect 10980 29084 11008 29115
rect 10704 29056 11008 29084
rect 11072 29084 11100 29192
rect 11238 29180 11244 29232
rect 11296 29220 11302 29232
rect 12621 29223 12679 29229
rect 11296 29192 12572 29220
rect 11296 29180 11302 29192
rect 11514 29112 11520 29164
rect 11572 29152 11578 29164
rect 12544 29161 12572 29192
rect 12621 29189 12633 29223
rect 12667 29220 12679 29223
rect 13538 29220 13544 29232
rect 12667 29192 13544 29220
rect 12667 29189 12679 29192
rect 12621 29183 12679 29189
rect 13538 29180 13544 29192
rect 13596 29180 13602 29232
rect 13722 29220 13728 29232
rect 13683 29192 13728 29220
rect 13722 29180 13728 29192
rect 13780 29180 13786 29232
rect 13832 29229 13860 29260
rect 17604 29260 19156 29288
rect 13817 29223 13875 29229
rect 13817 29189 13829 29223
rect 13863 29220 13875 29223
rect 14461 29223 14519 29229
rect 14461 29220 14473 29223
rect 13863 29192 14473 29220
rect 13863 29189 13875 29192
rect 13817 29183 13875 29189
rect 14461 29189 14473 29192
rect 14507 29189 14519 29223
rect 14461 29183 14519 29189
rect 14550 29180 14556 29232
rect 14608 29220 14614 29232
rect 15746 29220 15752 29232
rect 14608 29192 14653 29220
rect 15707 29192 15752 29220
rect 14608 29180 14614 29192
rect 15746 29180 15752 29192
rect 15804 29180 15810 29232
rect 15930 29180 15936 29232
rect 15988 29220 15994 29232
rect 16298 29220 16304 29232
rect 15988 29192 16304 29220
rect 15988 29180 15994 29192
rect 16298 29180 16304 29192
rect 16356 29180 16362 29232
rect 17604 29220 17632 29260
rect 19150 29248 19156 29260
rect 19208 29248 19214 29300
rect 19352 29260 20576 29288
rect 16500 29192 17632 29220
rect 17681 29223 17739 29229
rect 11885 29155 11943 29161
rect 11885 29152 11897 29155
rect 11572 29124 11897 29152
rect 11572 29112 11578 29124
rect 11885 29121 11897 29124
rect 11931 29121 11943 29155
rect 12529 29155 12587 29161
rect 11885 29115 11943 29121
rect 11992 29124 12480 29152
rect 11698 29084 11704 29096
rect 11072 29056 11704 29084
rect 10704 29016 10732 29056
rect 11698 29044 11704 29056
rect 11756 29044 11762 29096
rect 11054 29016 11060 29028
rect 7331 28988 7980 29016
rect 8128 28994 9076 29016
rect 10428 28994 10732 29016
rect 8036 28988 9076 28994
rect 7331 28985 7343 28988
rect 7285 28979 7343 28985
rect 8036 28966 8156 28988
rect 8036 28948 8064 28966
rect 7208 28920 8064 28948
rect 9048 28948 9076 28988
rect 10244 28988 10732 28994
rect 11015 28988 11060 29016
rect 10244 28966 10456 28988
rect 11054 28976 11060 28988
rect 11112 28976 11118 29028
rect 11330 28976 11336 29028
rect 11388 29016 11394 29028
rect 11790 29016 11796 29028
rect 11388 28988 11796 29016
rect 11388 28976 11394 28988
rect 11790 28976 11796 28988
rect 11848 28976 11854 29028
rect 11992 29025 12020 29124
rect 12452 29084 12480 29124
rect 12529 29121 12541 29155
rect 12575 29121 12587 29155
rect 12529 29115 12587 29121
rect 13170 29084 13176 29096
rect 12452 29056 13176 29084
rect 13170 29044 13176 29056
rect 13228 29044 13234 29096
rect 13541 29087 13599 29093
rect 13541 29053 13553 29087
rect 13587 29053 13599 29087
rect 13541 29047 13599 29053
rect 11977 29019 12035 29025
rect 11977 28985 11989 29019
rect 12023 28985 12035 29019
rect 13556 29016 13584 29047
rect 14458 29044 14464 29096
rect 14516 29084 14522 29096
rect 15657 29087 15715 29093
rect 15657 29084 15669 29087
rect 14516 29056 15669 29084
rect 14516 29044 14522 29056
rect 15657 29053 15669 29056
rect 15703 29084 15715 29087
rect 16500 29084 16528 29192
rect 17681 29189 17693 29223
rect 17727 29220 17739 29223
rect 18414 29220 18420 29232
rect 17727 29192 18420 29220
rect 17727 29189 17739 29192
rect 17681 29183 17739 29189
rect 18414 29180 18420 29192
rect 18472 29180 18478 29232
rect 19242 29220 19248 29232
rect 19203 29192 19248 29220
rect 19242 29180 19248 29192
rect 19300 29180 19306 29232
rect 19352 29229 19380 29260
rect 19337 29223 19395 29229
rect 19337 29189 19349 29223
rect 19383 29189 19395 29223
rect 19337 29183 19395 29189
rect 19518 29180 19524 29232
rect 19576 29220 19582 29232
rect 19889 29223 19947 29229
rect 19889 29220 19901 29223
rect 19576 29192 19901 29220
rect 19576 29180 19582 29192
rect 19889 29189 19901 29192
rect 19935 29189 19947 29223
rect 20438 29220 20444 29232
rect 20399 29192 20444 29220
rect 19889 29183 19947 29189
rect 20438 29180 20444 29192
rect 20496 29180 20502 29232
rect 20548 29229 20576 29260
rect 20990 29248 20996 29300
rect 21048 29288 21054 29300
rect 21177 29291 21235 29297
rect 21177 29288 21189 29291
rect 21048 29260 21189 29288
rect 21048 29248 21054 29260
rect 21177 29257 21189 29260
rect 21223 29257 21235 29291
rect 21177 29251 21235 29257
rect 23198 29248 23204 29300
rect 23256 29288 23262 29300
rect 23385 29291 23443 29297
rect 23385 29288 23397 29291
rect 23256 29260 23397 29288
rect 23256 29248 23262 29260
rect 23385 29257 23397 29260
rect 23431 29257 23443 29291
rect 23385 29251 23443 29257
rect 20533 29223 20591 29229
rect 20533 29189 20545 29223
rect 20579 29220 20591 29223
rect 21726 29220 21732 29232
rect 20579 29192 21732 29220
rect 20579 29189 20591 29192
rect 20533 29183 20591 29189
rect 21726 29180 21732 29192
rect 21784 29180 21790 29232
rect 16666 29112 16672 29164
rect 16724 29152 16730 29164
rect 17037 29155 17095 29161
rect 17037 29152 17049 29155
rect 16724 29124 17049 29152
rect 16724 29112 16730 29124
rect 17037 29121 17049 29124
rect 17083 29121 17095 29155
rect 17037 29115 17095 29121
rect 20806 29112 20812 29164
rect 20864 29152 20870 29164
rect 21085 29155 21143 29161
rect 21085 29152 21097 29155
rect 20864 29124 21097 29152
rect 20864 29112 20870 29124
rect 21085 29121 21097 29124
rect 21131 29121 21143 29155
rect 21085 29115 21143 29121
rect 22189 29155 22247 29161
rect 22189 29121 22201 29155
rect 22235 29152 22247 29155
rect 23201 29155 23259 29161
rect 22235 29124 22784 29152
rect 22235 29121 22247 29124
rect 22189 29115 22247 29121
rect 15703 29056 16528 29084
rect 15703 29053 15715 29056
rect 15657 29047 15715 29053
rect 16574 29044 16580 29096
rect 16632 29084 16638 29096
rect 17589 29087 17647 29093
rect 17589 29084 17601 29087
rect 16632 29056 17601 29084
rect 16632 29044 16638 29056
rect 17589 29053 17601 29056
rect 17635 29053 17647 29087
rect 17589 29047 17647 29053
rect 18690 29044 18696 29096
rect 18748 29084 18754 29096
rect 22097 29087 22155 29093
rect 22097 29084 22109 29087
rect 18748 29056 22109 29084
rect 18748 29044 18754 29056
rect 22097 29053 22109 29056
rect 22143 29053 22155 29087
rect 22097 29047 22155 29053
rect 15013 29019 15071 29025
rect 13556 28988 14964 29016
rect 11977 28979 12035 28985
rect 10244 28948 10272 28966
rect 9048 28920 10272 28948
rect 14936 28948 14964 28988
rect 15013 28985 15025 29019
rect 15059 29016 15071 29019
rect 16206 29016 16212 29028
rect 15059 28988 16212 29016
rect 15059 28985 15071 28988
rect 15013 28979 15071 28985
rect 16206 28976 16212 28988
rect 16264 28976 16270 29028
rect 16942 29016 16948 29028
rect 16903 28988 16948 29016
rect 16942 28976 16948 28988
rect 17000 28976 17006 29028
rect 17770 28976 17776 29028
rect 17828 29016 17834 29028
rect 18141 29019 18199 29025
rect 18141 29016 18153 29019
rect 17828 28988 18153 29016
rect 17828 28976 17834 28988
rect 18141 28985 18153 28988
rect 18187 29016 18199 29019
rect 18785 29019 18843 29025
rect 18187 28988 18736 29016
rect 18187 28985 18199 28988
rect 18141 28979 18199 28985
rect 15286 28948 15292 28960
rect 14936 28920 15292 28948
rect 15286 28908 15292 28920
rect 15344 28908 15350 28960
rect 15378 28908 15384 28960
rect 15436 28948 15442 28960
rect 18322 28948 18328 28960
rect 15436 28920 18328 28948
rect 15436 28908 15442 28920
rect 18322 28908 18328 28920
rect 18380 28908 18386 28960
rect 18708 28948 18736 28988
rect 18785 28985 18797 29019
rect 18831 29016 18843 29019
rect 19334 29016 19340 29028
rect 18831 28988 19340 29016
rect 18831 28985 18843 28988
rect 18785 28979 18843 28985
rect 19334 28976 19340 28988
rect 19392 28976 19398 29028
rect 21542 29016 21548 29028
rect 20272 28988 21548 29016
rect 20272 28948 20300 28988
rect 21542 28976 21548 28988
rect 21600 28976 21606 29028
rect 22756 29025 22784 29124
rect 23201 29121 23213 29155
rect 23247 29152 23259 29155
rect 23247 29124 23428 29152
rect 23247 29121 23259 29124
rect 23201 29115 23259 29121
rect 23400 29028 23428 29124
rect 24118 29112 24124 29164
rect 24176 29152 24182 29164
rect 30101 29155 30159 29161
rect 30101 29152 30113 29155
rect 24176 29124 30113 29152
rect 24176 29112 24182 29124
rect 30101 29121 30113 29124
rect 30147 29121 30159 29155
rect 30101 29115 30159 29121
rect 38010 29084 38016 29096
rect 37971 29056 38016 29084
rect 38010 29044 38016 29056
rect 38068 29044 38074 29096
rect 38286 29084 38292 29096
rect 38247 29056 38292 29084
rect 38286 29044 38292 29056
rect 38344 29044 38350 29096
rect 22741 29019 22799 29025
rect 22741 28985 22753 29019
rect 22787 29016 22799 29019
rect 23198 29016 23204 29028
rect 22787 28988 23204 29016
rect 22787 28985 22799 28988
rect 22741 28979 22799 28985
rect 23198 28976 23204 28988
rect 23256 28976 23262 29028
rect 23382 28976 23388 29028
rect 23440 29016 23446 29028
rect 23845 29019 23903 29025
rect 23845 29016 23857 29019
rect 23440 28988 23857 29016
rect 23440 28976 23446 28988
rect 23845 28985 23857 28988
rect 23891 28985 23903 29019
rect 23845 28979 23903 28985
rect 30193 29019 30251 29025
rect 30193 28985 30205 29019
rect 30239 29016 30251 29019
rect 36630 29016 36636 29028
rect 30239 28988 36636 29016
rect 30239 28985 30251 28988
rect 30193 28979 30251 28985
rect 36630 28976 36636 28988
rect 36688 28976 36694 29028
rect 18708 28920 20300 28948
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 2225 28747 2283 28753
rect 2225 28713 2237 28747
rect 2271 28744 2283 28747
rect 4614 28744 4620 28756
rect 2271 28716 4620 28744
rect 2271 28713 2283 28716
rect 2225 28707 2283 28713
rect 4614 28704 4620 28716
rect 4672 28704 4678 28756
rect 4709 28747 4767 28753
rect 4709 28713 4721 28747
rect 4755 28744 4767 28747
rect 11790 28744 11796 28756
rect 4755 28716 11796 28744
rect 4755 28713 4767 28716
rect 4709 28707 4767 28713
rect 11790 28704 11796 28716
rect 11848 28704 11854 28756
rect 14366 28744 14372 28756
rect 14327 28716 14372 28744
rect 14366 28704 14372 28716
rect 14424 28704 14430 28756
rect 14826 28704 14832 28756
rect 14884 28744 14890 28756
rect 17218 28744 17224 28756
rect 14884 28716 17224 28744
rect 14884 28704 14890 28716
rect 17218 28704 17224 28716
rect 17276 28704 17282 28756
rect 17678 28704 17684 28756
rect 17736 28744 17742 28756
rect 18509 28747 18567 28753
rect 17736 28716 17908 28744
rect 17736 28704 17742 28716
rect 3970 28636 3976 28688
rect 4028 28676 4034 28688
rect 4065 28679 4123 28685
rect 4065 28676 4077 28679
rect 4028 28648 4077 28676
rect 4028 28636 4034 28648
rect 4065 28645 4077 28648
rect 4111 28645 4123 28679
rect 4065 28639 4123 28645
rect 4154 28636 4160 28688
rect 4212 28676 4218 28688
rect 4982 28676 4988 28688
rect 4212 28648 4988 28676
rect 4212 28636 4218 28648
rect 4982 28636 4988 28648
rect 5040 28636 5046 28688
rect 5350 28676 5356 28688
rect 5311 28648 5356 28676
rect 5350 28636 5356 28648
rect 5408 28636 5414 28688
rect 5997 28679 6055 28685
rect 5997 28645 6009 28679
rect 6043 28676 6055 28679
rect 7006 28676 7012 28688
rect 6043 28648 7012 28676
rect 6043 28645 6055 28648
rect 5997 28639 6055 28645
rect 7006 28636 7012 28648
rect 7064 28636 7070 28688
rect 7282 28636 7288 28688
rect 7340 28636 7346 28688
rect 7837 28679 7895 28685
rect 7837 28645 7849 28679
rect 7883 28676 7895 28679
rect 10226 28676 10232 28688
rect 7883 28648 10232 28676
rect 7883 28645 7895 28648
rect 7837 28639 7895 28645
rect 10226 28636 10232 28648
rect 10284 28636 10290 28688
rect 16114 28636 16120 28688
rect 16172 28676 16178 28688
rect 17770 28676 17776 28688
rect 16172 28648 17776 28676
rect 16172 28636 16178 28648
rect 17770 28636 17776 28648
rect 17828 28636 17834 28688
rect 17880 28685 17908 28716
rect 18509 28713 18521 28747
rect 18555 28744 18567 28747
rect 19242 28744 19248 28756
rect 18555 28716 19248 28744
rect 18555 28713 18567 28716
rect 18509 28707 18567 28713
rect 19242 28704 19248 28716
rect 19300 28704 19306 28756
rect 19521 28747 19579 28753
rect 19521 28713 19533 28747
rect 19567 28744 19579 28747
rect 20438 28744 20444 28756
rect 19567 28716 20444 28744
rect 19567 28713 19579 28716
rect 19521 28707 19579 28713
rect 20438 28704 20444 28716
rect 20496 28704 20502 28756
rect 22554 28704 22560 28756
rect 22612 28744 22618 28756
rect 23290 28744 23296 28756
rect 22612 28716 23296 28744
rect 22612 28704 22618 28716
rect 23290 28704 23296 28716
rect 23348 28704 23354 28756
rect 17865 28679 17923 28685
rect 17865 28645 17877 28679
rect 17911 28645 17923 28679
rect 17865 28639 17923 28645
rect 17954 28636 17960 28688
rect 18012 28676 18018 28688
rect 22189 28679 22247 28685
rect 22189 28676 22201 28679
rect 18012 28648 22201 28676
rect 18012 28636 18018 28648
rect 2869 28611 2927 28617
rect 2869 28577 2881 28611
rect 2915 28608 2927 28611
rect 4706 28608 4712 28620
rect 2915 28580 4712 28608
rect 2915 28577 2927 28580
rect 2869 28571 2927 28577
rect 4706 28568 4712 28580
rect 4764 28568 4770 28620
rect 6638 28568 6644 28620
rect 6696 28568 6702 28620
rect 7300 28608 7328 28636
rect 6932 28580 7328 28608
rect 2133 28543 2191 28549
rect 2133 28509 2145 28543
rect 2179 28540 2191 28543
rect 2406 28540 2412 28552
rect 2179 28512 2412 28540
rect 2179 28509 2191 28512
rect 2133 28503 2191 28509
rect 2406 28500 2412 28512
rect 2464 28540 2470 28552
rect 2777 28543 2835 28549
rect 2777 28540 2789 28543
rect 2464 28512 2789 28540
rect 2464 28500 2470 28512
rect 2777 28509 2789 28512
rect 2823 28540 2835 28543
rect 3973 28543 4031 28549
rect 3973 28540 3985 28543
rect 2823 28512 3985 28540
rect 2823 28509 2835 28512
rect 2777 28503 2835 28509
rect 3973 28509 3985 28512
rect 4019 28509 4031 28543
rect 4614 28540 4620 28552
rect 4575 28512 4620 28540
rect 3973 28503 4031 28509
rect 3988 28472 4016 28503
rect 4614 28500 4620 28512
rect 4672 28540 4678 28552
rect 5258 28540 5264 28552
rect 4672 28512 5264 28540
rect 4672 28500 4678 28512
rect 5258 28500 5264 28512
rect 5316 28500 5322 28552
rect 5905 28543 5963 28549
rect 5905 28509 5917 28543
rect 5951 28540 5963 28543
rect 6656 28540 6684 28568
rect 6932 28549 6960 28580
rect 8662 28568 8668 28620
rect 8720 28608 8726 28620
rect 11422 28608 11428 28620
rect 8720 28580 11428 28608
rect 8720 28568 8726 28580
rect 11422 28568 11428 28580
rect 11480 28568 11486 28620
rect 11698 28568 11704 28620
rect 11756 28608 11762 28620
rect 12069 28611 12127 28617
rect 12069 28608 12081 28611
rect 11756 28580 12081 28608
rect 11756 28568 11762 28580
rect 12069 28577 12081 28580
rect 12115 28577 12127 28611
rect 12069 28571 12127 28577
rect 14921 28611 14979 28617
rect 14921 28577 14933 28611
rect 14967 28608 14979 28611
rect 15102 28608 15108 28620
rect 14967 28580 15108 28608
rect 14967 28577 14979 28580
rect 14921 28571 14979 28577
rect 15102 28568 15108 28580
rect 15160 28568 15166 28620
rect 15565 28611 15623 28617
rect 15565 28577 15577 28611
rect 15611 28608 15623 28611
rect 15746 28608 15752 28620
rect 15611 28580 15752 28608
rect 15611 28577 15623 28580
rect 15565 28571 15623 28577
rect 15746 28568 15752 28580
rect 15804 28608 15810 28620
rect 16574 28608 16580 28620
rect 15804 28580 16580 28608
rect 15804 28568 15810 28580
rect 16574 28568 16580 28580
rect 16632 28568 16638 28620
rect 16669 28611 16727 28617
rect 16669 28577 16681 28611
rect 16715 28608 16727 28611
rect 16850 28608 16856 28620
rect 16715 28580 16856 28608
rect 16715 28577 16727 28580
rect 16669 28571 16727 28577
rect 16850 28568 16856 28580
rect 16908 28568 16914 28620
rect 19886 28608 19892 28620
rect 19352 28580 19892 28608
rect 6917 28543 6975 28549
rect 6917 28540 6929 28543
rect 5951 28512 6929 28540
rect 5951 28509 5963 28512
rect 5905 28503 5963 28509
rect 6917 28509 6929 28512
rect 6963 28509 6975 28543
rect 6917 28503 6975 28509
rect 5920 28472 5948 28503
rect 7282 28500 7288 28552
rect 7340 28540 7346 28552
rect 7745 28543 7803 28549
rect 7745 28540 7757 28543
rect 7340 28512 7757 28540
rect 7340 28500 7346 28512
rect 7745 28509 7757 28512
rect 7791 28540 7803 28543
rect 7926 28540 7932 28552
rect 7791 28512 7932 28540
rect 7791 28509 7803 28512
rect 7745 28503 7803 28509
rect 7926 28500 7932 28512
rect 7984 28500 7990 28552
rect 8018 28500 8024 28552
rect 8076 28540 8082 28552
rect 8573 28543 8631 28549
rect 8573 28540 8585 28543
rect 8076 28512 8585 28540
rect 8076 28500 8082 28512
rect 8573 28509 8585 28512
rect 8619 28540 8631 28543
rect 9030 28540 9036 28552
rect 8619 28512 9036 28540
rect 8619 28509 8631 28512
rect 8573 28503 8631 28509
rect 9030 28500 9036 28512
rect 9088 28500 9094 28552
rect 9609 28543 9667 28549
rect 9609 28509 9621 28543
rect 9655 28540 9667 28543
rect 9655 28509 9674 28540
rect 9609 28503 9674 28509
rect 3988 28444 5948 28472
rect 6730 28432 6736 28484
rect 6788 28472 6794 28484
rect 7009 28475 7067 28481
rect 6788 28444 6960 28472
rect 6788 28432 6794 28444
rect 1670 28404 1676 28416
rect 1631 28376 1676 28404
rect 1670 28364 1676 28376
rect 1728 28364 1734 28416
rect 2590 28364 2596 28416
rect 2648 28404 2654 28416
rect 2774 28404 2780 28416
rect 2648 28376 2780 28404
rect 2648 28364 2654 28376
rect 2774 28364 2780 28376
rect 2832 28364 2838 28416
rect 4246 28364 4252 28416
rect 4304 28404 4310 28416
rect 6822 28404 6828 28416
rect 4304 28376 6828 28404
rect 4304 28364 4310 28376
rect 6822 28364 6828 28376
rect 6880 28364 6886 28416
rect 6932 28404 6960 28444
rect 7009 28441 7021 28475
rect 7055 28472 7067 28475
rect 9214 28472 9220 28484
rect 7055 28444 9220 28472
rect 7055 28441 7067 28444
rect 7009 28435 7067 28441
rect 9214 28432 9220 28444
rect 9272 28432 9278 28484
rect 9306 28432 9312 28484
rect 9364 28472 9370 28484
rect 9646 28472 9674 28503
rect 12250 28500 12256 28552
rect 12308 28540 12314 28552
rect 12897 28543 12955 28549
rect 12897 28540 12909 28543
rect 12308 28512 12909 28540
rect 12308 28500 12314 28512
rect 12897 28509 12909 28512
rect 12943 28509 12955 28543
rect 12897 28503 12955 28509
rect 12986 28500 12992 28552
rect 13044 28540 13050 28552
rect 13262 28540 13268 28552
rect 13044 28512 13268 28540
rect 13044 28500 13050 28512
rect 13262 28500 13268 28512
rect 13320 28540 13326 28552
rect 13541 28543 13599 28549
rect 13541 28540 13553 28543
rect 13320 28512 13553 28540
rect 13320 28500 13326 28512
rect 13541 28509 13553 28512
rect 13587 28509 13599 28543
rect 18417 28543 18475 28549
rect 18417 28540 18429 28543
rect 13541 28503 13599 28509
rect 17972 28512 18429 28540
rect 9364 28444 9674 28472
rect 9364 28432 9370 28444
rect 11146 28432 11152 28484
rect 11204 28432 11210 28484
rect 11793 28475 11851 28481
rect 11793 28441 11805 28475
rect 11839 28472 11851 28475
rect 11839 28444 12848 28472
rect 11839 28441 11851 28444
rect 11793 28435 11851 28441
rect 8481 28407 8539 28413
rect 8481 28404 8493 28407
rect 6932 28376 8493 28404
rect 8481 28373 8493 28376
rect 8527 28373 8539 28407
rect 8481 28367 8539 28373
rect 9677 28407 9735 28413
rect 9677 28373 9689 28407
rect 9723 28404 9735 28407
rect 9766 28404 9772 28416
rect 9723 28376 9772 28404
rect 9723 28373 9735 28376
rect 9677 28367 9735 28373
rect 9766 28364 9772 28376
rect 9824 28364 9830 28416
rect 9950 28364 9956 28416
rect 10008 28404 10014 28416
rect 10321 28407 10379 28413
rect 10321 28404 10333 28407
rect 10008 28376 10333 28404
rect 10008 28364 10014 28376
rect 10321 28373 10333 28376
rect 10367 28404 10379 28407
rect 10962 28404 10968 28416
rect 10367 28376 10968 28404
rect 10367 28373 10379 28376
rect 10321 28367 10379 28373
rect 10962 28364 10968 28376
rect 11020 28364 11026 28416
rect 11698 28364 11704 28416
rect 11756 28404 11762 28416
rect 11900 28404 11928 28444
rect 12820 28416 12848 28444
rect 13170 28432 13176 28484
rect 13228 28472 13234 28484
rect 15013 28475 15071 28481
rect 15013 28472 15025 28475
rect 13228 28444 15025 28472
rect 13228 28432 13234 28444
rect 15013 28441 15025 28444
rect 15059 28441 15071 28475
rect 15013 28435 15071 28441
rect 15194 28432 15200 28484
rect 15252 28472 15258 28484
rect 16025 28475 16083 28481
rect 16025 28472 16037 28475
rect 15252 28444 16037 28472
rect 15252 28432 15258 28444
rect 16025 28441 16037 28444
rect 16071 28441 16083 28475
rect 16025 28435 16083 28441
rect 16390 28432 16396 28484
rect 16448 28472 16454 28484
rect 16577 28475 16635 28481
rect 16577 28472 16589 28475
rect 16448 28444 16589 28472
rect 16448 28432 16454 28444
rect 16577 28441 16589 28444
rect 16623 28441 16635 28475
rect 16577 28435 16635 28441
rect 17313 28475 17371 28481
rect 17313 28441 17325 28475
rect 17359 28441 17371 28475
rect 17313 28435 17371 28441
rect 17405 28475 17463 28481
rect 17405 28441 17417 28475
rect 17451 28441 17463 28475
rect 17405 28435 17463 28441
rect 11756 28376 11928 28404
rect 11756 28364 11762 28376
rect 12802 28364 12808 28416
rect 12860 28364 12866 28416
rect 12989 28407 13047 28413
rect 12989 28373 13001 28407
rect 13035 28404 13047 28407
rect 13354 28404 13360 28416
rect 13035 28376 13360 28404
rect 13035 28373 13047 28376
rect 12989 28367 13047 28373
rect 13354 28364 13360 28376
rect 13412 28364 13418 28416
rect 13633 28407 13691 28413
rect 13633 28373 13645 28407
rect 13679 28404 13691 28407
rect 13722 28404 13728 28416
rect 13679 28376 13728 28404
rect 13679 28373 13691 28376
rect 13633 28367 13691 28373
rect 13722 28364 13728 28376
rect 13780 28364 13786 28416
rect 15562 28364 15568 28416
rect 15620 28404 15626 28416
rect 17328 28404 17356 28435
rect 15620 28376 17356 28404
rect 17420 28404 17448 28435
rect 17678 28432 17684 28484
rect 17736 28472 17742 28484
rect 17972 28472 18000 28512
rect 18417 28509 18429 28512
rect 18463 28540 18475 28543
rect 19352 28540 19380 28580
rect 19886 28568 19892 28580
rect 19944 28568 19950 28620
rect 19978 28568 19984 28620
rect 20036 28608 20042 28620
rect 20441 28611 20499 28617
rect 20441 28608 20453 28611
rect 20036 28580 20453 28608
rect 20036 28568 20042 28580
rect 20441 28577 20453 28580
rect 20487 28577 20499 28611
rect 20441 28571 20499 28577
rect 18463 28512 19380 28540
rect 19429 28543 19487 28549
rect 18463 28509 18475 28512
rect 18417 28503 18475 28509
rect 19429 28509 19441 28543
rect 19475 28540 19487 28543
rect 19518 28540 19524 28552
rect 19475 28512 19524 28540
rect 19475 28509 19487 28512
rect 19429 28503 19487 28509
rect 19518 28500 19524 28512
rect 19576 28500 19582 28552
rect 19610 28500 19616 28552
rect 19668 28540 19674 28552
rect 20162 28540 20168 28552
rect 19668 28512 20168 28540
rect 19668 28500 19674 28512
rect 20162 28500 20168 28512
rect 20220 28500 20226 28552
rect 20533 28543 20591 28549
rect 20533 28509 20545 28543
rect 20579 28540 20591 28543
rect 20806 28540 20812 28552
rect 20579 28512 20812 28540
rect 20579 28509 20591 28512
rect 20533 28503 20591 28509
rect 20806 28500 20812 28512
rect 20864 28500 20870 28552
rect 21192 28549 21220 28648
rect 22189 28645 22201 28648
rect 22235 28676 22247 28679
rect 23750 28676 23756 28688
rect 22235 28648 23756 28676
rect 22235 28645 22247 28648
rect 22189 28639 22247 28645
rect 23750 28636 23756 28648
rect 23808 28636 23814 28688
rect 38286 28676 38292 28688
rect 38247 28648 38292 28676
rect 38286 28636 38292 28648
rect 38344 28636 38350 28688
rect 21726 28608 21732 28620
rect 21639 28580 21732 28608
rect 21726 28568 21732 28580
rect 21784 28608 21790 28620
rect 21784 28580 28994 28608
rect 21784 28568 21790 28580
rect 21177 28543 21235 28549
rect 21177 28509 21189 28543
rect 21223 28509 21235 28543
rect 21177 28503 21235 28509
rect 21085 28475 21143 28481
rect 21085 28472 21097 28475
rect 17736 28444 18000 28472
rect 18156 28444 21097 28472
rect 17736 28432 17742 28444
rect 18156 28404 18184 28444
rect 21085 28441 21097 28444
rect 21131 28441 21143 28475
rect 22741 28475 22799 28481
rect 22741 28472 22753 28475
rect 21085 28435 21143 28441
rect 22204 28444 22753 28472
rect 17420 28376 18184 28404
rect 15620 28364 15626 28376
rect 19518 28364 19524 28416
rect 19576 28404 19582 28416
rect 20530 28404 20536 28416
rect 19576 28376 20536 28404
rect 19576 28364 19582 28376
rect 20530 28364 20536 28376
rect 20588 28404 20594 28416
rect 22204 28404 22232 28444
rect 22741 28441 22753 28444
rect 22787 28441 22799 28475
rect 22741 28435 22799 28441
rect 20588 28376 22232 28404
rect 28966 28404 28994 28580
rect 38010 28472 38016 28484
rect 31726 28444 38016 28472
rect 31726 28404 31754 28444
rect 38010 28432 38016 28444
rect 38068 28432 38074 28484
rect 28966 28376 31754 28404
rect 20588 28364 20594 28376
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 2774 28160 2780 28212
rect 2832 28200 2838 28212
rect 4985 28203 5043 28209
rect 4985 28200 4997 28203
rect 2832 28172 4997 28200
rect 2832 28160 2838 28172
rect 4985 28169 4997 28172
rect 5031 28169 5043 28203
rect 4985 28163 5043 28169
rect 5258 28160 5264 28212
rect 5316 28200 5322 28212
rect 7466 28200 7472 28212
rect 5316 28172 7472 28200
rect 5316 28160 5322 28172
rect 2409 28135 2467 28141
rect 2409 28101 2421 28135
rect 2455 28132 2467 28135
rect 4062 28132 4068 28144
rect 2455 28104 4068 28132
rect 2455 28101 2467 28104
rect 2409 28095 2467 28101
rect 4062 28092 4068 28104
rect 4120 28092 4126 28144
rect 1673 28067 1731 28073
rect 1673 28033 1685 28067
rect 1719 28064 1731 28067
rect 1762 28064 1768 28076
rect 1719 28036 1768 28064
rect 1719 28033 1731 28036
rect 1673 28027 1731 28033
rect 1762 28024 1768 28036
rect 1820 28024 1826 28076
rect 2317 28067 2375 28073
rect 2317 28033 2329 28067
rect 2363 28064 2375 28067
rect 2961 28067 3019 28073
rect 2363 28036 2452 28064
rect 2363 28033 2375 28036
rect 2317 28027 2375 28033
rect 2424 28008 2452 28036
rect 2961 28033 2973 28067
rect 3007 28064 3019 28067
rect 3234 28064 3240 28076
rect 3007 28036 3240 28064
rect 3007 28033 3019 28036
rect 2961 28027 3019 28033
rect 3234 28024 3240 28036
rect 3292 28024 3298 28076
rect 3605 28067 3663 28073
rect 3605 28033 3617 28067
rect 3651 28064 3663 28067
rect 3786 28064 3792 28076
rect 3651 28036 3792 28064
rect 3651 28033 3663 28036
rect 3605 28027 3663 28033
rect 2406 27956 2412 28008
rect 2464 27996 2470 28008
rect 2590 27996 2596 28008
rect 2464 27968 2596 27996
rect 2464 27956 2470 27968
rect 2590 27956 2596 27968
rect 2648 27956 2654 28008
rect 2866 27956 2872 28008
rect 2924 27996 2930 28008
rect 3620 27996 3648 28027
rect 3786 28024 3792 28036
rect 3844 28024 3850 28076
rect 4249 28067 4307 28073
rect 4249 28033 4261 28067
rect 4295 28064 4307 28067
rect 4614 28064 4620 28076
rect 4295 28036 4620 28064
rect 4295 28033 4307 28036
rect 4249 28027 4307 28033
rect 4614 28024 4620 28036
rect 4672 28024 4678 28076
rect 5077 28067 5135 28073
rect 5077 28033 5089 28067
rect 5123 28064 5135 28067
rect 5258 28064 5264 28076
rect 5123 28036 5264 28064
rect 5123 28033 5135 28036
rect 5077 28027 5135 28033
rect 5258 28024 5264 28036
rect 5316 28024 5322 28076
rect 5736 28062 5764 28172
rect 7466 28160 7472 28172
rect 7524 28160 7530 28212
rect 7561 28203 7619 28209
rect 7561 28169 7573 28203
rect 7607 28200 7619 28203
rect 7650 28200 7656 28212
rect 7607 28172 7656 28200
rect 7607 28169 7619 28172
rect 7561 28163 7619 28169
rect 7650 28160 7656 28172
rect 7708 28160 7714 28212
rect 9766 28160 9772 28212
rect 9824 28200 9830 28212
rect 9824 28172 12434 28200
rect 9824 28160 9830 28172
rect 6917 28135 6975 28141
rect 6917 28101 6929 28135
rect 6963 28132 6975 28135
rect 8294 28132 8300 28144
rect 6963 28104 8300 28132
rect 6963 28101 6975 28104
rect 6917 28095 6975 28101
rect 8294 28092 8300 28104
rect 8352 28092 8358 28144
rect 10042 28092 10048 28144
rect 10100 28092 10106 28144
rect 10226 28092 10232 28144
rect 10284 28132 10290 28144
rect 11885 28135 11943 28141
rect 11885 28132 11897 28135
rect 10284 28104 11897 28132
rect 10284 28092 10290 28104
rect 11885 28101 11897 28104
rect 11931 28101 11943 28135
rect 12406 28132 12434 28172
rect 12526 28160 12532 28212
rect 12584 28200 12590 28212
rect 16114 28200 16120 28212
rect 12584 28172 16120 28200
rect 12584 28160 12590 28172
rect 16114 28160 16120 28172
rect 16172 28160 16178 28212
rect 22005 28203 22063 28209
rect 22005 28200 22017 28203
rect 17512 28172 22017 28200
rect 13449 28135 13507 28141
rect 13449 28132 13461 28135
rect 12406 28104 13461 28132
rect 11885 28095 11943 28101
rect 13449 28101 13461 28104
rect 13495 28101 13507 28135
rect 13449 28095 13507 28101
rect 13541 28135 13599 28141
rect 13541 28101 13553 28135
rect 13587 28132 13599 28135
rect 14918 28132 14924 28144
rect 13587 28104 14924 28132
rect 13587 28101 13599 28104
rect 13541 28095 13599 28101
rect 14918 28092 14924 28104
rect 14976 28092 14982 28144
rect 15013 28135 15071 28141
rect 15013 28101 15025 28135
rect 15059 28132 15071 28135
rect 15059 28104 16068 28132
rect 15059 28101 15071 28104
rect 15013 28095 15071 28101
rect 5813 28067 5871 28073
rect 5813 28062 5825 28067
rect 5736 28034 5825 28062
rect 5813 28033 5825 28034
rect 5859 28033 5871 28067
rect 6822 28064 6828 28076
rect 6735 28036 6828 28064
rect 5813 28027 5871 28033
rect 6822 28024 6828 28036
rect 6880 28064 6886 28076
rect 7282 28064 7288 28076
rect 6880 28036 7288 28064
rect 6880 28024 6886 28036
rect 7282 28024 7288 28036
rect 7340 28024 7346 28076
rect 7466 28064 7472 28076
rect 7427 28036 7472 28064
rect 7466 28024 7472 28036
rect 7524 28024 7530 28076
rect 10781 28067 10839 28073
rect 10781 28033 10793 28067
rect 10827 28064 10839 28067
rect 11606 28064 11612 28076
rect 10827 28036 11612 28064
rect 10827 28033 10839 28036
rect 10781 28027 10839 28033
rect 11606 28024 11612 28036
rect 11664 28024 11670 28076
rect 12437 28067 12495 28073
rect 12437 28033 12449 28067
rect 12483 28064 12495 28067
rect 12483 28036 12940 28064
rect 12483 28033 12495 28036
rect 12437 28027 12495 28033
rect 2924 27968 3648 27996
rect 3697 27999 3755 28005
rect 2924 27956 2930 27968
rect 3697 27965 3709 27999
rect 3743 27996 3755 27999
rect 7190 27996 7196 28008
rect 3743 27968 7196 27996
rect 3743 27965 3755 27968
rect 3697 27959 3755 27965
rect 7190 27956 7196 27968
rect 7248 27956 7254 28008
rect 8573 27999 8631 28005
rect 8573 27965 8585 27999
rect 8619 27996 8631 27999
rect 10410 27996 10416 28008
rect 8619 27968 10416 27996
rect 8619 27965 8631 27968
rect 8573 27959 8631 27965
rect 10410 27956 10416 27968
rect 10468 27956 10474 28008
rect 10505 27999 10563 28005
rect 10505 27965 10517 27999
rect 10551 27996 10563 27999
rect 11238 27996 11244 28008
rect 10551 27968 11244 27996
rect 10551 27965 10563 27968
rect 10505 27959 10563 27965
rect 11238 27956 11244 27968
rect 11296 27956 11302 28008
rect 11330 27956 11336 28008
rect 11388 27996 11394 28008
rect 11793 27999 11851 28005
rect 11793 27996 11805 27999
rect 11388 27968 11805 27996
rect 11388 27956 11394 27968
rect 11793 27965 11805 27968
rect 11839 27965 11851 27999
rect 12912 27996 12940 28036
rect 15105 27999 15163 28005
rect 12912 27968 15056 27996
rect 11793 27959 11851 27965
rect 1857 27931 1915 27937
rect 1857 27897 1869 27931
rect 1903 27928 1915 27931
rect 3053 27931 3111 27937
rect 1903 27900 2774 27928
rect 1903 27897 1915 27900
rect 1857 27891 1915 27897
rect 2746 27860 2774 27900
rect 3053 27897 3065 27931
rect 3099 27928 3111 27931
rect 5074 27928 5080 27940
rect 3099 27900 5080 27928
rect 3099 27897 3111 27900
rect 3053 27891 3111 27897
rect 5074 27888 5080 27900
rect 5132 27888 5138 27940
rect 6270 27928 6276 27940
rect 5828 27900 6276 27928
rect 4246 27860 4252 27872
rect 2746 27832 4252 27860
rect 4246 27820 4252 27832
rect 4304 27820 4310 27872
rect 4341 27863 4399 27869
rect 4341 27829 4353 27863
rect 4387 27860 4399 27863
rect 5828 27860 5856 27900
rect 6270 27888 6276 27900
rect 6328 27888 6334 27940
rect 8662 27928 8668 27940
rect 7300 27900 8668 27928
rect 4387 27832 5856 27860
rect 5905 27863 5963 27869
rect 4387 27829 4399 27832
rect 4341 27823 4399 27829
rect 5905 27829 5917 27863
rect 5951 27860 5963 27863
rect 7300 27860 7328 27900
rect 8662 27888 8668 27900
rect 8720 27888 8726 27940
rect 11146 27888 11152 27940
rect 11204 27928 11210 27940
rect 12989 27931 13047 27937
rect 12989 27928 13001 27931
rect 11204 27900 13001 27928
rect 11204 27888 11210 27900
rect 12989 27897 13001 27900
rect 13035 27897 13047 27931
rect 12989 27891 13047 27897
rect 13630 27888 13636 27940
rect 13688 27928 13694 27940
rect 14553 27931 14611 27937
rect 14553 27928 14565 27931
rect 13688 27900 14565 27928
rect 13688 27888 13694 27900
rect 14553 27897 14565 27900
rect 14599 27928 14611 27931
rect 14826 27928 14832 27940
rect 14599 27900 14832 27928
rect 14599 27897 14611 27900
rect 14553 27891 14611 27897
rect 14826 27888 14832 27900
rect 14884 27888 14890 27940
rect 15028 27928 15056 27968
rect 15105 27965 15117 27999
rect 15151 27996 15163 27999
rect 15378 27996 15384 28008
rect 15151 27968 15384 27996
rect 15151 27965 15163 27968
rect 15105 27959 15163 27965
rect 15378 27956 15384 27968
rect 15436 27956 15442 28008
rect 15654 27928 15660 27940
rect 15028 27900 15660 27928
rect 15654 27888 15660 27900
rect 15712 27888 15718 27940
rect 9030 27860 9036 27872
rect 5951 27832 7328 27860
rect 8991 27832 9036 27860
rect 5951 27829 5963 27832
rect 5905 27823 5963 27829
rect 9030 27820 9036 27832
rect 9088 27820 9094 27872
rect 9950 27820 9956 27872
rect 10008 27860 10014 27872
rect 11514 27860 11520 27872
rect 10008 27832 11520 27860
rect 10008 27820 10014 27832
rect 11514 27820 11520 27832
rect 11572 27860 11578 27872
rect 12342 27860 12348 27872
rect 11572 27832 12348 27860
rect 11572 27820 11578 27832
rect 12342 27820 12348 27832
rect 12400 27820 12406 27872
rect 13078 27820 13084 27872
rect 13136 27860 13142 27872
rect 15194 27860 15200 27872
rect 13136 27832 15200 27860
rect 13136 27820 13142 27832
rect 15194 27820 15200 27832
rect 15252 27820 15258 27872
rect 16040 27860 16068 28104
rect 16132 28073 16160 28160
rect 17402 28132 17408 28144
rect 17363 28104 17408 28132
rect 17402 28092 17408 28104
rect 17460 28092 17466 28144
rect 17512 28141 17540 28172
rect 22005 28169 22017 28172
rect 22051 28169 22063 28203
rect 23750 28200 23756 28212
rect 23711 28172 23756 28200
rect 22005 28163 22063 28169
rect 23750 28160 23756 28172
rect 23808 28160 23814 28212
rect 17497 28135 17555 28141
rect 17497 28101 17509 28135
rect 17543 28101 17555 28135
rect 18417 28135 18475 28141
rect 18417 28132 18429 28135
rect 17497 28095 17555 28101
rect 17696 28104 18429 28132
rect 16117 28067 16175 28073
rect 16117 28033 16129 28067
rect 16163 28033 16175 28067
rect 16117 28027 16175 28033
rect 16209 27999 16267 28005
rect 16209 27965 16221 27999
rect 16255 27996 16267 27999
rect 17696 27996 17724 28104
rect 18417 28101 18429 28104
rect 18463 28101 18475 28135
rect 18417 28095 18475 28101
rect 18969 28135 19027 28141
rect 18969 28101 18981 28135
rect 19015 28132 19027 28135
rect 19426 28132 19432 28144
rect 19015 28104 19432 28132
rect 19015 28101 19027 28104
rect 18969 28095 19027 28101
rect 19426 28092 19432 28104
rect 19484 28092 19490 28144
rect 23382 28132 23388 28144
rect 19628 28104 23388 28132
rect 19628 28073 19656 28104
rect 23382 28092 23388 28104
rect 23440 28092 23446 28144
rect 19613 28067 19671 28073
rect 19613 28033 19625 28067
rect 19659 28033 19671 28067
rect 19613 28027 19671 28033
rect 20257 28067 20315 28073
rect 20257 28033 20269 28067
rect 20303 28064 20315 28067
rect 20438 28064 20444 28076
rect 20303 28036 20444 28064
rect 20303 28033 20315 28036
rect 20257 28027 20315 28033
rect 20438 28024 20444 28036
rect 20496 28024 20502 28076
rect 20714 28024 20720 28076
rect 20772 28064 20778 28076
rect 20809 28067 20867 28073
rect 20809 28064 20821 28067
rect 20772 28036 20821 28064
rect 20772 28024 20778 28036
rect 20809 28033 20821 28036
rect 20855 28033 20867 28067
rect 20809 28027 20867 28033
rect 20901 28067 20959 28073
rect 20901 28033 20913 28067
rect 20947 28064 20959 28067
rect 21726 28064 21732 28076
rect 20947 28036 21732 28064
rect 20947 28033 20959 28036
rect 20901 28027 20959 28033
rect 21726 28024 21732 28036
rect 21784 28024 21790 28076
rect 22741 28067 22799 28073
rect 22741 28033 22753 28067
rect 22787 28064 22799 28067
rect 24670 28064 24676 28076
rect 22787 28036 24676 28064
rect 22787 28033 22799 28036
rect 22741 28027 22799 28033
rect 18322 27996 18328 28008
rect 16255 27968 17724 27996
rect 18235 27968 18328 27996
rect 16255 27965 16267 27968
rect 16209 27959 16267 27965
rect 18322 27956 18328 27968
rect 18380 27996 18386 28008
rect 18506 27996 18512 28008
rect 18380 27968 18512 27996
rect 18380 27956 18386 27968
rect 18506 27956 18512 27968
rect 18564 27956 18570 28008
rect 18598 27956 18604 28008
rect 18656 27996 18662 28008
rect 21358 27996 21364 28008
rect 18656 27968 21364 27996
rect 18656 27956 18662 27968
rect 21358 27956 21364 27968
rect 21416 27956 21422 28008
rect 16482 27888 16488 27940
rect 16540 27928 16546 27940
rect 16945 27931 17003 27937
rect 16945 27928 16957 27931
rect 16540 27900 16957 27928
rect 16540 27888 16546 27900
rect 16945 27897 16957 27900
rect 16991 27897 17003 27931
rect 18874 27928 18880 27940
rect 16945 27891 17003 27897
rect 17512 27900 18880 27928
rect 17512 27860 17540 27900
rect 18874 27888 18880 27900
rect 18932 27888 18938 27940
rect 20165 27931 20223 27937
rect 20165 27928 20177 27931
rect 18984 27900 20177 27928
rect 16040 27832 17540 27860
rect 17586 27820 17592 27872
rect 17644 27860 17650 27872
rect 18984 27860 19012 27900
rect 20165 27897 20177 27900
rect 20211 27897 20223 27931
rect 20165 27891 20223 27897
rect 20438 27888 20444 27940
rect 20496 27928 20502 27940
rect 22756 27928 22784 28027
rect 24670 28024 24676 28036
rect 24728 28024 24734 28076
rect 20496 27900 22784 27928
rect 23293 27931 23351 27937
rect 20496 27888 20502 27900
rect 23293 27897 23305 27931
rect 23339 27928 23351 27931
rect 23382 27928 23388 27940
rect 23339 27900 23388 27928
rect 23339 27897 23351 27900
rect 23293 27891 23351 27897
rect 23382 27888 23388 27900
rect 23440 27928 23446 27940
rect 37734 27928 37740 27940
rect 23440 27900 37740 27928
rect 23440 27888 23446 27900
rect 37734 27888 37740 27900
rect 37792 27888 37798 27940
rect 19518 27860 19524 27872
rect 17644 27832 19012 27860
rect 19479 27832 19524 27860
rect 17644 27820 17650 27832
rect 19518 27820 19524 27832
rect 19576 27820 19582 27872
rect 19978 27820 19984 27872
rect 20036 27860 20042 27872
rect 22554 27860 22560 27872
rect 20036 27832 22560 27860
rect 20036 27820 20042 27832
rect 22554 27820 22560 27832
rect 22612 27820 22618 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 3418 27616 3424 27668
rect 3476 27656 3482 27668
rect 10134 27656 10140 27668
rect 3476 27628 10140 27656
rect 3476 27616 3482 27628
rect 10134 27616 10140 27628
rect 10192 27616 10198 27668
rect 10410 27616 10416 27668
rect 10468 27656 10474 27668
rect 12986 27656 12992 27668
rect 10468 27628 12992 27656
rect 10468 27616 10474 27628
rect 12986 27616 12992 27628
rect 13044 27656 13050 27668
rect 13044 27628 15148 27656
rect 13044 27616 13050 27628
rect 2133 27591 2191 27597
rect 2133 27557 2145 27591
rect 2179 27588 2191 27591
rect 3050 27588 3056 27600
rect 2179 27560 3056 27588
rect 2179 27557 2191 27560
rect 2133 27551 2191 27557
rect 3050 27548 3056 27560
rect 3108 27548 3114 27600
rect 4062 27588 4068 27600
rect 4023 27560 4068 27588
rect 4062 27548 4068 27560
rect 4120 27548 4126 27600
rect 4709 27591 4767 27597
rect 4709 27557 4721 27591
rect 4755 27588 4767 27591
rect 5718 27588 5724 27600
rect 4755 27560 5724 27588
rect 4755 27557 4767 27560
rect 4709 27551 4767 27557
rect 5718 27548 5724 27560
rect 5776 27548 5782 27600
rect 6086 27548 6092 27600
rect 6144 27588 6150 27600
rect 6825 27591 6883 27597
rect 6825 27588 6837 27591
rect 6144 27560 6837 27588
rect 6144 27548 6150 27560
rect 6825 27557 6837 27560
rect 6871 27557 6883 27591
rect 6825 27551 6883 27557
rect 9401 27591 9459 27597
rect 9401 27557 9413 27591
rect 9447 27588 9459 27591
rect 10042 27588 10048 27600
rect 9447 27560 10048 27588
rect 9447 27557 9459 27560
rect 9401 27551 9459 27557
rect 2682 27480 2688 27532
rect 2740 27520 2746 27532
rect 2777 27523 2835 27529
rect 2777 27520 2789 27523
rect 2740 27492 2789 27520
rect 2740 27480 2746 27492
rect 2777 27489 2789 27492
rect 2823 27489 2835 27523
rect 2777 27483 2835 27489
rect 3786 27480 3792 27532
rect 3844 27520 3850 27532
rect 5258 27520 5264 27532
rect 3844 27492 5264 27520
rect 3844 27480 3850 27492
rect 1670 27412 1676 27464
rect 1728 27452 1734 27464
rect 2041 27455 2099 27461
rect 2041 27452 2053 27455
rect 1728 27424 2053 27452
rect 1728 27412 1734 27424
rect 2041 27421 2053 27424
rect 2087 27452 2099 27455
rect 2869 27455 2927 27461
rect 2869 27452 2881 27455
rect 2087 27424 2881 27452
rect 2087 27421 2099 27424
rect 2041 27415 2099 27421
rect 2869 27421 2881 27424
rect 2915 27421 2927 27455
rect 2869 27415 2927 27421
rect 3973 27455 4031 27461
rect 3973 27421 3985 27455
rect 4019 27452 4031 27455
rect 4338 27452 4344 27464
rect 4019 27424 4344 27452
rect 4019 27421 4031 27424
rect 3973 27415 4031 27421
rect 2682 27344 2688 27396
rect 2740 27384 2746 27396
rect 2884 27384 2912 27415
rect 4338 27412 4344 27424
rect 4396 27412 4402 27464
rect 4632 27461 4660 27492
rect 5258 27480 5264 27492
rect 5316 27480 5322 27532
rect 4617 27455 4675 27461
rect 4617 27421 4629 27455
rect 4663 27421 4675 27455
rect 6840 27452 6868 27551
rect 10042 27548 10048 27560
rect 10100 27548 10106 27600
rect 12158 27588 12164 27600
rect 10152 27560 12164 27588
rect 8021 27523 8079 27529
rect 8021 27489 8033 27523
rect 8067 27520 8079 27523
rect 9858 27520 9864 27532
rect 8067 27492 9864 27520
rect 8067 27489 8079 27492
rect 8021 27483 8079 27489
rect 9858 27480 9864 27492
rect 9916 27480 9922 27532
rect 10152 27520 10180 27560
rect 12158 27548 12164 27560
rect 12216 27588 12222 27600
rect 13633 27591 13691 27597
rect 12216 27560 13584 27588
rect 12216 27548 12222 27560
rect 9968 27492 10180 27520
rect 10321 27523 10379 27529
rect 8110 27452 8116 27464
rect 6840 27424 8116 27452
rect 4617 27415 4675 27421
rect 8110 27412 8116 27424
rect 8168 27452 8174 27464
rect 9309 27455 9367 27461
rect 9309 27452 9321 27455
rect 8168 27424 9321 27452
rect 8168 27412 8174 27424
rect 9309 27421 9321 27424
rect 9355 27421 9367 27455
rect 9309 27415 9367 27421
rect 3234 27384 3240 27396
rect 2740 27356 3240 27384
rect 2740 27344 2746 27356
rect 3234 27344 3240 27356
rect 3292 27384 3298 27396
rect 3421 27387 3479 27393
rect 3421 27384 3433 27387
rect 3292 27356 3433 27384
rect 3292 27344 3298 27356
rect 3421 27353 3433 27356
rect 3467 27384 3479 27387
rect 3786 27384 3792 27396
rect 3467 27356 3792 27384
rect 3467 27353 3479 27356
rect 3421 27347 3479 27353
rect 3786 27344 3792 27356
rect 3844 27384 3850 27396
rect 6822 27384 6828 27396
rect 3844 27356 6828 27384
rect 3844 27344 3850 27356
rect 6822 27344 6828 27356
rect 6880 27344 6886 27396
rect 8573 27387 8631 27393
rect 8573 27353 8585 27387
rect 8619 27384 8631 27387
rect 8754 27384 8760 27396
rect 8619 27356 8760 27384
rect 8619 27353 8631 27356
rect 8573 27347 8631 27353
rect 8754 27344 8760 27356
rect 8812 27384 8818 27396
rect 9968 27384 9996 27492
rect 10321 27489 10333 27523
rect 10367 27520 10379 27523
rect 11422 27520 11428 27532
rect 10367 27492 11428 27520
rect 10367 27489 10379 27492
rect 10321 27483 10379 27489
rect 11422 27480 11428 27492
rect 11480 27480 11486 27532
rect 12434 27480 12440 27532
rect 12492 27520 12498 27532
rect 12802 27520 12808 27532
rect 12492 27492 12808 27520
rect 12492 27480 12498 27492
rect 12802 27480 12808 27492
rect 12860 27480 12866 27532
rect 12894 27452 12900 27464
rect 12855 27424 12900 27452
rect 12894 27412 12900 27424
rect 12952 27412 12958 27464
rect 13556 27461 13584 27560
rect 13633 27557 13645 27591
rect 13679 27588 13691 27591
rect 14550 27588 14556 27600
rect 13679 27560 14556 27588
rect 13679 27557 13691 27560
rect 13633 27551 13691 27557
rect 14550 27548 14556 27560
rect 14608 27548 14614 27600
rect 15120 27588 15148 27628
rect 16850 27616 16856 27668
rect 16908 27656 16914 27668
rect 20346 27656 20352 27668
rect 16908 27628 20352 27656
rect 16908 27616 16914 27628
rect 20346 27616 20352 27628
rect 20404 27616 20410 27668
rect 15378 27588 15384 27600
rect 15120 27560 15384 27588
rect 15378 27548 15384 27560
rect 15436 27548 15442 27600
rect 16390 27588 16396 27600
rect 16351 27560 16396 27588
rect 16390 27548 16396 27560
rect 16448 27548 16454 27600
rect 18782 27548 18788 27600
rect 18840 27588 18846 27600
rect 18840 27560 21220 27588
rect 18840 27548 18846 27560
rect 14366 27520 14372 27532
rect 14279 27492 14372 27520
rect 14366 27480 14372 27492
rect 14424 27520 14430 27532
rect 17586 27520 17592 27532
rect 14424 27492 16436 27520
rect 17547 27492 17592 27520
rect 14424 27480 14430 27492
rect 13541 27455 13599 27461
rect 13541 27421 13553 27455
rect 13587 27452 13599 27455
rect 14182 27452 14188 27464
rect 13587 27424 14188 27452
rect 13587 27421 13599 27424
rect 13541 27415 13599 27421
rect 14182 27412 14188 27424
rect 14240 27412 14246 27464
rect 16114 27412 16120 27464
rect 16172 27452 16178 27464
rect 16301 27455 16359 27461
rect 16301 27452 16313 27455
rect 16172 27424 16313 27452
rect 16172 27412 16178 27424
rect 16301 27421 16313 27424
rect 16347 27421 16359 27455
rect 16301 27415 16359 27421
rect 16408 27396 16436 27492
rect 17586 27480 17592 27492
rect 17644 27480 17650 27532
rect 19518 27480 19524 27532
rect 19576 27520 19582 27532
rect 20533 27523 20591 27529
rect 20533 27520 20545 27523
rect 19576 27492 20545 27520
rect 19576 27480 19582 27492
rect 20533 27489 20545 27492
rect 20579 27489 20591 27523
rect 20533 27483 20591 27489
rect 20622 27480 20628 27532
rect 20680 27520 20686 27532
rect 20809 27523 20867 27529
rect 20809 27520 20821 27523
rect 20680 27492 20821 27520
rect 20680 27480 20686 27492
rect 20809 27489 20821 27492
rect 20855 27489 20867 27523
rect 20809 27483 20867 27489
rect 19429 27455 19487 27461
rect 19429 27421 19441 27455
rect 19475 27452 19487 27455
rect 19978 27452 19984 27464
rect 19475 27424 19984 27452
rect 19475 27421 19487 27424
rect 19429 27415 19487 27421
rect 19978 27412 19984 27424
rect 20036 27412 20042 27464
rect 10502 27384 10508 27396
rect 8812 27356 9996 27384
rect 10463 27356 10508 27384
rect 8812 27344 8818 27356
rect 10502 27344 10508 27356
rect 10560 27344 10566 27396
rect 10597 27387 10655 27393
rect 10597 27353 10609 27387
rect 10643 27384 10655 27387
rect 11514 27384 11520 27396
rect 10643 27356 11520 27384
rect 10643 27353 10655 27356
rect 10597 27347 10655 27353
rect 11514 27344 11520 27356
rect 11572 27344 11578 27396
rect 11701 27387 11759 27393
rect 11701 27353 11713 27387
rect 11747 27353 11759 27387
rect 11701 27347 11759 27353
rect 11793 27387 11851 27393
rect 11793 27353 11805 27387
rect 11839 27384 11851 27387
rect 13078 27384 13084 27396
rect 11839 27356 13084 27384
rect 11839 27353 11851 27356
rect 11793 27347 11851 27353
rect 5534 27276 5540 27328
rect 5592 27316 5598 27328
rect 5721 27319 5779 27325
rect 5721 27316 5733 27319
rect 5592 27288 5733 27316
rect 5592 27276 5598 27288
rect 5721 27285 5733 27288
rect 5767 27285 5779 27319
rect 5721 27279 5779 27285
rect 6365 27319 6423 27325
rect 6365 27285 6377 27319
rect 6411 27316 6423 27319
rect 6638 27316 6644 27328
rect 6411 27288 6644 27316
rect 6411 27285 6423 27288
rect 6365 27279 6423 27285
rect 6638 27276 6644 27288
rect 6696 27276 6702 27328
rect 6914 27276 6920 27328
rect 6972 27316 6978 27328
rect 7374 27316 7380 27328
rect 6972 27288 7380 27316
rect 6972 27276 6978 27288
rect 7374 27276 7380 27288
rect 7432 27276 7438 27328
rect 7469 27319 7527 27325
rect 7469 27285 7481 27319
rect 7515 27316 7527 27319
rect 9122 27316 9128 27328
rect 7515 27288 9128 27316
rect 7515 27285 7527 27288
rect 7469 27279 7527 27285
rect 9122 27276 9128 27288
rect 9180 27276 9186 27328
rect 9766 27276 9772 27328
rect 9824 27316 9830 27328
rect 11716 27316 11744 27347
rect 13078 27344 13084 27356
rect 13136 27384 13142 27396
rect 13262 27384 13268 27396
rect 13136 27356 13268 27384
rect 13136 27344 13142 27356
rect 13262 27344 13268 27356
rect 13320 27344 13326 27396
rect 13354 27344 13360 27396
rect 13412 27384 13418 27396
rect 14461 27387 14519 27393
rect 13412 27356 14320 27384
rect 13412 27344 13418 27356
rect 9824 27288 11744 27316
rect 12437 27319 12495 27325
rect 9824 27276 9830 27288
rect 12437 27285 12449 27319
rect 12483 27316 12495 27319
rect 12526 27316 12532 27328
rect 12483 27288 12532 27316
rect 12483 27285 12495 27288
rect 12437 27279 12495 27285
rect 12526 27276 12532 27288
rect 12584 27316 12590 27328
rect 12710 27316 12716 27328
rect 12584 27288 12716 27316
rect 12584 27276 12590 27288
rect 12710 27276 12716 27288
rect 12768 27276 12774 27328
rect 12989 27319 13047 27325
rect 12989 27285 13001 27319
rect 13035 27316 13047 27319
rect 13446 27316 13452 27328
rect 13035 27288 13452 27316
rect 13035 27285 13047 27288
rect 12989 27279 13047 27285
rect 13446 27276 13452 27288
rect 13504 27276 13510 27328
rect 14292 27316 14320 27356
rect 14461 27353 14473 27387
rect 14507 27353 14519 27387
rect 14461 27347 14519 27353
rect 15381 27387 15439 27393
rect 15381 27353 15393 27387
rect 15427 27384 15439 27387
rect 15562 27384 15568 27396
rect 15427 27356 15568 27384
rect 15427 27353 15439 27356
rect 15381 27347 15439 27353
rect 14476 27316 14504 27347
rect 15562 27344 15568 27356
rect 15620 27344 15626 27396
rect 16390 27344 16396 27396
rect 16448 27384 16454 27396
rect 16945 27387 17003 27393
rect 16945 27384 16957 27387
rect 16448 27356 16957 27384
rect 16448 27344 16454 27356
rect 16945 27353 16957 27356
rect 16991 27353 17003 27387
rect 17494 27384 17500 27396
rect 17455 27356 17500 27384
rect 16945 27347 17003 27353
rect 17494 27344 17500 27356
rect 17552 27344 17558 27396
rect 18141 27387 18199 27393
rect 18141 27353 18153 27387
rect 18187 27353 18199 27387
rect 18690 27384 18696 27396
rect 18651 27356 18696 27384
rect 18141 27347 18199 27353
rect 14292 27288 14504 27316
rect 15286 27276 15292 27328
rect 15344 27316 15350 27328
rect 18156 27316 18184 27347
rect 18690 27344 18696 27356
rect 18748 27344 18754 27396
rect 18785 27387 18843 27393
rect 18785 27353 18797 27387
rect 18831 27384 18843 27387
rect 20530 27384 20536 27396
rect 18831 27356 20536 27384
rect 18831 27353 18843 27356
rect 18785 27347 18843 27353
rect 20530 27344 20536 27356
rect 20588 27344 20594 27396
rect 20625 27387 20683 27393
rect 20625 27353 20637 27387
rect 20671 27384 20683 27387
rect 20990 27384 20996 27396
rect 20671 27356 20996 27384
rect 20671 27353 20683 27356
rect 20625 27347 20683 27353
rect 20990 27344 20996 27356
rect 21048 27344 21054 27396
rect 21192 27384 21220 27560
rect 21266 27548 21272 27600
rect 21324 27588 21330 27600
rect 22002 27588 22008 27600
rect 21324 27560 22008 27588
rect 21324 27548 21330 27560
rect 22002 27548 22008 27560
rect 22060 27588 22066 27600
rect 22833 27591 22891 27597
rect 22833 27588 22845 27591
rect 22060 27560 22845 27588
rect 22060 27548 22066 27560
rect 22833 27557 22845 27560
rect 22879 27557 22891 27591
rect 22833 27551 22891 27557
rect 21634 27412 21640 27464
rect 21692 27452 21698 27464
rect 23937 27455 23995 27461
rect 23937 27452 23949 27455
rect 21692 27424 23949 27452
rect 21692 27412 21698 27424
rect 23937 27421 23949 27424
rect 23983 27421 23995 27455
rect 23937 27415 23995 27421
rect 22373 27387 22431 27393
rect 22373 27384 22385 27387
rect 21192 27356 22385 27384
rect 22373 27353 22385 27356
rect 22419 27384 22431 27387
rect 34514 27384 34520 27396
rect 22419 27356 34520 27384
rect 22419 27353 22431 27356
rect 22373 27347 22431 27353
rect 34514 27344 34520 27356
rect 34572 27344 34578 27396
rect 15344 27288 18184 27316
rect 15344 27276 15350 27288
rect 19334 27276 19340 27328
rect 19392 27316 19398 27328
rect 19521 27319 19579 27325
rect 19521 27316 19533 27319
rect 19392 27288 19533 27316
rect 19392 27276 19398 27288
rect 19521 27285 19533 27288
rect 19567 27285 19579 27319
rect 19521 27279 19579 27285
rect 19978 27276 19984 27328
rect 20036 27316 20042 27328
rect 21266 27316 21272 27328
rect 20036 27288 21272 27316
rect 20036 27276 20042 27288
rect 21266 27276 21272 27288
rect 21324 27276 21330 27328
rect 21818 27316 21824 27328
rect 21779 27288 21824 27316
rect 21818 27276 21824 27288
rect 21876 27276 21882 27328
rect 23382 27316 23388 27328
rect 23343 27288 23388 27316
rect 23382 27276 23388 27288
rect 23440 27276 23446 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 2222 27072 2228 27124
rect 2280 27112 2286 27124
rect 2409 27115 2467 27121
rect 2409 27112 2421 27115
rect 2280 27084 2421 27112
rect 2280 27072 2286 27084
rect 2409 27081 2421 27084
rect 2455 27081 2467 27115
rect 3694 27112 3700 27124
rect 3655 27084 3700 27112
rect 2409 27075 2467 27081
rect 3694 27072 3700 27084
rect 3752 27072 3758 27124
rect 6917 27115 6975 27121
rect 6917 27081 6929 27115
rect 6963 27112 6975 27115
rect 7098 27112 7104 27124
rect 6963 27084 7104 27112
rect 6963 27081 6975 27084
rect 6917 27075 6975 27081
rect 7098 27072 7104 27084
rect 7156 27112 7162 27124
rect 7558 27112 7564 27124
rect 7156 27084 7564 27112
rect 7156 27072 7162 27084
rect 7558 27072 7564 27084
rect 7616 27072 7622 27124
rect 8021 27115 8079 27121
rect 8021 27081 8033 27115
rect 8067 27112 8079 27115
rect 10502 27112 10508 27124
rect 8067 27084 10508 27112
rect 8067 27081 8079 27084
rect 8021 27075 8079 27081
rect 10502 27072 10508 27084
rect 10560 27072 10566 27124
rect 11057 27115 11115 27121
rect 11057 27081 11069 27115
rect 11103 27112 11115 27115
rect 12066 27112 12072 27124
rect 11103 27084 12072 27112
rect 11103 27081 11115 27084
rect 11057 27075 11115 27081
rect 12066 27072 12072 27084
rect 12124 27072 12130 27124
rect 15102 27112 15108 27124
rect 13832 27084 15108 27112
rect 3053 27047 3111 27053
rect 3053 27013 3065 27047
rect 3099 27044 3111 27047
rect 8478 27044 8484 27056
rect 3099 27016 8484 27044
rect 3099 27013 3111 27016
rect 3053 27007 3111 27013
rect 8478 27004 8484 27016
rect 8536 27004 8542 27056
rect 8570 27004 8576 27056
rect 8628 27004 8634 27056
rect 9490 27044 9496 27056
rect 9451 27016 9496 27044
rect 9490 27004 9496 27016
rect 9548 27004 9554 27056
rect 9585 27047 9643 27053
rect 9585 27013 9597 27047
rect 9631 27044 9643 27047
rect 11146 27044 11152 27056
rect 9631 27016 11152 27044
rect 9631 27013 9643 27016
rect 9585 27007 9643 27013
rect 11146 27004 11152 27016
rect 11204 27004 11210 27056
rect 12434 27004 12440 27056
rect 12492 27044 12498 27056
rect 13722 27044 13728 27056
rect 12492 27016 12537 27044
rect 13683 27016 13728 27044
rect 12492 27004 12498 27016
rect 13722 27004 13728 27016
rect 13780 27004 13786 27056
rect 13832 27053 13860 27084
rect 15102 27072 15108 27084
rect 15160 27112 15166 27124
rect 20714 27112 20720 27124
rect 15160 27084 15700 27112
rect 15160 27072 15166 27084
rect 13817 27047 13875 27053
rect 13817 27013 13829 27047
rect 13863 27013 13875 27047
rect 14550 27044 14556 27056
rect 14511 27016 14556 27044
rect 13817 27007 13875 27013
rect 14550 27004 14556 27016
rect 14608 27004 14614 27056
rect 15672 27053 15700 27084
rect 18984 27084 20720 27112
rect 15657 27047 15715 27053
rect 15657 27013 15669 27047
rect 15703 27013 15715 27047
rect 15657 27007 15715 27013
rect 15749 27047 15807 27053
rect 15749 27013 15761 27047
rect 15795 27044 15807 27047
rect 16942 27044 16948 27056
rect 15795 27016 16948 27044
rect 15795 27013 15807 27016
rect 15749 27007 15807 27013
rect 16942 27004 16948 27016
rect 17000 27004 17006 27056
rect 17589 27047 17647 27053
rect 17589 27013 17601 27047
rect 17635 27044 17647 27047
rect 17862 27044 17868 27056
rect 17635 27016 17868 27044
rect 17635 27013 17647 27016
rect 17589 27007 17647 27013
rect 17862 27004 17868 27016
rect 17920 27004 17926 27056
rect 18984 27053 19012 27084
rect 20714 27072 20720 27084
rect 20772 27072 20778 27124
rect 18969 27047 19027 27053
rect 18969 27013 18981 27047
rect 19015 27013 19027 27047
rect 18969 27007 19027 27013
rect 19334 27004 19340 27056
rect 19392 27044 19398 27056
rect 19794 27044 19800 27056
rect 19392 27016 19800 27044
rect 19392 27004 19398 27016
rect 19794 27004 19800 27016
rect 19852 27004 19858 27056
rect 20165 27047 20223 27053
rect 20165 27013 20177 27047
rect 20211 27044 20223 27047
rect 21269 27047 21327 27053
rect 21269 27044 21281 27047
rect 20211 27016 21281 27044
rect 20211 27013 20223 27016
rect 20165 27007 20223 27013
rect 21269 27013 21281 27016
rect 21315 27013 21327 27047
rect 21269 27007 21327 27013
rect 22557 27047 22615 27053
rect 22557 27013 22569 27047
rect 22603 27044 22615 27047
rect 22646 27044 22652 27056
rect 22603 27016 22652 27044
rect 22603 27013 22615 27016
rect 22557 27007 22615 27013
rect 22646 27004 22652 27016
rect 22704 27004 22710 27056
rect 23290 27004 23296 27056
rect 23348 27044 23354 27056
rect 23385 27047 23443 27053
rect 23385 27044 23397 27047
rect 23348 27016 23397 27044
rect 23348 27004 23354 27016
rect 23385 27013 23397 27016
rect 23431 27013 23443 27047
rect 23385 27007 23443 27013
rect 1857 26979 1915 26985
rect 1857 26945 1869 26979
rect 1903 26945 1915 26979
rect 1857 26939 1915 26945
rect 2317 26979 2375 26985
rect 2317 26945 2329 26979
rect 2363 26976 2375 26979
rect 2866 26976 2872 26988
rect 2363 26948 2872 26976
rect 2363 26945 2375 26948
rect 2317 26939 2375 26945
rect 1872 26840 1900 26939
rect 2866 26936 2872 26948
rect 2924 26976 2930 26988
rect 2961 26979 3019 26985
rect 2961 26976 2973 26979
rect 2924 26948 2973 26976
rect 2924 26936 2930 26948
rect 2961 26945 2973 26948
rect 3007 26945 3019 26979
rect 3786 26976 3792 26988
rect 3747 26948 3792 26976
rect 2961 26939 3019 26945
rect 3786 26936 3792 26948
rect 3844 26936 3850 26988
rect 7929 26979 7987 26985
rect 7929 26945 7941 26979
rect 7975 26976 7987 26979
rect 8588 26976 8616 27004
rect 7975 26948 8616 26976
rect 7975 26945 7987 26948
rect 7929 26939 7987 26945
rect 10226 26936 10232 26988
rect 10284 26976 10290 26988
rect 10321 26979 10379 26985
rect 10321 26976 10333 26979
rect 10284 26948 10333 26976
rect 10284 26936 10290 26948
rect 10321 26945 10333 26948
rect 10367 26945 10379 26979
rect 10962 26976 10968 26988
rect 10923 26948 10968 26976
rect 10321 26939 10379 26945
rect 10962 26936 10968 26948
rect 11020 26936 11026 26988
rect 16301 26979 16359 26985
rect 16301 26945 16313 26979
rect 16347 26976 16359 26979
rect 16390 26976 16396 26988
rect 16347 26948 16396 26976
rect 16347 26945 16359 26948
rect 16301 26939 16359 26945
rect 16390 26936 16396 26948
rect 16448 26936 16454 26988
rect 21358 26976 21364 26988
rect 21319 26948 21364 26976
rect 21358 26936 21364 26948
rect 21416 26936 21422 26988
rect 22005 26979 22063 26985
rect 22005 26976 22017 26979
rect 21836 26948 22017 26976
rect 5074 26868 5080 26920
rect 5132 26908 5138 26920
rect 8018 26908 8024 26920
rect 5132 26880 8024 26908
rect 5132 26868 5138 26880
rect 8018 26868 8024 26880
rect 8076 26868 8082 26920
rect 9309 26911 9367 26917
rect 9309 26877 9321 26911
rect 9355 26908 9367 26911
rect 9858 26908 9864 26920
rect 9355 26880 9864 26908
rect 9355 26877 9367 26880
rect 9309 26871 9367 26877
rect 9858 26868 9864 26880
rect 9916 26868 9922 26920
rect 11146 26868 11152 26920
rect 11204 26908 11210 26920
rect 11885 26911 11943 26917
rect 11885 26908 11897 26911
rect 11204 26880 11897 26908
rect 11204 26868 11210 26880
rect 11885 26877 11897 26880
rect 11931 26877 11943 26911
rect 11885 26871 11943 26877
rect 12529 26911 12587 26917
rect 12529 26877 12541 26911
rect 12575 26908 12587 26911
rect 14274 26908 14280 26920
rect 12575 26880 14280 26908
rect 12575 26877 12587 26880
rect 12529 26871 12587 26877
rect 14274 26868 14280 26880
rect 14332 26868 14338 26920
rect 14461 26911 14519 26917
rect 14461 26877 14473 26911
rect 14507 26877 14519 26911
rect 14461 26871 14519 26877
rect 6822 26840 6828 26852
rect 1872 26812 6828 26840
rect 6822 26800 6828 26812
rect 6880 26800 6886 26852
rect 7466 26840 7472 26852
rect 7427 26812 7472 26840
rect 7466 26800 7472 26812
rect 7524 26800 7530 26852
rect 9048 26812 12020 26840
rect 1670 26772 1676 26784
rect 1631 26744 1676 26772
rect 1670 26732 1676 26744
rect 1728 26732 1734 26784
rect 4338 26772 4344 26784
rect 4251 26744 4344 26772
rect 4338 26732 4344 26744
rect 4396 26772 4402 26784
rect 4614 26772 4620 26784
rect 4396 26744 4620 26772
rect 4396 26732 4402 26744
rect 4614 26732 4620 26744
rect 4672 26732 4678 26784
rect 4893 26775 4951 26781
rect 4893 26741 4905 26775
rect 4939 26772 4951 26775
rect 5074 26772 5080 26784
rect 4939 26744 5080 26772
rect 4939 26741 4951 26744
rect 4893 26735 4951 26741
rect 5074 26732 5080 26744
rect 5132 26732 5138 26784
rect 5350 26772 5356 26784
rect 5311 26744 5356 26772
rect 5350 26732 5356 26744
rect 5408 26732 5414 26784
rect 5534 26732 5540 26784
rect 5592 26772 5598 26784
rect 5905 26775 5963 26781
rect 5905 26772 5917 26775
rect 5592 26744 5917 26772
rect 5592 26732 5598 26744
rect 5905 26741 5917 26744
rect 5951 26741 5963 26775
rect 5905 26735 5963 26741
rect 5994 26732 6000 26784
rect 6052 26772 6058 26784
rect 9048 26772 9076 26812
rect 6052 26744 9076 26772
rect 6052 26732 6058 26744
rect 9122 26732 9128 26784
rect 9180 26772 9186 26784
rect 9950 26772 9956 26784
rect 9180 26744 9956 26772
rect 9180 26732 9186 26744
rect 9950 26732 9956 26744
rect 10008 26732 10014 26784
rect 10413 26775 10471 26781
rect 10413 26741 10425 26775
rect 10459 26772 10471 26775
rect 10686 26772 10692 26784
rect 10459 26744 10692 26772
rect 10459 26741 10471 26744
rect 10413 26735 10471 26741
rect 10686 26732 10692 26744
rect 10744 26732 10750 26784
rect 11992 26772 12020 26812
rect 12066 26800 12072 26852
rect 12124 26840 12130 26852
rect 13265 26843 13323 26849
rect 13265 26840 13277 26843
rect 12124 26812 13277 26840
rect 12124 26800 12130 26812
rect 13265 26809 13277 26812
rect 13311 26809 13323 26843
rect 13265 26803 13323 26809
rect 12526 26772 12532 26784
rect 11992 26744 12532 26772
rect 12526 26732 12532 26744
rect 12584 26732 12590 26784
rect 13078 26732 13084 26784
rect 13136 26772 13142 26784
rect 14476 26772 14504 26871
rect 16114 26868 16120 26920
rect 16172 26908 16178 26920
rect 16172 26880 17264 26908
rect 16172 26868 16178 26880
rect 15013 26843 15071 26849
rect 15013 26809 15025 26843
rect 15059 26840 15071 26843
rect 15059 26812 15792 26840
rect 15059 26809 15071 26812
rect 15013 26803 15071 26809
rect 13136 26744 14504 26772
rect 13136 26732 13142 26744
rect 14734 26732 14740 26784
rect 14792 26772 14798 26784
rect 15286 26772 15292 26784
rect 14792 26744 15292 26772
rect 14792 26732 14798 26744
rect 15286 26732 15292 26744
rect 15344 26732 15350 26784
rect 15764 26772 15792 26812
rect 15838 26800 15844 26852
rect 15896 26840 15902 26852
rect 17129 26843 17187 26849
rect 17129 26840 17141 26843
rect 15896 26812 17141 26840
rect 15896 26800 15902 26812
rect 17129 26809 17141 26812
rect 17175 26809 17187 26843
rect 17236 26840 17264 26880
rect 17586 26868 17592 26920
rect 17644 26908 17650 26920
rect 17681 26911 17739 26917
rect 17681 26908 17693 26911
rect 17644 26880 17693 26908
rect 17644 26868 17650 26880
rect 17681 26877 17693 26880
rect 17727 26877 17739 26911
rect 18414 26908 18420 26920
rect 18375 26880 18420 26908
rect 17681 26871 17739 26877
rect 18414 26868 18420 26880
rect 18472 26908 18478 26920
rect 18966 26908 18972 26920
rect 18472 26880 18972 26908
rect 18472 26868 18478 26880
rect 18966 26868 18972 26880
rect 19024 26868 19030 26920
rect 19061 26911 19119 26917
rect 19061 26877 19073 26911
rect 19107 26908 19119 26911
rect 19426 26908 19432 26920
rect 19107 26880 19432 26908
rect 19107 26877 19119 26880
rect 19061 26871 19119 26877
rect 19426 26868 19432 26880
rect 19484 26868 19490 26920
rect 20254 26908 20260 26920
rect 19628 26880 19840 26908
rect 20215 26880 20260 26908
rect 19628 26840 19656 26880
rect 17236 26812 19656 26840
rect 19705 26843 19763 26849
rect 17129 26803 17187 26809
rect 19705 26809 19717 26843
rect 19751 26809 19763 26843
rect 19812 26840 19840 26880
rect 20254 26868 20260 26880
rect 20312 26868 20318 26920
rect 20622 26868 20628 26920
rect 20680 26908 20686 26920
rect 21836 26908 21864 26948
rect 22005 26945 22017 26948
rect 22051 26945 22063 26979
rect 22005 26939 22063 26945
rect 36630 26936 36636 26988
rect 36688 26976 36694 26988
rect 38013 26979 38071 26985
rect 38013 26976 38025 26979
rect 36688 26948 38025 26976
rect 36688 26936 36694 26948
rect 38013 26945 38025 26948
rect 38059 26945 38071 26979
rect 38013 26939 38071 26945
rect 22649 26911 22707 26917
rect 22649 26908 22661 26911
rect 20680 26880 21864 26908
rect 22066 26880 22661 26908
rect 20680 26868 20686 26880
rect 21634 26840 21640 26852
rect 19812 26812 21640 26840
rect 19705 26803 19763 26809
rect 19518 26772 19524 26784
rect 15764 26744 19524 26772
rect 19518 26732 19524 26744
rect 19576 26772 19582 26784
rect 19720 26772 19748 26803
rect 21634 26800 21640 26812
rect 21692 26800 21698 26852
rect 21818 26800 21824 26852
rect 21876 26840 21882 26852
rect 22066 26840 22094 26880
rect 22649 26877 22661 26880
rect 22695 26877 22707 26911
rect 22649 26871 22707 26877
rect 23293 26911 23351 26917
rect 23293 26877 23305 26911
rect 23339 26877 23351 26911
rect 23566 26908 23572 26920
rect 23527 26880 23572 26908
rect 23293 26871 23351 26877
rect 21876 26812 22094 26840
rect 21876 26800 21882 26812
rect 22462 26800 22468 26852
rect 22520 26840 22526 26852
rect 23308 26840 23336 26871
rect 23566 26868 23572 26880
rect 23624 26868 23630 26920
rect 22520 26812 23336 26840
rect 22520 26800 22526 26812
rect 19576 26744 19748 26772
rect 19576 26732 19582 26744
rect 20254 26732 20260 26784
rect 20312 26772 20318 26784
rect 29822 26772 29828 26784
rect 20312 26744 29828 26772
rect 20312 26732 20318 26744
rect 29822 26732 29828 26744
rect 29880 26732 29886 26784
rect 38194 26772 38200 26784
rect 38155 26744 38200 26772
rect 38194 26732 38200 26744
rect 38252 26732 38258 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 1949 26571 2007 26577
rect 1949 26537 1961 26571
rect 1995 26568 2007 26571
rect 2038 26568 2044 26580
rect 1995 26540 2044 26568
rect 1995 26537 2007 26540
rect 1949 26531 2007 26537
rect 2038 26528 2044 26540
rect 2096 26528 2102 26580
rect 2130 26528 2136 26580
rect 2188 26568 2194 26580
rect 2593 26571 2651 26577
rect 2593 26568 2605 26571
rect 2188 26540 2605 26568
rect 2188 26528 2194 26540
rect 2593 26537 2605 26540
rect 2639 26537 2651 26571
rect 2593 26531 2651 26537
rect 3237 26571 3295 26577
rect 3237 26537 3249 26571
rect 3283 26568 3295 26571
rect 3326 26568 3332 26580
rect 3283 26540 3332 26568
rect 3283 26537 3295 26540
rect 3237 26531 3295 26537
rect 3326 26528 3332 26540
rect 3384 26528 3390 26580
rect 4798 26528 4804 26580
rect 4856 26568 4862 26580
rect 7101 26571 7159 26577
rect 7101 26568 7113 26571
rect 4856 26540 7113 26568
rect 4856 26528 4862 26540
rect 7101 26537 7113 26540
rect 7147 26537 7159 26571
rect 7101 26531 7159 26537
rect 8481 26571 8539 26577
rect 8481 26537 8493 26571
rect 8527 26568 8539 26571
rect 12434 26568 12440 26580
rect 8527 26540 12440 26568
rect 8527 26537 8539 26540
rect 8481 26531 8539 26537
rect 12434 26528 12440 26540
rect 12492 26528 12498 26580
rect 12526 26528 12532 26580
rect 12584 26568 12590 26580
rect 12584 26540 12629 26568
rect 12584 26528 12590 26540
rect 12710 26528 12716 26580
rect 12768 26568 12774 26580
rect 16209 26571 16267 26577
rect 12768 26540 13216 26568
rect 12768 26528 12774 26540
rect 13078 26500 13084 26512
rect 10796 26472 13084 26500
rect 10796 26444 10824 26472
rect 13078 26460 13084 26472
rect 13136 26460 13142 26512
rect 13188 26500 13216 26540
rect 16209 26537 16221 26571
rect 16255 26568 16267 26571
rect 17402 26568 17408 26580
rect 16255 26540 17408 26568
rect 16255 26537 16267 26540
rect 16209 26531 16267 26537
rect 17402 26528 17408 26540
rect 17460 26528 17466 26580
rect 18049 26571 18107 26577
rect 18049 26537 18061 26571
rect 18095 26568 18107 26571
rect 18230 26568 18236 26580
rect 18095 26540 18236 26568
rect 18095 26537 18107 26540
rect 18049 26531 18107 26537
rect 18230 26528 18236 26540
rect 18288 26528 18294 26580
rect 18414 26528 18420 26580
rect 18472 26568 18478 26580
rect 22462 26568 22468 26580
rect 18472 26540 22468 26568
rect 18472 26528 18478 26540
rect 22462 26528 22468 26540
rect 22520 26528 22526 26580
rect 22646 26568 22652 26580
rect 22607 26540 22652 26568
rect 22646 26528 22652 26540
rect 22704 26528 22710 26580
rect 23290 26568 23296 26580
rect 23251 26540 23296 26568
rect 23290 26528 23296 26540
rect 23348 26528 23354 26580
rect 29822 26568 29828 26580
rect 29783 26540 29828 26568
rect 29822 26528 29828 26540
rect 29880 26528 29886 26580
rect 13188 26472 13952 26500
rect 4985 26435 5043 26441
rect 4985 26401 4997 26435
rect 5031 26432 5043 26435
rect 6546 26432 6552 26444
rect 5031 26404 6552 26432
rect 5031 26401 5043 26404
rect 4985 26395 5043 26401
rect 6546 26392 6552 26404
rect 6604 26392 6610 26444
rect 7837 26435 7895 26441
rect 7837 26401 7849 26435
rect 7883 26432 7895 26435
rect 7883 26404 10364 26432
rect 7883 26401 7895 26404
rect 7837 26395 7895 26401
rect 1857 26367 1915 26373
rect 1857 26333 1869 26367
rect 1903 26364 1915 26367
rect 2222 26364 2228 26376
rect 1903 26336 2228 26364
rect 1903 26333 1915 26336
rect 1857 26327 1915 26333
rect 2222 26324 2228 26336
rect 2280 26364 2286 26376
rect 2682 26364 2688 26376
rect 2280 26336 2688 26364
rect 2280 26324 2286 26336
rect 2682 26324 2688 26336
rect 2740 26324 2746 26376
rect 2866 26324 2872 26376
rect 2924 26364 2930 26376
rect 3145 26367 3203 26373
rect 3145 26364 3157 26367
rect 2924 26336 3157 26364
rect 2924 26324 2930 26336
rect 3145 26333 3157 26336
rect 3191 26333 3203 26367
rect 3145 26327 3203 26333
rect 6089 26367 6147 26373
rect 6089 26333 6101 26367
rect 6135 26364 6147 26367
rect 7282 26364 7288 26376
rect 6135 26336 7288 26364
rect 6135 26333 6147 26336
rect 6089 26327 6147 26333
rect 7282 26324 7288 26336
rect 7340 26324 7346 26376
rect 7929 26367 7987 26373
rect 7929 26333 7941 26367
rect 7975 26333 7987 26367
rect 8386 26364 8392 26376
rect 8299 26336 8392 26364
rect 7929 26327 7987 26333
rect 2590 26256 2596 26308
rect 2648 26296 2654 26308
rect 4433 26299 4491 26305
rect 2648 26268 2774 26296
rect 2648 26256 2654 26268
rect 2746 26228 2774 26268
rect 4433 26265 4445 26299
rect 4479 26296 4491 26299
rect 5534 26296 5540 26308
rect 4479 26268 5540 26296
rect 4479 26265 4491 26268
rect 4433 26259 4491 26265
rect 5534 26256 5540 26268
rect 5592 26256 5598 26308
rect 7944 26296 7972 26327
rect 8386 26324 8392 26336
rect 8444 26364 8450 26376
rect 9030 26364 9036 26376
rect 8444 26336 9036 26364
rect 8444 26324 8450 26336
rect 9030 26324 9036 26336
rect 9088 26324 9094 26376
rect 8938 26296 8944 26308
rect 7944 26268 8944 26296
rect 8938 26256 8944 26268
rect 8996 26256 9002 26308
rect 9214 26296 9220 26308
rect 9175 26268 9220 26296
rect 9214 26256 9220 26268
rect 9272 26256 9278 26308
rect 9306 26256 9312 26308
rect 9364 26296 9370 26308
rect 9364 26268 9409 26296
rect 9364 26256 9370 26268
rect 9858 26256 9864 26308
rect 9916 26296 9922 26308
rect 10226 26296 10232 26308
rect 9916 26268 10232 26296
rect 9916 26256 9922 26268
rect 10226 26256 10232 26268
rect 10284 26256 10290 26308
rect 10336 26296 10364 26404
rect 10502 26392 10508 26444
rect 10560 26432 10566 26444
rect 10689 26435 10747 26441
rect 10689 26432 10701 26435
rect 10560 26404 10701 26432
rect 10560 26392 10566 26404
rect 10689 26401 10701 26404
rect 10735 26401 10747 26435
rect 10689 26395 10747 26401
rect 10778 26392 10784 26444
rect 10836 26392 10842 26444
rect 11330 26432 11336 26444
rect 11291 26404 11336 26432
rect 11330 26392 11336 26404
rect 11388 26392 11394 26444
rect 11790 26392 11796 26444
rect 11848 26432 11854 26444
rect 11848 26404 13860 26432
rect 11848 26392 11854 26404
rect 11977 26367 12035 26373
rect 11977 26333 11989 26367
rect 12023 26364 12035 26367
rect 12710 26364 12716 26376
rect 12023 26336 12716 26364
rect 12023 26333 12035 26336
rect 11977 26327 12035 26333
rect 12710 26324 12716 26336
rect 12768 26324 12774 26376
rect 11425 26299 11483 26305
rect 11425 26296 11437 26299
rect 10336 26268 11437 26296
rect 11425 26265 11437 26268
rect 11471 26265 11483 26299
rect 13078 26296 13084 26308
rect 13039 26268 13084 26296
rect 11425 26259 11483 26265
rect 13078 26256 13084 26268
rect 13136 26256 13142 26308
rect 13173 26299 13231 26305
rect 13173 26265 13185 26299
rect 13219 26296 13231 26299
rect 13354 26296 13360 26308
rect 13219 26268 13360 26296
rect 13219 26265 13231 26268
rect 13173 26259 13231 26265
rect 13354 26256 13360 26268
rect 13412 26256 13418 26308
rect 13722 26296 13728 26308
rect 13683 26268 13728 26296
rect 13722 26256 13728 26268
rect 13780 26256 13786 26308
rect 13832 26296 13860 26404
rect 13924 26364 13952 26472
rect 13998 26460 14004 26512
rect 14056 26500 14062 26512
rect 15378 26500 15384 26512
rect 14056 26472 15384 26500
rect 14056 26460 14062 26472
rect 15378 26460 15384 26472
rect 15436 26460 15442 26512
rect 15565 26503 15623 26509
rect 15565 26469 15577 26503
rect 15611 26500 15623 26503
rect 15746 26500 15752 26512
rect 15611 26472 15752 26500
rect 15611 26469 15623 26472
rect 15565 26463 15623 26469
rect 15746 26460 15752 26472
rect 15804 26500 15810 26512
rect 16853 26503 16911 26509
rect 16853 26500 16865 26503
rect 15804 26472 16865 26500
rect 15804 26460 15810 26472
rect 16853 26469 16865 26472
rect 16899 26469 16911 26503
rect 18785 26503 18843 26509
rect 16853 26463 16911 26469
rect 16960 26472 17724 26500
rect 14461 26435 14519 26441
rect 14461 26401 14473 26435
rect 14507 26432 14519 26435
rect 16482 26432 16488 26444
rect 14507 26404 16488 26432
rect 14507 26401 14519 26404
rect 14461 26395 14519 26401
rect 16482 26392 16488 26404
rect 16540 26392 16546 26444
rect 16960 26432 16988 26472
rect 16592 26404 16988 26432
rect 17405 26435 17463 26441
rect 14734 26364 14740 26376
rect 13924 26336 14740 26364
rect 14734 26324 14740 26336
rect 14792 26324 14798 26376
rect 16117 26367 16175 26373
rect 16117 26333 16129 26367
rect 16163 26333 16175 26367
rect 16117 26327 16175 26333
rect 13832 26268 14780 26296
rect 4982 26228 4988 26240
rect 2746 26200 4988 26228
rect 4982 26188 4988 26200
rect 5040 26188 5046 26240
rect 5350 26188 5356 26240
rect 5408 26228 5414 26240
rect 6641 26231 6699 26237
rect 6641 26228 6653 26231
rect 5408 26200 6653 26228
rect 5408 26188 5414 26200
rect 6641 26197 6653 26200
rect 6687 26228 6699 26231
rect 8386 26228 8392 26240
rect 6687 26200 8392 26228
rect 6687 26197 6699 26200
rect 6641 26191 6699 26197
rect 8386 26188 8392 26200
rect 8444 26188 8450 26240
rect 9122 26188 9128 26240
rect 9180 26228 9186 26240
rect 11330 26228 11336 26240
rect 9180 26200 11336 26228
rect 9180 26188 9186 26200
rect 11330 26188 11336 26200
rect 11388 26188 11394 26240
rect 14752 26228 14780 26268
rect 14826 26256 14832 26308
rect 14884 26296 14890 26308
rect 15013 26299 15071 26305
rect 15013 26296 15025 26299
rect 14884 26268 15025 26296
rect 14884 26256 14890 26268
rect 15013 26265 15025 26268
rect 15059 26265 15071 26299
rect 15013 26259 15071 26265
rect 15105 26299 15163 26305
rect 15105 26265 15117 26299
rect 15151 26265 15163 26299
rect 15105 26259 15163 26265
rect 15120 26228 15148 26259
rect 15378 26256 15384 26308
rect 15436 26296 15442 26308
rect 16132 26296 16160 26327
rect 16298 26324 16304 26376
rect 16356 26364 16362 26376
rect 16592 26364 16620 26404
rect 17405 26401 17417 26435
rect 17451 26432 17463 26435
rect 17586 26432 17592 26444
rect 17451 26404 17592 26432
rect 17451 26401 17463 26404
rect 17405 26395 17463 26401
rect 17586 26392 17592 26404
rect 17644 26392 17650 26444
rect 17696 26432 17724 26472
rect 18785 26469 18797 26503
rect 18831 26500 18843 26503
rect 20073 26503 20131 26509
rect 18831 26472 19472 26500
rect 18831 26469 18843 26472
rect 18785 26463 18843 26469
rect 19444 26432 19472 26472
rect 20073 26469 20085 26503
rect 20119 26500 20131 26503
rect 20622 26500 20628 26512
rect 20119 26472 20628 26500
rect 20119 26469 20131 26472
rect 20073 26463 20131 26469
rect 20622 26460 20628 26472
rect 20680 26460 20686 26512
rect 19510 26435 19568 26441
rect 19510 26432 19522 26435
rect 17696 26404 19334 26432
rect 19444 26404 19522 26432
rect 19306 26376 19334 26404
rect 19510 26401 19522 26404
rect 19556 26401 19568 26435
rect 19510 26395 19568 26401
rect 20530 26392 20536 26444
rect 20588 26432 20594 26444
rect 21545 26435 21603 26441
rect 21545 26432 21557 26435
rect 20588 26404 21557 26432
rect 20588 26392 20594 26404
rect 21545 26401 21557 26404
rect 21591 26432 21603 26435
rect 26234 26432 26240 26444
rect 21591 26404 26240 26432
rect 21591 26401 21603 26404
rect 21545 26395 21603 26401
rect 26234 26392 26240 26404
rect 26292 26392 26298 26444
rect 18782 26364 18788 26376
rect 16356 26336 16620 26364
rect 18743 26336 18788 26364
rect 16356 26324 16362 26336
rect 18782 26324 18788 26336
rect 18840 26324 18846 26376
rect 19306 26336 19340 26376
rect 19334 26324 19340 26336
rect 19392 26324 19398 26376
rect 20898 26364 20904 26376
rect 20859 26336 20904 26364
rect 20898 26324 20904 26336
rect 20956 26324 20962 26376
rect 22738 26364 22744 26376
rect 22699 26336 22744 26364
rect 22738 26324 22744 26336
rect 22796 26324 22802 26376
rect 23198 26364 23204 26376
rect 23111 26336 23204 26364
rect 23198 26324 23204 26336
rect 23256 26364 23262 26376
rect 24581 26367 24639 26373
rect 24581 26364 24593 26367
rect 23256 26336 24593 26364
rect 23256 26324 23262 26336
rect 24581 26333 24593 26336
rect 24627 26333 24639 26367
rect 24581 26327 24639 26333
rect 29917 26367 29975 26373
rect 29917 26333 29929 26367
rect 29963 26364 29975 26367
rect 37918 26364 37924 26376
rect 29963 26336 37924 26364
rect 29963 26333 29975 26336
rect 29917 26327 29975 26333
rect 37918 26324 37924 26336
rect 37976 26324 37982 26376
rect 17310 26296 17316 26308
rect 15436 26268 17172 26296
rect 17271 26268 17316 26296
rect 15436 26256 15442 26268
rect 14752 26200 15148 26228
rect 17144 26228 17172 26268
rect 17310 26256 17316 26268
rect 17368 26256 17374 26308
rect 19613 26299 19671 26305
rect 17420 26268 19288 26296
rect 17420 26228 17448 26268
rect 17144 26200 17448 26228
rect 18230 26188 18236 26240
rect 18288 26228 18294 26240
rect 19150 26228 19156 26240
rect 18288 26200 19156 26228
rect 18288 26188 18294 26200
rect 19150 26188 19156 26200
rect 19208 26188 19214 26240
rect 19260 26228 19288 26268
rect 19613 26265 19625 26299
rect 19659 26296 19671 26299
rect 19659 26268 19748 26296
rect 19659 26265 19671 26268
rect 19613 26259 19671 26265
rect 19518 26228 19524 26240
rect 19260 26200 19524 26228
rect 19518 26188 19524 26200
rect 19576 26188 19582 26240
rect 19720 26228 19748 26268
rect 21358 26256 21364 26308
rect 21416 26296 21422 26308
rect 21453 26299 21511 26305
rect 21453 26296 21465 26299
rect 21416 26268 21465 26296
rect 21416 26256 21422 26268
rect 21453 26265 21465 26268
rect 21499 26265 21511 26299
rect 22756 26296 22784 26324
rect 23845 26299 23903 26305
rect 23845 26296 23857 26299
rect 22756 26268 23857 26296
rect 21453 26259 21511 26265
rect 23845 26265 23857 26268
rect 23891 26265 23903 26299
rect 23845 26259 23903 26265
rect 19794 26228 19800 26240
rect 19720 26200 19800 26228
rect 19794 26188 19800 26200
rect 19852 26188 19858 26240
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 1302 25984 1308 26036
rect 1360 26024 1366 26036
rect 1949 26027 2007 26033
rect 1949 26024 1961 26027
rect 1360 25996 1961 26024
rect 1360 25984 1366 25996
rect 1949 25993 1961 25996
rect 1995 25993 2007 26027
rect 1949 25987 2007 25993
rect 2498 25984 2504 26036
rect 2556 26024 2562 26036
rect 2593 26027 2651 26033
rect 2593 26024 2605 26027
rect 2556 25996 2605 26024
rect 2556 25984 2562 25996
rect 2593 25993 2605 25996
rect 2639 25993 2651 26027
rect 2593 25987 2651 25993
rect 6641 26027 6699 26033
rect 6641 25993 6653 26027
rect 6687 26024 6699 26027
rect 7742 26024 7748 26036
rect 6687 25996 7748 26024
rect 6687 25993 6699 25996
rect 6641 25987 6699 25993
rect 7742 25984 7748 25996
rect 7800 25984 7806 26036
rect 7837 26027 7895 26033
rect 7837 25993 7849 26027
rect 7883 26024 7895 26027
rect 11790 26024 11796 26036
rect 7883 25996 10640 26024
rect 11751 25996 11796 26024
rect 7883 25993 7895 25996
rect 7837 25987 7895 25993
rect 3878 25916 3884 25968
rect 3936 25956 3942 25968
rect 3936 25928 7880 25956
rect 3936 25916 3942 25928
rect 1857 25891 1915 25897
rect 1857 25857 1869 25891
rect 1903 25888 1915 25891
rect 2501 25891 2559 25897
rect 2501 25888 2513 25891
rect 1903 25860 2513 25888
rect 1903 25857 1915 25860
rect 1857 25851 1915 25857
rect 2501 25857 2513 25860
rect 2547 25888 2559 25891
rect 2866 25888 2872 25900
rect 2547 25860 2872 25888
rect 2547 25857 2559 25860
rect 2501 25851 2559 25857
rect 2866 25848 2872 25860
rect 2924 25848 2930 25900
rect 5810 25888 5816 25900
rect 5771 25860 5816 25888
rect 5810 25848 5816 25860
rect 5868 25848 5874 25900
rect 7098 25888 7104 25900
rect 7059 25860 7104 25888
rect 7098 25848 7104 25860
rect 7156 25848 7162 25900
rect 7650 25848 7656 25900
rect 7708 25888 7714 25900
rect 7745 25891 7803 25897
rect 7745 25888 7757 25891
rect 7708 25860 7757 25888
rect 7708 25848 7714 25860
rect 7745 25857 7757 25860
rect 7791 25857 7803 25891
rect 7852 25888 7880 25928
rect 7926 25916 7932 25968
rect 7984 25956 7990 25968
rect 9217 25959 9275 25965
rect 9217 25956 9229 25959
rect 7984 25928 9229 25956
rect 7984 25916 7990 25928
rect 9217 25925 9229 25928
rect 9263 25925 9275 25959
rect 9217 25919 9275 25925
rect 9398 25916 9404 25968
rect 9456 25956 9462 25968
rect 10502 25956 10508 25968
rect 9456 25928 10508 25956
rect 9456 25916 9462 25928
rect 10502 25916 10508 25928
rect 10560 25916 10566 25968
rect 10612 25965 10640 25996
rect 11790 25984 11796 25996
rect 11848 25984 11854 26036
rect 11882 25984 11888 26036
rect 11940 26024 11946 26036
rect 17221 26027 17279 26033
rect 11940 25996 15884 26024
rect 11940 25984 11946 25996
rect 10597 25959 10655 25965
rect 10597 25925 10609 25959
rect 10643 25925 10655 25959
rect 11146 25956 11152 25968
rect 11107 25928 11152 25956
rect 10597 25919 10655 25925
rect 11146 25916 11152 25928
rect 11204 25916 11210 25968
rect 12526 25956 12532 25968
rect 11256 25928 11836 25956
rect 12487 25928 12532 25956
rect 8389 25891 8447 25897
rect 8389 25888 8401 25891
rect 7852 25860 8401 25888
rect 7745 25851 7803 25857
rect 8389 25857 8401 25860
rect 8435 25857 8447 25891
rect 8389 25851 8447 25857
rect 3697 25823 3755 25829
rect 3697 25789 3709 25823
rect 3743 25820 3755 25823
rect 6178 25820 6184 25832
rect 3743 25792 6184 25820
rect 3743 25789 3755 25792
rect 3697 25783 3755 25789
rect 6178 25780 6184 25792
rect 6236 25780 6242 25832
rect 7760 25820 7788 25851
rect 8570 25820 8576 25832
rect 7760 25792 8576 25820
rect 8570 25780 8576 25792
rect 8628 25780 8634 25832
rect 9122 25820 9128 25832
rect 9083 25792 9128 25820
rect 9122 25780 9128 25792
rect 9180 25780 9186 25832
rect 9858 25780 9864 25832
rect 9916 25820 9922 25832
rect 10505 25823 10563 25829
rect 10505 25820 10517 25823
rect 9916 25792 10517 25820
rect 9916 25780 9922 25792
rect 10505 25789 10517 25792
rect 10551 25820 10563 25823
rect 11256 25820 11284 25928
rect 11701 25891 11759 25897
rect 11701 25857 11713 25891
rect 11747 25857 11759 25891
rect 11701 25851 11759 25857
rect 10551 25792 11284 25820
rect 10551 25789 10563 25792
rect 10505 25783 10563 25789
rect 4801 25755 4859 25761
rect 4801 25721 4813 25755
rect 4847 25752 4859 25755
rect 5810 25752 5816 25764
rect 4847 25724 5816 25752
rect 4847 25721 4859 25724
rect 4801 25715 4859 25721
rect 5810 25712 5816 25724
rect 5868 25712 5874 25764
rect 5905 25755 5963 25761
rect 5905 25721 5917 25755
rect 5951 25752 5963 25755
rect 8202 25752 8208 25764
rect 5951 25724 8208 25752
rect 5951 25721 5963 25724
rect 5905 25715 5963 25721
rect 8202 25712 8208 25724
rect 8260 25712 8266 25764
rect 9214 25712 9220 25764
rect 9272 25752 9278 25764
rect 9677 25755 9735 25761
rect 9677 25752 9689 25755
rect 9272 25724 9689 25752
rect 9272 25712 9278 25724
rect 9677 25721 9689 25724
rect 9723 25752 9735 25755
rect 11146 25752 11152 25764
rect 9723 25724 11152 25752
rect 9723 25721 9735 25724
rect 9677 25715 9735 25721
rect 11146 25712 11152 25724
rect 11204 25712 11210 25764
rect 11716 25752 11744 25851
rect 11808 25820 11836 25928
rect 12526 25916 12532 25928
rect 12584 25916 12590 25968
rect 13446 25916 13452 25968
rect 13504 25956 13510 25968
rect 13725 25959 13783 25965
rect 13725 25956 13737 25959
rect 13504 25928 13737 25956
rect 13504 25916 13510 25928
rect 13725 25925 13737 25928
rect 13771 25925 13783 25959
rect 13725 25919 13783 25925
rect 14277 25959 14335 25965
rect 14277 25925 14289 25959
rect 14323 25956 14335 25959
rect 14366 25956 14372 25968
rect 14323 25928 14372 25956
rect 14323 25925 14335 25928
rect 14277 25919 14335 25925
rect 14366 25916 14372 25928
rect 14424 25916 14430 25968
rect 14458 25916 14464 25968
rect 14516 25956 14522 25968
rect 14737 25959 14795 25965
rect 14737 25956 14749 25959
rect 14516 25928 14749 25956
rect 14516 25916 14522 25928
rect 14737 25925 14749 25928
rect 14783 25925 14795 25959
rect 15286 25956 15292 25968
rect 15247 25928 15292 25956
rect 14737 25919 14795 25925
rect 15286 25916 15292 25928
rect 15344 25916 15350 25968
rect 15381 25959 15439 25965
rect 15381 25925 15393 25959
rect 15427 25956 15439 25959
rect 15746 25956 15752 25968
rect 15427 25928 15752 25956
rect 15427 25925 15439 25928
rect 15381 25919 15439 25925
rect 15746 25916 15752 25928
rect 15804 25916 15810 25968
rect 15856 25956 15884 25996
rect 17221 25993 17233 26027
rect 17267 26024 17279 26027
rect 17310 26024 17316 26036
rect 17267 25996 17316 26024
rect 17267 25993 17279 25996
rect 17221 25987 17279 25993
rect 17310 25984 17316 25996
rect 17368 25984 17374 26036
rect 17494 25984 17500 26036
rect 17552 26024 17558 26036
rect 17865 26027 17923 26033
rect 17865 26024 17877 26027
rect 17552 25996 17877 26024
rect 17552 25984 17558 25996
rect 17865 25993 17877 25996
rect 17911 25993 17923 26027
rect 17865 25987 17923 25993
rect 18509 26027 18567 26033
rect 18509 25993 18521 26027
rect 18555 26024 18567 26027
rect 18690 26024 18696 26036
rect 18555 25996 18696 26024
rect 18555 25993 18567 25996
rect 18509 25987 18567 25993
rect 18690 25984 18696 25996
rect 18748 25984 18754 26036
rect 20714 26024 20720 26036
rect 20675 25996 20720 26024
rect 20714 25984 20720 25996
rect 20772 25984 20778 26036
rect 20990 25984 20996 26036
rect 21048 26024 21054 26036
rect 21361 26027 21419 26033
rect 21361 26024 21373 26027
rect 21048 25996 21373 26024
rect 21048 25984 21054 25996
rect 21361 25993 21373 25996
rect 21407 25993 21419 26027
rect 22738 26024 22744 26036
rect 21361 25987 21419 25993
rect 22066 25996 22744 26024
rect 19245 25959 19303 25965
rect 19245 25956 19257 25959
rect 15856 25928 19257 25956
rect 19245 25925 19257 25928
rect 19291 25925 19303 25959
rect 19245 25919 19303 25925
rect 19334 25916 19340 25968
rect 19392 25956 19398 25968
rect 20070 25956 20076 25968
rect 19392 25928 20076 25956
rect 19392 25916 19398 25928
rect 20070 25916 20076 25928
rect 20128 25956 20134 25968
rect 22066 25956 22094 25996
rect 22738 25984 22744 25996
rect 22796 26024 22802 26036
rect 23198 26024 23204 26036
rect 22796 25996 23204 26024
rect 22796 25984 22802 25996
rect 23198 25984 23204 25996
rect 23256 25984 23262 26036
rect 20128 25928 22094 25956
rect 22557 25959 22615 25965
rect 20128 25916 20134 25928
rect 14642 25848 14648 25900
rect 14700 25848 14706 25900
rect 16206 25848 16212 25900
rect 16264 25888 16270 25900
rect 16301 25891 16359 25897
rect 16301 25888 16313 25891
rect 16264 25860 16313 25888
rect 16264 25848 16270 25860
rect 16301 25857 16313 25860
rect 16347 25857 16359 25891
rect 16301 25851 16359 25857
rect 16850 25848 16856 25900
rect 16908 25888 16914 25900
rect 17126 25888 17132 25900
rect 16908 25860 17132 25888
rect 16908 25848 16914 25860
rect 17126 25848 17132 25860
rect 17184 25848 17190 25900
rect 17954 25888 17960 25900
rect 17915 25860 17960 25888
rect 17954 25848 17960 25860
rect 18012 25848 18018 25900
rect 18138 25848 18144 25900
rect 18196 25888 18202 25900
rect 18417 25891 18475 25897
rect 18417 25888 18429 25891
rect 18196 25860 18429 25888
rect 18196 25848 18202 25860
rect 18417 25857 18429 25860
rect 18463 25857 18475 25891
rect 20622 25888 20628 25900
rect 20583 25860 20628 25888
rect 18417 25851 18475 25857
rect 20622 25848 20628 25860
rect 20680 25848 20686 25900
rect 21468 25897 21496 25928
rect 22557 25925 22569 25959
rect 22603 25956 22615 25959
rect 23293 25959 23351 25965
rect 23293 25956 23305 25959
rect 22603 25928 23305 25956
rect 22603 25925 22615 25928
rect 22557 25919 22615 25925
rect 23293 25925 23305 25928
rect 23339 25925 23351 25959
rect 23293 25919 23351 25925
rect 21453 25891 21511 25897
rect 21453 25857 21465 25891
rect 21499 25857 21511 25891
rect 21453 25851 21511 25857
rect 22830 25848 22836 25900
rect 22888 25888 22894 25900
rect 23385 25891 23443 25897
rect 23385 25888 23397 25891
rect 22888 25860 23397 25888
rect 22888 25848 22894 25860
rect 23385 25857 23397 25860
rect 23431 25888 23443 25891
rect 23845 25891 23903 25897
rect 23845 25888 23857 25891
rect 23431 25860 23857 25888
rect 23431 25857 23443 25860
rect 23385 25851 23443 25857
rect 23845 25857 23857 25860
rect 23891 25857 23903 25891
rect 23845 25851 23903 25857
rect 12437 25823 12495 25829
rect 12437 25820 12449 25823
rect 11808 25792 12449 25820
rect 12437 25789 12449 25792
rect 12483 25789 12495 25823
rect 13633 25823 13691 25829
rect 13633 25820 13645 25823
rect 12437 25783 12495 25789
rect 12544 25792 13645 25820
rect 11716 25724 12112 25752
rect 4249 25687 4307 25693
rect 4249 25653 4261 25687
rect 4295 25684 4307 25687
rect 4614 25684 4620 25696
rect 4295 25656 4620 25684
rect 4295 25653 4307 25656
rect 4249 25647 4307 25653
rect 4614 25644 4620 25656
rect 4672 25644 4678 25696
rect 5353 25687 5411 25693
rect 5353 25653 5365 25687
rect 5399 25684 5411 25687
rect 5534 25684 5540 25696
rect 5399 25656 5540 25684
rect 5399 25653 5411 25656
rect 5353 25647 5411 25653
rect 5534 25644 5540 25656
rect 5592 25644 5598 25696
rect 7190 25684 7196 25696
rect 7151 25656 7196 25684
rect 7190 25644 7196 25656
rect 7248 25644 7254 25696
rect 8481 25687 8539 25693
rect 8481 25653 8493 25687
rect 8527 25684 8539 25687
rect 9766 25684 9772 25696
rect 8527 25656 9772 25684
rect 8527 25653 8539 25656
rect 8481 25647 8539 25653
rect 9766 25644 9772 25656
rect 9824 25644 9830 25696
rect 12084 25684 12112 25724
rect 12158 25712 12164 25764
rect 12216 25752 12222 25764
rect 12544 25752 12572 25792
rect 13633 25789 13645 25792
rect 13679 25820 13691 25823
rect 14660 25820 14688 25848
rect 19153 25823 19211 25829
rect 13679 25792 14688 25820
rect 14844 25808 15332 25820
rect 15672 25808 19104 25820
rect 14844 25792 19104 25808
rect 13679 25789 13691 25792
rect 13633 25783 13691 25789
rect 12216 25724 12572 25752
rect 12989 25755 13047 25761
rect 12216 25712 12222 25724
rect 12989 25721 13001 25755
rect 13035 25721 13047 25755
rect 12989 25715 13047 25721
rect 12710 25684 12716 25696
rect 12084 25656 12716 25684
rect 12710 25644 12716 25656
rect 12768 25644 12774 25696
rect 13004 25684 13032 25715
rect 13446 25712 13452 25764
rect 13504 25752 13510 25764
rect 14458 25752 14464 25764
rect 13504 25724 14464 25752
rect 13504 25712 13510 25724
rect 14458 25712 14464 25724
rect 14516 25712 14522 25764
rect 14734 25712 14740 25764
rect 14792 25752 14798 25764
rect 14844 25752 14872 25792
rect 15304 25780 15700 25792
rect 16022 25752 16028 25764
rect 14792 25724 14872 25752
rect 14936 25724 16028 25752
rect 14792 25712 14798 25724
rect 14642 25684 14648 25696
rect 13004 25656 14648 25684
rect 14642 25644 14648 25656
rect 14700 25684 14706 25696
rect 14936 25684 14964 25724
rect 16022 25712 16028 25724
rect 16080 25712 16086 25764
rect 19076 25752 19104 25792
rect 19153 25789 19165 25823
rect 19199 25820 19211 25823
rect 20070 25820 20076 25832
rect 19199 25792 20076 25820
rect 19199 25789 19211 25792
rect 19153 25783 19211 25789
rect 20070 25780 20076 25792
rect 20128 25780 20134 25832
rect 20162 25780 20168 25832
rect 20220 25820 20226 25832
rect 22646 25820 22652 25832
rect 20220 25792 20265 25820
rect 22607 25792 22652 25820
rect 20220 25780 20226 25792
rect 22646 25780 22652 25792
rect 22704 25780 22710 25832
rect 19334 25752 19340 25764
rect 19076 25724 19340 25752
rect 19334 25712 19340 25724
rect 19392 25712 19398 25764
rect 22097 25755 22155 25761
rect 22097 25721 22109 25755
rect 22143 25752 22155 25755
rect 23566 25752 23572 25764
rect 22143 25724 23572 25752
rect 22143 25721 22155 25724
rect 22097 25715 22155 25721
rect 23566 25712 23572 25724
rect 23624 25712 23630 25764
rect 14700 25656 14964 25684
rect 14700 25644 14706 25656
rect 15378 25644 15384 25696
rect 15436 25684 15442 25696
rect 16209 25687 16267 25693
rect 16209 25684 16221 25687
rect 15436 25656 16221 25684
rect 15436 25644 15442 25656
rect 16209 25653 16221 25656
rect 16255 25653 16267 25687
rect 16209 25647 16267 25653
rect 17402 25644 17408 25696
rect 17460 25684 17466 25696
rect 23106 25684 23112 25696
rect 17460 25656 23112 25684
rect 17460 25644 17466 25656
rect 23106 25644 23112 25656
rect 23164 25644 23170 25696
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 2222 25480 2228 25492
rect 2183 25452 2228 25480
rect 2222 25440 2228 25452
rect 2280 25480 2286 25492
rect 2777 25483 2835 25489
rect 2777 25480 2789 25483
rect 2280 25452 2789 25480
rect 2280 25440 2286 25452
rect 2777 25449 2789 25452
rect 2823 25449 2835 25483
rect 4982 25480 4988 25492
rect 4943 25452 4988 25480
rect 2777 25443 2835 25449
rect 4982 25440 4988 25452
rect 5040 25440 5046 25492
rect 5074 25440 5080 25492
rect 5132 25480 5138 25492
rect 5537 25483 5595 25489
rect 5537 25480 5549 25483
rect 5132 25452 5549 25480
rect 5132 25440 5138 25452
rect 5537 25449 5549 25452
rect 5583 25449 5595 25483
rect 5537 25443 5595 25449
rect 7285 25483 7343 25489
rect 7285 25449 7297 25483
rect 7331 25480 7343 25483
rect 9122 25480 9128 25492
rect 7331 25452 9128 25480
rect 7331 25449 7343 25452
rect 7285 25443 7343 25449
rect 9122 25440 9128 25452
rect 9180 25440 9186 25492
rect 9309 25483 9367 25489
rect 9309 25449 9321 25483
rect 9355 25480 9367 25483
rect 12526 25480 12532 25492
rect 9355 25452 12532 25480
rect 9355 25449 9367 25452
rect 9309 25443 9367 25449
rect 12526 25440 12532 25452
rect 12584 25440 12590 25492
rect 12618 25440 12624 25492
rect 12676 25480 12682 25492
rect 14734 25480 14740 25492
rect 12676 25452 14740 25480
rect 12676 25440 12682 25452
rect 14734 25440 14740 25452
rect 14792 25440 14798 25492
rect 15010 25440 15016 25492
rect 15068 25480 15074 25492
rect 15068 25452 18460 25480
rect 15068 25440 15074 25452
rect 7190 25372 7196 25424
rect 7248 25412 7254 25424
rect 12158 25412 12164 25424
rect 7248 25384 12164 25412
rect 7248 25372 7254 25384
rect 6733 25347 6791 25353
rect 6733 25313 6745 25347
rect 6779 25344 6791 25347
rect 7929 25347 7987 25353
rect 6779 25316 7880 25344
rect 6779 25313 6791 25316
rect 6733 25307 6791 25313
rect 5626 25236 5632 25288
rect 5684 25276 5690 25288
rect 7193 25279 7251 25285
rect 7193 25276 7205 25279
rect 5684 25248 7205 25276
rect 5684 25236 5690 25248
rect 7193 25245 7205 25248
rect 7239 25245 7251 25279
rect 7852 25276 7880 25316
rect 7929 25313 7941 25347
rect 7975 25344 7987 25347
rect 8386 25344 8392 25356
rect 7975 25316 8392 25344
rect 7975 25313 7987 25316
rect 7929 25307 7987 25313
rect 8386 25304 8392 25316
rect 8444 25344 8450 25356
rect 9398 25344 9404 25356
rect 8444 25316 9404 25344
rect 8444 25304 8450 25316
rect 9398 25304 9404 25316
rect 9456 25304 9462 25356
rect 10134 25344 10140 25356
rect 9692 25316 10140 25344
rect 9217 25279 9275 25285
rect 9217 25276 9229 25279
rect 7852 25248 9229 25276
rect 7193 25239 7251 25245
rect 9217 25245 9229 25248
rect 9263 25276 9275 25279
rect 9692 25276 9720 25316
rect 10134 25304 10140 25316
rect 10192 25304 10198 25356
rect 10229 25347 10287 25353
rect 10229 25313 10241 25347
rect 10275 25344 10287 25347
rect 10410 25344 10416 25356
rect 10275 25316 10416 25344
rect 10275 25313 10287 25316
rect 10229 25307 10287 25313
rect 10410 25304 10416 25316
rect 10468 25304 10474 25356
rect 11532 25353 11560 25384
rect 12158 25372 12164 25384
rect 12216 25372 12222 25424
rect 18432 25412 18460 25452
rect 18874 25440 18880 25492
rect 18932 25480 18938 25492
rect 21453 25483 21511 25489
rect 21453 25480 21465 25483
rect 18932 25452 21465 25480
rect 18932 25440 18938 25452
rect 21453 25449 21465 25452
rect 21499 25449 21511 25483
rect 21453 25443 21511 25449
rect 22646 25440 22652 25492
rect 22704 25480 22710 25492
rect 29825 25483 29883 25489
rect 29825 25480 29837 25483
rect 22704 25452 29837 25480
rect 22704 25440 22710 25452
rect 29825 25449 29837 25452
rect 29871 25449 29883 25483
rect 29825 25443 29883 25449
rect 20622 25412 20628 25424
rect 18432 25384 20628 25412
rect 20622 25372 20628 25384
rect 20680 25372 20686 25424
rect 11517 25347 11575 25353
rect 11517 25313 11529 25347
rect 11563 25313 11575 25347
rect 11517 25307 11575 25313
rect 11606 25304 11612 25356
rect 11664 25344 11670 25356
rect 13081 25347 13139 25353
rect 13081 25344 13093 25347
rect 11664 25316 13093 25344
rect 11664 25304 11670 25316
rect 13081 25313 13093 25316
rect 13127 25344 13139 25347
rect 15289 25347 15347 25353
rect 15289 25344 15301 25347
rect 13127 25316 15301 25344
rect 13127 25313 13139 25316
rect 13081 25307 13139 25313
rect 15289 25313 15301 25316
rect 15335 25313 15347 25347
rect 15289 25307 15347 25313
rect 15933 25347 15991 25353
rect 15933 25313 15945 25347
rect 15979 25344 15991 25347
rect 16298 25344 16304 25356
rect 15979 25316 16304 25344
rect 15979 25313 15991 25316
rect 15933 25307 15991 25313
rect 16298 25304 16304 25316
rect 16356 25304 16362 25356
rect 16482 25344 16488 25356
rect 16443 25316 16488 25344
rect 16482 25304 16488 25316
rect 16540 25304 16546 25356
rect 16758 25344 16764 25356
rect 16719 25316 16764 25344
rect 16758 25304 16764 25316
rect 16816 25304 16822 25356
rect 18414 25304 18420 25356
rect 18472 25344 18478 25356
rect 18601 25347 18659 25353
rect 18601 25344 18613 25347
rect 18472 25316 18613 25344
rect 18472 25304 18478 25316
rect 18601 25313 18613 25316
rect 18647 25313 18659 25347
rect 18601 25307 18659 25313
rect 19518 25304 19524 25356
rect 19576 25344 19582 25356
rect 22664 25344 22692 25440
rect 19576 25316 22692 25344
rect 19576 25304 19582 25316
rect 9263 25248 9720 25276
rect 9263 25245 9275 25248
rect 9217 25239 9275 25245
rect 14274 25236 14280 25288
rect 14332 25276 14338 25288
rect 14369 25279 14427 25285
rect 14369 25276 14381 25279
rect 14332 25248 14381 25276
rect 14332 25236 14338 25248
rect 14369 25245 14381 25248
rect 14415 25245 14427 25279
rect 14369 25239 14427 25245
rect 19150 25236 19156 25288
rect 19208 25276 19214 25288
rect 19334 25276 19340 25288
rect 19208 25248 19340 25276
rect 19208 25236 19214 25248
rect 19334 25236 19340 25248
rect 19392 25276 19398 25288
rect 19429 25279 19487 25285
rect 19429 25276 19441 25279
rect 19392 25248 19441 25276
rect 19392 25236 19398 25248
rect 19429 25245 19441 25248
rect 19475 25245 19487 25279
rect 19429 25239 19487 25245
rect 21545 25279 21603 25285
rect 21545 25245 21557 25279
rect 21591 25276 21603 25279
rect 22094 25276 22100 25288
rect 21591 25248 22100 25276
rect 21591 25245 21603 25248
rect 21545 25239 21603 25245
rect 22094 25236 22100 25248
rect 22152 25276 22158 25288
rect 29917 25279 29975 25285
rect 22152 25248 22245 25276
rect 22152 25236 22158 25248
rect 29917 25245 29929 25279
rect 29963 25276 29975 25279
rect 37826 25276 37832 25288
rect 29963 25248 37832 25276
rect 29963 25245 29975 25248
rect 29917 25239 29975 25245
rect 37826 25236 37832 25248
rect 37884 25236 37890 25288
rect 1765 25211 1823 25217
rect 1765 25177 1777 25211
rect 1811 25208 1823 25211
rect 2866 25208 2872 25220
rect 1811 25180 2872 25208
rect 1811 25177 1823 25180
rect 1765 25171 1823 25177
rect 2866 25168 2872 25180
rect 2924 25168 2930 25220
rect 8478 25168 8484 25220
rect 8536 25208 8542 25220
rect 10413 25211 10471 25217
rect 10413 25208 10425 25211
rect 8536 25180 10425 25208
rect 8536 25168 8542 25180
rect 10413 25177 10425 25180
rect 10459 25177 10471 25211
rect 10413 25171 10471 25177
rect 10505 25211 10563 25217
rect 10505 25177 10517 25211
rect 10551 25208 10563 25211
rect 11618 25211 11676 25217
rect 10551 25180 11560 25208
rect 10551 25177 10563 25180
rect 10505 25171 10563 25177
rect 3418 25140 3424 25152
rect 3379 25112 3424 25140
rect 3418 25100 3424 25112
rect 3476 25100 3482 25152
rect 4525 25143 4583 25149
rect 4525 25109 4537 25143
rect 4571 25140 4583 25143
rect 4614 25140 4620 25152
rect 4571 25112 4620 25140
rect 4571 25109 4583 25112
rect 4525 25103 4583 25109
rect 4614 25100 4620 25112
rect 4672 25100 4678 25152
rect 6178 25140 6184 25152
rect 6091 25112 6184 25140
rect 6178 25100 6184 25112
rect 6236 25140 6242 25152
rect 6730 25140 6736 25152
rect 6236 25112 6736 25140
rect 6236 25100 6242 25112
rect 6730 25100 6736 25112
rect 6788 25100 6794 25152
rect 8573 25143 8631 25149
rect 8573 25109 8585 25143
rect 8619 25140 8631 25143
rect 10594 25140 10600 25152
rect 8619 25112 10600 25140
rect 8619 25109 8631 25112
rect 8573 25103 8631 25109
rect 10594 25100 10600 25112
rect 10652 25100 10658 25152
rect 11532 25140 11560 25180
rect 11618 25177 11630 25211
rect 11664 25208 11676 25211
rect 11790 25208 11796 25220
rect 11664 25180 11796 25208
rect 11664 25177 11676 25180
rect 11618 25171 11676 25177
rect 11790 25168 11796 25180
rect 11848 25168 11854 25220
rect 12161 25211 12219 25217
rect 12161 25177 12173 25211
rect 12207 25177 12219 25211
rect 12161 25171 12219 25177
rect 12066 25140 12072 25152
rect 11532 25112 12072 25140
rect 12066 25100 12072 25112
rect 12124 25140 12130 25152
rect 12176 25140 12204 25171
rect 12434 25168 12440 25220
rect 12492 25208 12498 25220
rect 13173 25211 13231 25217
rect 13173 25208 13185 25211
rect 12492 25180 13185 25208
rect 12492 25168 12498 25180
rect 13173 25177 13185 25180
rect 13219 25177 13231 25211
rect 13722 25208 13728 25220
rect 13683 25180 13728 25208
rect 13173 25171 13231 25177
rect 13722 25168 13728 25180
rect 13780 25168 13786 25220
rect 15010 25208 15016 25220
rect 13832 25180 15016 25208
rect 12124 25112 12204 25140
rect 12124 25100 12130 25112
rect 12250 25100 12256 25152
rect 12308 25140 12314 25152
rect 12618 25140 12624 25152
rect 12308 25112 12624 25140
rect 12308 25100 12314 25112
rect 12618 25100 12624 25112
rect 12676 25100 12682 25152
rect 12710 25100 12716 25152
rect 12768 25140 12774 25152
rect 13832 25140 13860 25180
rect 15010 25168 15016 25180
rect 15068 25168 15074 25220
rect 15378 25168 15384 25220
rect 15436 25208 15442 25220
rect 16577 25211 16635 25217
rect 15436 25180 15481 25208
rect 15436 25168 15442 25180
rect 16577 25177 16589 25211
rect 16623 25177 16635 25211
rect 16577 25171 16635 25177
rect 14458 25140 14464 25152
rect 12768 25112 13860 25140
rect 14419 25112 14464 25140
rect 12768 25100 12774 25112
rect 14458 25100 14464 25112
rect 14516 25100 14522 25152
rect 16592 25140 16620 25171
rect 16666 25168 16672 25220
rect 16724 25208 16730 25220
rect 17957 25211 18015 25217
rect 17957 25208 17969 25211
rect 16724 25180 17969 25208
rect 16724 25168 16730 25180
rect 17957 25177 17969 25180
rect 18003 25177 18015 25211
rect 18506 25208 18512 25220
rect 18467 25180 18512 25208
rect 17957 25171 18015 25177
rect 18506 25168 18512 25180
rect 18564 25168 18570 25220
rect 20254 25208 20260 25220
rect 20215 25180 20260 25208
rect 20254 25168 20260 25180
rect 20312 25168 20318 25220
rect 20349 25211 20407 25217
rect 20349 25177 20361 25211
rect 20395 25177 20407 25211
rect 20349 25171 20407 25177
rect 20901 25211 20959 25217
rect 20901 25177 20913 25211
rect 20947 25208 20959 25211
rect 22186 25208 22192 25220
rect 20947 25180 22192 25208
rect 20947 25177 20959 25180
rect 20901 25171 20959 25177
rect 19242 25140 19248 25152
rect 16592 25112 19248 25140
rect 19242 25100 19248 25112
rect 19300 25100 19306 25152
rect 19521 25143 19579 25149
rect 19521 25109 19533 25143
rect 19567 25140 19579 25143
rect 20364 25140 20392 25171
rect 22186 25168 22192 25180
rect 22244 25208 22250 25220
rect 23017 25211 23075 25217
rect 23017 25208 23029 25211
rect 22244 25180 23029 25208
rect 22244 25168 22250 25180
rect 23017 25177 23029 25180
rect 23063 25177 23075 25211
rect 23017 25171 23075 25177
rect 23106 25168 23112 25220
rect 23164 25208 23170 25220
rect 24026 25208 24032 25220
rect 23164 25180 23209 25208
rect 23939 25180 24032 25208
rect 23164 25168 23170 25180
rect 24026 25168 24032 25180
rect 24084 25208 24090 25220
rect 32950 25208 32956 25220
rect 24084 25180 32956 25208
rect 24084 25168 24090 25180
rect 32950 25168 32956 25180
rect 33008 25168 33014 25220
rect 38286 25140 38292 25152
rect 19567 25112 20392 25140
rect 38247 25112 38292 25140
rect 19567 25109 19579 25112
rect 19521 25103 19579 25109
rect 38286 25100 38292 25112
rect 38344 25100 38350 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 4709 24939 4767 24945
rect 4709 24905 4721 24939
rect 4755 24936 4767 24939
rect 4982 24936 4988 24948
rect 4755 24908 4988 24936
rect 4755 24905 4767 24908
rect 4709 24899 4767 24905
rect 4982 24896 4988 24908
rect 5040 24896 5046 24948
rect 9858 24936 9864 24948
rect 9819 24908 9864 24936
rect 9858 24896 9864 24908
rect 9916 24896 9922 24948
rect 11606 24936 11612 24948
rect 10428 24908 11612 24936
rect 10428 24868 10456 24908
rect 11606 24896 11612 24908
rect 11664 24896 11670 24948
rect 11808 24908 12112 24936
rect 7668 24840 8156 24868
rect 1578 24800 1584 24812
rect 1539 24772 1584 24800
rect 1578 24760 1584 24772
rect 1636 24800 1642 24812
rect 2225 24803 2283 24809
rect 2225 24800 2237 24803
rect 1636 24772 2237 24800
rect 1636 24760 1642 24772
rect 2225 24769 2237 24772
rect 2271 24769 2283 24803
rect 2866 24800 2872 24812
rect 2827 24772 2872 24800
rect 2225 24763 2283 24769
rect 2866 24760 2872 24772
rect 2924 24800 2930 24812
rect 3326 24800 3332 24812
rect 2924 24772 3332 24800
rect 2924 24760 2930 24772
rect 3326 24760 3332 24772
rect 3384 24800 3390 24812
rect 3421 24803 3479 24809
rect 3421 24800 3433 24803
rect 3384 24772 3433 24800
rect 3384 24760 3390 24772
rect 3421 24769 3433 24772
rect 3467 24769 3479 24803
rect 3421 24763 3479 24769
rect 4890 24760 4896 24812
rect 4948 24800 4954 24812
rect 5721 24803 5779 24809
rect 5721 24800 5733 24803
rect 4948 24772 5733 24800
rect 4948 24760 4954 24772
rect 5721 24769 5733 24772
rect 5767 24769 5779 24803
rect 5721 24763 5779 24769
rect 6454 24760 6460 24812
rect 6512 24800 6518 24812
rect 6549 24803 6607 24809
rect 6549 24800 6561 24803
rect 6512 24772 6561 24800
rect 6512 24760 6518 24772
rect 6549 24769 6561 24772
rect 6595 24769 6607 24803
rect 6549 24763 6607 24769
rect 6730 24760 6736 24812
rect 6788 24800 6794 24812
rect 7668 24800 7696 24840
rect 7834 24800 7840 24812
rect 6788 24772 7696 24800
rect 7795 24772 7840 24800
rect 6788 24760 6794 24772
rect 7834 24760 7840 24772
rect 7892 24760 7898 24812
rect 7926 24760 7932 24812
rect 7984 24800 7990 24812
rect 8128 24800 8156 24840
rect 9646 24840 10456 24868
rect 8481 24803 8539 24809
rect 8481 24800 8493 24803
rect 7984 24772 8029 24800
rect 8128 24772 8493 24800
rect 7984 24760 7990 24772
rect 8481 24769 8493 24772
rect 8527 24800 8539 24803
rect 8662 24800 8668 24812
rect 8527 24772 8668 24800
rect 8527 24769 8539 24772
rect 8481 24763 8539 24769
rect 8662 24760 8668 24772
rect 8720 24760 8726 24812
rect 8846 24760 8852 24812
rect 8904 24800 8910 24812
rect 9125 24803 9183 24809
rect 9125 24800 9137 24803
rect 8904 24772 9137 24800
rect 8904 24760 8910 24772
rect 9125 24769 9137 24772
rect 9171 24769 9183 24803
rect 9125 24763 9183 24769
rect 9217 24803 9275 24809
rect 9217 24769 9229 24803
rect 9263 24800 9275 24803
rect 9646 24800 9674 24840
rect 10502 24828 10508 24880
rect 10560 24868 10566 24880
rect 11808 24877 11836 24908
rect 10597 24871 10655 24877
rect 10597 24868 10609 24871
rect 10560 24840 10609 24868
rect 10560 24828 10566 24840
rect 10597 24837 10609 24840
rect 10643 24837 10655 24871
rect 10597 24831 10655 24837
rect 11793 24871 11851 24877
rect 11793 24837 11805 24871
rect 11839 24837 11851 24871
rect 11793 24831 11851 24837
rect 11882 24828 11888 24880
rect 11940 24868 11946 24880
rect 12084 24868 12112 24908
rect 12158 24896 12164 24948
rect 12216 24936 12222 24948
rect 13906 24936 13912 24948
rect 12216 24908 13912 24936
rect 12216 24896 12222 24908
rect 13906 24896 13912 24908
rect 13964 24896 13970 24948
rect 15930 24936 15936 24948
rect 14108 24908 15936 24936
rect 12618 24868 12624 24880
rect 11940 24840 11985 24868
rect 12084 24840 12624 24868
rect 11940 24828 11946 24840
rect 12618 24828 12624 24840
rect 12676 24828 12682 24880
rect 13081 24871 13139 24877
rect 13081 24868 13093 24871
rect 12820 24840 13093 24868
rect 9263 24772 9674 24800
rect 9769 24803 9827 24809
rect 9263 24769 9275 24772
rect 9217 24763 9275 24769
rect 9769 24769 9781 24803
rect 9815 24800 9827 24803
rect 10318 24800 10324 24812
rect 9815 24772 10324 24800
rect 9815 24769 9827 24772
rect 9769 24763 9827 24769
rect 10318 24760 10324 24772
rect 10376 24760 10382 24812
rect 12526 24760 12532 24812
rect 12584 24800 12590 24812
rect 12820 24800 12848 24840
rect 13081 24837 13093 24840
rect 13127 24837 13139 24871
rect 13081 24831 13139 24837
rect 12584 24772 12848 24800
rect 13633 24803 13691 24809
rect 12584 24760 12590 24772
rect 13633 24769 13645 24803
rect 13679 24800 13691 24803
rect 13814 24800 13820 24812
rect 13679 24772 13820 24800
rect 13679 24769 13691 24772
rect 13633 24763 13691 24769
rect 13814 24760 13820 24772
rect 13872 24760 13878 24812
rect 5813 24735 5871 24741
rect 5813 24701 5825 24735
rect 5859 24732 5871 24735
rect 9306 24732 9312 24744
rect 5859 24704 9312 24732
rect 5859 24701 5871 24704
rect 5813 24695 5871 24701
rect 9306 24692 9312 24704
rect 9364 24692 9370 24744
rect 10042 24692 10048 24744
rect 10100 24732 10106 24744
rect 10505 24735 10563 24741
rect 10505 24732 10517 24735
rect 10100 24704 10517 24732
rect 10100 24692 10106 24704
rect 10505 24701 10517 24704
rect 10551 24701 10563 24735
rect 10505 24695 10563 24701
rect 11149 24735 11207 24741
rect 11149 24701 11161 24735
rect 11195 24732 11207 24735
rect 12158 24732 12164 24744
rect 11195 24704 12164 24732
rect 11195 24701 11207 24704
rect 11149 24695 11207 24701
rect 12158 24692 12164 24704
rect 12216 24692 12222 24744
rect 12989 24735 13047 24741
rect 12989 24732 13001 24735
rect 12268 24704 13001 24732
rect 1765 24667 1823 24673
rect 1765 24633 1777 24667
rect 1811 24664 1823 24667
rect 1946 24664 1952 24676
rect 1811 24636 1952 24664
rect 1811 24633 1823 24636
rect 1765 24627 1823 24633
rect 1946 24624 1952 24636
rect 2004 24664 2010 24676
rect 5626 24664 5632 24676
rect 2004 24636 5632 24664
rect 2004 24624 2010 24636
rect 5626 24624 5632 24636
rect 5684 24624 5690 24676
rect 6641 24667 6699 24673
rect 6641 24633 6653 24667
rect 6687 24664 6699 24667
rect 8573 24667 8631 24673
rect 6687 24636 8064 24664
rect 6687 24633 6699 24636
rect 6641 24627 6699 24633
rect 3418 24556 3424 24608
rect 3476 24596 3482 24608
rect 4157 24599 4215 24605
rect 4157 24596 4169 24599
rect 3476 24568 4169 24596
rect 3476 24556 3482 24568
rect 4157 24565 4169 24568
rect 4203 24596 4215 24599
rect 4614 24596 4620 24608
rect 4203 24568 4620 24596
rect 4203 24565 4215 24568
rect 4157 24559 4215 24565
rect 4614 24556 4620 24568
rect 4672 24596 4678 24608
rect 5169 24599 5227 24605
rect 5169 24596 5181 24599
rect 4672 24568 5181 24596
rect 4672 24556 4678 24568
rect 5169 24565 5181 24568
rect 5215 24565 5227 24599
rect 5169 24559 5227 24565
rect 7377 24599 7435 24605
rect 7377 24565 7389 24599
rect 7423 24596 7435 24599
rect 7926 24596 7932 24608
rect 7423 24568 7932 24596
rect 7423 24565 7435 24568
rect 7377 24559 7435 24565
rect 7926 24556 7932 24568
rect 7984 24556 7990 24608
rect 8036 24596 8064 24636
rect 8573 24633 8585 24667
rect 8619 24664 8631 24667
rect 8619 24636 9674 24664
rect 8619 24633 8631 24636
rect 8573 24627 8631 24633
rect 9490 24596 9496 24608
rect 8036 24568 9496 24596
rect 9490 24556 9496 24568
rect 9548 24556 9554 24608
rect 9646 24596 9674 24636
rect 10594 24624 10600 24676
rect 10652 24664 10658 24676
rect 12268 24664 12296 24704
rect 12989 24701 13001 24704
rect 13035 24701 13047 24735
rect 14108 24732 14136 24908
rect 15930 24896 15936 24908
rect 15988 24936 15994 24948
rect 16482 24936 16488 24948
rect 15988 24908 16488 24936
rect 15988 24896 15994 24908
rect 16482 24896 16488 24908
rect 16540 24896 16546 24948
rect 18325 24939 18383 24945
rect 18325 24905 18337 24939
rect 18371 24936 18383 24939
rect 18506 24936 18512 24948
rect 18371 24908 18512 24936
rect 18371 24905 18383 24908
rect 18325 24899 18383 24905
rect 18506 24896 18512 24908
rect 18564 24896 18570 24948
rect 20162 24936 20168 24948
rect 18708 24908 20168 24936
rect 14366 24828 14372 24880
rect 14424 24868 14430 24880
rect 14461 24871 14519 24877
rect 14461 24868 14473 24871
rect 14424 24840 14473 24868
rect 14424 24828 14430 24840
rect 14461 24837 14473 24840
rect 14507 24837 14519 24871
rect 18708 24868 18736 24908
rect 20162 24896 20168 24908
rect 20220 24896 20226 24948
rect 22738 24936 22744 24948
rect 22699 24908 22744 24936
rect 22738 24896 22744 24908
rect 22796 24896 22802 24948
rect 23106 24896 23112 24948
rect 23164 24936 23170 24948
rect 23201 24939 23259 24945
rect 23201 24936 23213 24939
rect 23164 24908 23213 24936
rect 23164 24896 23170 24908
rect 23201 24905 23213 24908
rect 23247 24905 23259 24939
rect 23201 24899 23259 24905
rect 19429 24871 19487 24877
rect 19429 24868 19441 24871
rect 14461 24831 14519 24837
rect 16546 24840 18736 24868
rect 18892 24840 19441 24868
rect 15654 24760 15660 24812
rect 15712 24800 15718 24812
rect 16301 24803 16359 24809
rect 16301 24800 16313 24803
rect 15712 24772 16313 24800
rect 15712 24760 15718 24772
rect 16301 24769 16313 24772
rect 16347 24800 16359 24803
rect 16390 24800 16396 24812
rect 16347 24772 16396 24800
rect 16347 24769 16359 24772
rect 16301 24763 16359 24769
rect 16390 24760 16396 24772
rect 16448 24760 16454 24812
rect 14366 24732 14372 24744
rect 12989 24695 13047 24701
rect 13372 24704 14136 24732
rect 14327 24704 14372 24732
rect 10652 24636 12296 24664
rect 12345 24667 12403 24673
rect 10652 24624 10658 24636
rect 12345 24633 12357 24667
rect 12391 24664 12403 24667
rect 13372 24664 13400 24704
rect 14366 24692 14372 24704
rect 14424 24692 14430 24744
rect 15381 24735 15439 24741
rect 15381 24701 15393 24735
rect 15427 24732 15439 24735
rect 15562 24732 15568 24744
rect 15427 24704 15568 24732
rect 15427 24701 15439 24704
rect 15381 24695 15439 24701
rect 15562 24692 15568 24704
rect 15620 24732 15626 24744
rect 16546 24732 16574 24840
rect 17586 24800 17592 24812
rect 17547 24772 17592 24800
rect 17586 24760 17592 24772
rect 17644 24760 17650 24812
rect 18138 24760 18144 24812
rect 18196 24800 18202 24812
rect 18417 24803 18475 24809
rect 18417 24800 18429 24803
rect 18196 24772 18429 24800
rect 18196 24760 18202 24772
rect 18417 24769 18429 24772
rect 18463 24769 18475 24803
rect 18417 24763 18475 24769
rect 15620 24704 16574 24732
rect 17129 24735 17187 24741
rect 15620 24692 15626 24704
rect 17129 24701 17141 24735
rect 17175 24732 17187 24735
rect 17310 24732 17316 24744
rect 17175 24704 17316 24732
rect 17175 24701 17187 24704
rect 17129 24695 17187 24701
rect 17310 24692 17316 24704
rect 17368 24692 17374 24744
rect 17681 24735 17739 24741
rect 17681 24701 17693 24735
rect 17727 24732 17739 24735
rect 18892 24732 18920 24840
rect 19429 24837 19441 24840
rect 19475 24837 19487 24871
rect 20257 24871 20315 24877
rect 20257 24868 20269 24871
rect 19429 24831 19487 24837
rect 19996 24840 20269 24868
rect 19886 24760 19892 24812
rect 19944 24800 19950 24812
rect 19996 24800 20024 24840
rect 20257 24837 20269 24840
rect 20303 24837 20315 24871
rect 20257 24831 20315 24837
rect 21266 24800 21272 24812
rect 19944 24772 20024 24800
rect 21227 24772 21272 24800
rect 19944 24760 19950 24772
rect 21266 24760 21272 24772
rect 21324 24760 21330 24812
rect 21358 24760 21364 24812
rect 21416 24800 21422 24812
rect 21416 24772 21461 24800
rect 21416 24760 21422 24772
rect 21542 24760 21548 24812
rect 21600 24800 21606 24812
rect 29549 24803 29607 24809
rect 29549 24800 29561 24803
rect 21600 24772 29561 24800
rect 21600 24760 21606 24772
rect 29549 24769 29561 24772
rect 29595 24769 29607 24803
rect 29549 24763 29607 24769
rect 17727 24704 18920 24732
rect 17727 24701 17739 24704
rect 17681 24695 17739 24701
rect 19426 24692 19432 24744
rect 19484 24732 19490 24744
rect 19521 24735 19579 24741
rect 19521 24732 19533 24735
rect 19484 24704 19533 24732
rect 19484 24692 19490 24704
rect 19521 24701 19533 24704
rect 19567 24701 19579 24735
rect 19521 24695 19579 24701
rect 20165 24735 20223 24741
rect 20165 24701 20177 24735
rect 20211 24732 20223 24735
rect 20254 24732 20260 24744
rect 20211 24704 20260 24732
rect 20211 24701 20223 24704
rect 20165 24695 20223 24701
rect 20254 24692 20260 24704
rect 20312 24732 20318 24744
rect 20312 24704 20852 24732
rect 20312 24692 20318 24704
rect 12391 24636 13400 24664
rect 12391 24633 12403 24636
rect 12345 24627 12403 24633
rect 13906 24624 13912 24676
rect 13964 24664 13970 24676
rect 16298 24664 16304 24676
rect 13964 24636 16304 24664
rect 13964 24624 13970 24636
rect 16298 24624 16304 24636
rect 16356 24624 16362 24676
rect 17218 24624 17224 24676
rect 17276 24664 17282 24676
rect 18969 24667 19027 24673
rect 18969 24664 18981 24667
rect 17276 24636 18981 24664
rect 17276 24624 17282 24636
rect 18969 24633 18981 24636
rect 19015 24633 19027 24667
rect 18969 24627 19027 24633
rect 20070 24624 20076 24676
rect 20128 24664 20134 24676
rect 20714 24664 20720 24676
rect 20128 24636 20720 24664
rect 20128 24624 20134 24636
rect 20714 24624 20720 24636
rect 20772 24624 20778 24676
rect 20824 24664 20852 24704
rect 21910 24692 21916 24744
rect 21968 24732 21974 24744
rect 22005 24735 22063 24741
rect 22005 24732 22017 24735
rect 21968 24704 22017 24732
rect 21968 24692 21974 24704
rect 22005 24701 22017 24704
rect 22051 24701 22063 24735
rect 30006 24732 30012 24744
rect 22005 24695 22063 24701
rect 22480 24704 30012 24732
rect 22480 24664 22508 24704
rect 30006 24692 30012 24704
rect 30064 24692 30070 24744
rect 37918 24692 37924 24744
rect 37976 24732 37982 24744
rect 38013 24735 38071 24741
rect 38013 24732 38025 24735
rect 37976 24704 38025 24732
rect 37976 24692 37982 24704
rect 38013 24701 38025 24704
rect 38059 24701 38071 24735
rect 38286 24732 38292 24744
rect 38247 24704 38292 24732
rect 38013 24695 38071 24701
rect 38286 24692 38292 24704
rect 38344 24692 38350 24744
rect 23753 24667 23811 24673
rect 23753 24664 23765 24667
rect 20824 24636 22508 24664
rect 22572 24636 23765 24664
rect 11790 24596 11796 24608
rect 9646 24568 11796 24596
rect 11790 24556 11796 24568
rect 11848 24556 11854 24608
rect 14182 24556 14188 24608
rect 14240 24596 14246 24608
rect 15562 24596 15568 24608
rect 14240 24568 15568 24596
rect 14240 24556 14246 24568
rect 15562 24556 15568 24568
rect 15620 24556 15626 24608
rect 15746 24556 15752 24608
rect 15804 24596 15810 24608
rect 16206 24596 16212 24608
rect 15804 24568 16212 24596
rect 15804 24556 15810 24568
rect 16206 24556 16212 24568
rect 16264 24556 16270 24608
rect 17586 24556 17592 24608
rect 17644 24596 17650 24608
rect 22572 24596 22600 24636
rect 23753 24633 23765 24636
rect 23799 24633 23811 24667
rect 23753 24627 23811 24633
rect 17644 24568 22600 24596
rect 29641 24599 29699 24605
rect 17644 24556 17650 24568
rect 29641 24565 29653 24599
rect 29687 24596 29699 24599
rect 36538 24596 36544 24608
rect 29687 24568 36544 24596
rect 29687 24565 29699 24568
rect 29641 24559 29699 24565
rect 36538 24556 36544 24568
rect 36596 24556 36602 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 1670 24392 1676 24404
rect 1583 24364 1676 24392
rect 1670 24352 1676 24364
rect 1728 24392 1734 24404
rect 2590 24392 2596 24404
rect 1728 24364 2596 24392
rect 1728 24352 1734 24364
rect 2590 24352 2596 24364
rect 2648 24352 2654 24404
rect 3326 24392 3332 24404
rect 3287 24364 3332 24392
rect 3326 24352 3332 24364
rect 3384 24392 3390 24404
rect 3878 24392 3884 24404
rect 3384 24364 3884 24392
rect 3384 24352 3390 24364
rect 3878 24352 3884 24364
rect 3936 24392 3942 24404
rect 4893 24395 4951 24401
rect 4893 24392 4905 24395
rect 3936 24364 4905 24392
rect 3936 24352 3942 24364
rect 4893 24361 4905 24364
rect 4939 24361 4951 24395
rect 4893 24355 4951 24361
rect 6822 24352 6828 24404
rect 6880 24392 6886 24404
rect 7101 24395 7159 24401
rect 7101 24392 7113 24395
rect 6880 24364 7113 24392
rect 6880 24352 6886 24364
rect 7101 24361 7113 24364
rect 7147 24361 7159 24395
rect 7101 24355 7159 24361
rect 8481 24395 8539 24401
rect 8481 24361 8493 24395
rect 8527 24392 8539 24395
rect 10502 24392 10508 24404
rect 8527 24364 10508 24392
rect 8527 24361 8539 24364
rect 8481 24355 8539 24361
rect 10502 24352 10508 24364
rect 10560 24352 10566 24404
rect 13722 24352 13728 24404
rect 13780 24392 13786 24404
rect 15838 24392 15844 24404
rect 13780 24364 15844 24392
rect 13780 24352 13786 24364
rect 15838 24352 15844 24364
rect 15896 24352 15902 24404
rect 16390 24352 16396 24404
rect 16448 24392 16454 24404
rect 23017 24395 23075 24401
rect 23017 24392 23029 24395
rect 16448 24364 23029 24392
rect 16448 24352 16454 24364
rect 23017 24361 23029 24364
rect 23063 24361 23075 24395
rect 33594 24392 33600 24404
rect 33555 24364 33600 24392
rect 23017 24355 23075 24361
rect 33594 24352 33600 24364
rect 33652 24352 33658 24404
rect 2222 24324 2228 24336
rect 2183 24296 2228 24324
rect 2222 24284 2228 24296
rect 2280 24324 2286 24336
rect 5445 24327 5503 24333
rect 5445 24324 5457 24327
rect 2280 24296 5457 24324
rect 2280 24284 2286 24296
rect 5445 24293 5457 24296
rect 5491 24324 5503 24327
rect 5902 24324 5908 24336
rect 5491 24296 5908 24324
rect 5491 24293 5503 24296
rect 5445 24287 5503 24293
rect 5902 24284 5908 24296
rect 5960 24284 5966 24336
rect 9309 24327 9367 24333
rect 9309 24293 9321 24327
rect 9355 24324 9367 24327
rect 11882 24324 11888 24336
rect 9355 24296 11888 24324
rect 9355 24293 9367 24296
rect 9309 24287 9367 24293
rect 11882 24284 11888 24296
rect 11940 24284 11946 24336
rect 12618 24284 12624 24336
rect 12676 24324 12682 24336
rect 14918 24324 14924 24336
rect 12676 24296 14924 24324
rect 12676 24284 12682 24296
rect 14918 24284 14924 24296
rect 14976 24284 14982 24336
rect 15289 24327 15347 24333
rect 15289 24293 15301 24327
rect 15335 24324 15347 24327
rect 16758 24324 16764 24336
rect 15335 24296 16764 24324
rect 15335 24293 15347 24296
rect 15289 24287 15347 24293
rect 5718 24216 5724 24268
rect 5776 24256 5782 24268
rect 5776 24228 7788 24256
rect 5776 24216 5782 24228
rect 7760 24197 7788 24228
rect 7926 24216 7932 24268
rect 7984 24256 7990 24268
rect 9674 24256 9680 24268
rect 7984 24228 9680 24256
rect 7984 24216 7990 24228
rect 9674 24216 9680 24228
rect 9732 24216 9738 24268
rect 10229 24259 10287 24265
rect 10229 24225 10241 24259
rect 10275 24256 10287 24259
rect 10410 24256 10416 24268
rect 10275 24228 10416 24256
rect 10275 24225 10287 24228
rect 10229 24219 10287 24225
rect 10410 24216 10416 24228
rect 10468 24216 10474 24268
rect 10505 24259 10563 24265
rect 10505 24225 10517 24259
rect 10551 24256 10563 24259
rect 12158 24256 12164 24268
rect 10551 24228 12164 24256
rect 10551 24225 10563 24228
rect 10505 24219 10563 24225
rect 12158 24216 12164 24228
rect 12216 24216 12222 24268
rect 12345 24259 12403 24265
rect 12345 24225 12357 24259
rect 12391 24256 12403 24259
rect 13814 24256 13820 24268
rect 12391 24228 13820 24256
rect 12391 24225 12403 24228
rect 12345 24219 12403 24225
rect 13814 24216 13820 24228
rect 13872 24216 13878 24268
rect 14274 24216 14280 24268
rect 14332 24256 14338 24268
rect 15304 24256 15332 24287
rect 16758 24284 16764 24296
rect 16816 24284 16822 24336
rect 24026 24324 24032 24336
rect 17420 24296 24032 24324
rect 14332 24228 15332 24256
rect 14332 24216 14338 24228
rect 16390 24216 16396 24268
rect 16448 24256 16454 24268
rect 17420 24265 17448 24296
rect 24026 24284 24032 24296
rect 24084 24284 24090 24336
rect 17405 24259 17463 24265
rect 17405 24256 17417 24259
rect 16448 24228 17417 24256
rect 16448 24216 16454 24228
rect 17405 24225 17417 24228
rect 17451 24225 17463 24259
rect 17405 24219 17463 24225
rect 19242 24216 19248 24268
rect 19300 24256 19306 24268
rect 20717 24259 20775 24265
rect 20717 24256 20729 24259
rect 19300 24228 20729 24256
rect 19300 24216 19306 24228
rect 20717 24225 20729 24228
rect 20763 24225 20775 24259
rect 21266 24256 21272 24268
rect 21227 24228 21272 24256
rect 20717 24219 20775 24225
rect 21266 24216 21272 24228
rect 21324 24216 21330 24268
rect 21910 24256 21916 24268
rect 21871 24228 21916 24256
rect 21910 24216 21916 24228
rect 21968 24216 21974 24268
rect 22186 24256 22192 24268
rect 22147 24228 22192 24256
rect 22186 24216 22192 24228
rect 22244 24216 22250 24268
rect 7285 24191 7343 24197
rect 7285 24157 7297 24191
rect 7331 24157 7343 24191
rect 7285 24151 7343 24157
rect 7745 24191 7803 24197
rect 7745 24157 7757 24191
rect 7791 24157 7803 24191
rect 8386 24188 8392 24200
rect 8347 24160 8392 24188
rect 7745 24151 7803 24157
rect 6089 24123 6147 24129
rect 6089 24089 6101 24123
rect 6135 24120 6147 24123
rect 7300 24120 7328 24151
rect 8386 24148 8392 24160
rect 8444 24148 8450 24200
rect 8938 24148 8944 24200
rect 8996 24188 9002 24200
rect 9217 24191 9275 24197
rect 9217 24188 9229 24191
rect 8996 24160 9229 24188
rect 8996 24148 9002 24160
rect 9217 24157 9229 24160
rect 9263 24157 9275 24191
rect 9217 24151 9275 24157
rect 10962 24148 10968 24200
rect 11020 24188 11026 24200
rect 11057 24191 11115 24197
rect 11057 24188 11069 24191
rect 11020 24160 11069 24188
rect 11020 24148 11026 24160
rect 11057 24157 11069 24160
rect 11103 24157 11115 24191
rect 11057 24151 11115 24157
rect 19058 24148 19064 24200
rect 19116 24188 19122 24200
rect 19429 24191 19487 24197
rect 19429 24188 19441 24191
rect 19116 24160 19441 24188
rect 19116 24148 19122 24160
rect 19429 24157 19441 24160
rect 19475 24188 19487 24191
rect 19981 24191 20039 24197
rect 19981 24188 19993 24191
rect 19475 24160 19993 24188
rect 19475 24157 19487 24160
rect 19429 24151 19487 24157
rect 19981 24157 19993 24160
rect 20027 24157 20039 24191
rect 19981 24151 20039 24157
rect 20346 24148 20352 24200
rect 20404 24188 20410 24200
rect 20809 24191 20867 24197
rect 20809 24188 20821 24191
rect 20404 24160 20821 24188
rect 20404 24148 20410 24160
rect 20809 24157 20821 24160
rect 20855 24157 20867 24191
rect 20809 24151 20867 24157
rect 27246 24148 27252 24200
rect 27304 24188 27310 24200
rect 33781 24191 33839 24197
rect 33781 24188 33793 24191
rect 27304 24160 33793 24188
rect 27304 24148 27310 24160
rect 33781 24157 33793 24160
rect 33827 24188 33839 24191
rect 34241 24191 34299 24197
rect 34241 24188 34253 24191
rect 33827 24160 34253 24188
rect 33827 24157 33839 24160
rect 33781 24151 33839 24157
rect 34241 24157 34253 24160
rect 34287 24188 34299 24191
rect 37826 24188 37832 24200
rect 34287 24160 35894 24188
rect 37787 24160 37832 24188
rect 34287 24157 34299 24160
rect 34241 24151 34299 24157
rect 6135 24092 10088 24120
rect 6135 24089 6147 24092
rect 6089 24083 6147 24089
rect 2685 24055 2743 24061
rect 2685 24021 2697 24055
rect 2731 24052 2743 24055
rect 2866 24052 2872 24064
rect 2731 24024 2872 24052
rect 2731 24021 2743 24024
rect 2685 24015 2743 24021
rect 2866 24012 2872 24024
rect 2924 24012 2930 24064
rect 4341 24055 4399 24061
rect 4341 24021 4353 24055
rect 4387 24052 4399 24055
rect 4614 24052 4620 24064
rect 4387 24024 4620 24052
rect 4387 24021 4399 24024
rect 4341 24015 4399 24021
rect 4614 24012 4620 24024
rect 4672 24012 4678 24064
rect 6638 24052 6644 24064
rect 6599 24024 6644 24052
rect 6638 24012 6644 24024
rect 6696 24012 6702 24064
rect 7837 24055 7895 24061
rect 7837 24021 7849 24055
rect 7883 24052 7895 24055
rect 9950 24052 9956 24064
rect 7883 24024 9956 24052
rect 7883 24021 7895 24024
rect 7837 24015 7895 24021
rect 9950 24012 9956 24024
rect 10008 24012 10014 24064
rect 10060 24052 10088 24092
rect 10134 24080 10140 24132
rect 10192 24120 10198 24132
rect 10413 24123 10471 24129
rect 10413 24120 10425 24123
rect 10192 24092 10425 24120
rect 10192 24080 10198 24092
rect 10413 24089 10425 24092
rect 10459 24089 10471 24123
rect 11330 24120 11336 24132
rect 10413 24083 10471 24089
rect 10520 24092 11336 24120
rect 10520 24052 10548 24092
rect 11330 24080 11336 24092
rect 11388 24080 11394 24132
rect 11422 24080 11428 24132
rect 11480 24120 11486 24132
rect 11701 24123 11759 24129
rect 11701 24120 11713 24123
rect 11480 24092 11713 24120
rect 11480 24080 11486 24092
rect 11701 24089 11713 24092
rect 11747 24089 11759 24123
rect 12250 24120 12256 24132
rect 12211 24092 12256 24120
rect 11701 24083 11759 24089
rect 12250 24080 12256 24092
rect 12308 24080 12314 24132
rect 13078 24120 13084 24132
rect 13039 24092 13084 24120
rect 13078 24080 13084 24092
rect 13136 24080 13142 24132
rect 13173 24123 13231 24129
rect 13173 24089 13185 24123
rect 13219 24089 13231 24123
rect 13173 24083 13231 24089
rect 10060 24024 10548 24052
rect 11149 24055 11207 24061
rect 11149 24021 11161 24055
rect 11195 24052 11207 24055
rect 13188 24052 13216 24083
rect 13262 24080 13268 24132
rect 13320 24120 13326 24132
rect 13725 24123 13783 24129
rect 13725 24120 13737 24123
rect 13320 24092 13737 24120
rect 13320 24080 13326 24092
rect 13725 24089 13737 24092
rect 13771 24089 13783 24123
rect 14734 24120 14740 24132
rect 14695 24092 14740 24120
rect 13725 24083 13783 24089
rect 14734 24080 14740 24092
rect 14792 24080 14798 24132
rect 14826 24080 14832 24132
rect 14884 24120 14890 24132
rect 14884 24092 14929 24120
rect 14884 24080 14890 24092
rect 15838 24080 15844 24132
rect 15896 24120 15902 24132
rect 16393 24123 16451 24129
rect 16393 24120 16405 24123
rect 15896 24092 16405 24120
rect 15896 24080 15902 24092
rect 16393 24089 16405 24092
rect 16439 24089 16451 24123
rect 16393 24083 16451 24089
rect 16485 24123 16543 24129
rect 16485 24089 16497 24123
rect 16531 24089 16543 24123
rect 18598 24120 18604 24132
rect 18559 24092 18604 24120
rect 16485 24083 16543 24089
rect 11195 24024 13216 24052
rect 11195 24021 11207 24024
rect 11149 24015 11207 24021
rect 13538 24012 13544 24064
rect 13596 24052 13602 24064
rect 16500 24052 16528 24083
rect 18598 24080 18604 24092
rect 18656 24080 18662 24132
rect 19886 24080 19892 24132
rect 19944 24120 19950 24132
rect 20073 24123 20131 24129
rect 20073 24120 20085 24123
rect 19944 24092 20085 24120
rect 19944 24080 19950 24092
rect 20073 24089 20085 24092
rect 20119 24089 20131 24123
rect 20073 24083 20131 24089
rect 21174 24080 21180 24132
rect 21232 24120 21238 24132
rect 22005 24123 22063 24129
rect 22005 24120 22017 24123
rect 21232 24092 22017 24120
rect 21232 24080 21238 24092
rect 22005 24089 22017 24092
rect 22051 24089 22063 24123
rect 22005 24083 22063 24089
rect 13596 24024 16528 24052
rect 13596 24012 13602 24024
rect 16574 24012 16580 24064
rect 16632 24052 16638 24064
rect 17957 24055 18015 24061
rect 17957 24052 17969 24055
rect 16632 24024 17969 24052
rect 16632 24012 16638 24024
rect 17957 24021 17969 24024
rect 18003 24021 18015 24055
rect 18506 24052 18512 24064
rect 18467 24024 18512 24052
rect 17957 24015 18015 24021
rect 18506 24012 18512 24024
rect 18564 24012 18570 24064
rect 35866 24052 35894 24160
rect 37826 24148 37832 24160
rect 37884 24148 37890 24200
rect 37550 24052 37556 24064
rect 35866 24024 37556 24052
rect 37550 24012 37556 24024
rect 37608 24012 37614 24064
rect 38010 24052 38016 24064
rect 37971 24024 38016 24052
rect 38010 24012 38016 24024
rect 38068 24012 38074 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 2222 23808 2228 23860
rect 2280 23848 2286 23860
rect 2409 23851 2467 23857
rect 2409 23848 2421 23851
rect 2280 23820 2421 23848
rect 2280 23808 2286 23820
rect 2409 23817 2421 23820
rect 2455 23848 2467 23851
rect 2961 23851 3019 23857
rect 2961 23848 2973 23851
rect 2455 23820 2973 23848
rect 2455 23817 2467 23820
rect 2409 23811 2467 23817
rect 2961 23817 2973 23820
rect 3007 23848 3019 23851
rect 3234 23848 3240 23860
rect 3007 23820 3240 23848
rect 3007 23817 3019 23820
rect 2961 23811 3019 23817
rect 3234 23808 3240 23820
rect 3292 23808 3298 23860
rect 3878 23848 3884 23860
rect 3839 23820 3884 23848
rect 3878 23808 3884 23820
rect 3936 23848 3942 23860
rect 5169 23851 5227 23857
rect 5169 23848 5181 23851
rect 3936 23820 5181 23848
rect 3936 23808 3942 23820
rect 5169 23817 5181 23820
rect 5215 23817 5227 23851
rect 5902 23848 5908 23860
rect 5863 23820 5908 23848
rect 5169 23811 5227 23817
rect 5902 23808 5908 23820
rect 5960 23808 5966 23860
rect 7837 23851 7895 23857
rect 7837 23817 7849 23851
rect 7883 23848 7895 23851
rect 10134 23848 10140 23860
rect 7883 23820 10140 23848
rect 7883 23817 7895 23820
rect 7837 23811 7895 23817
rect 10134 23808 10140 23820
rect 10192 23808 10198 23860
rect 10962 23848 10968 23860
rect 10336 23820 10968 23848
rect 6638 23740 6644 23792
rect 6696 23780 6702 23792
rect 6696 23752 8248 23780
rect 6696 23740 6702 23752
rect 1946 23712 1952 23724
rect 1907 23684 1952 23712
rect 1946 23672 1952 23684
rect 2004 23672 2010 23724
rect 3602 23672 3608 23724
rect 3660 23712 3666 23724
rect 7745 23715 7803 23721
rect 7745 23712 7757 23715
rect 3660 23684 7757 23712
rect 3660 23672 3666 23684
rect 7745 23681 7757 23684
rect 7791 23681 7803 23715
rect 8220 23712 8248 23752
rect 8294 23740 8300 23792
rect 8352 23780 8358 23792
rect 10336 23780 10364 23820
rect 10962 23808 10968 23820
rect 11020 23808 11026 23860
rect 11057 23851 11115 23857
rect 11057 23817 11069 23851
rect 11103 23848 11115 23851
rect 12434 23848 12440 23860
rect 11103 23820 12440 23848
rect 11103 23817 11115 23820
rect 11057 23811 11115 23817
rect 12434 23808 12440 23820
rect 12492 23808 12498 23860
rect 14826 23848 14832 23860
rect 12544 23820 14832 23848
rect 8352 23752 10364 23780
rect 8352 23740 8358 23752
rect 9033 23715 9091 23721
rect 9033 23712 9045 23715
rect 8220 23684 9045 23712
rect 7745 23675 7803 23681
rect 9033 23681 9045 23684
rect 9079 23681 9091 23715
rect 9674 23712 9680 23724
rect 9635 23684 9680 23712
rect 9033 23675 9091 23681
rect 9674 23672 9680 23684
rect 9732 23672 9738 23724
rect 10336 23721 10364 23752
rect 10413 23783 10471 23789
rect 10413 23749 10425 23783
rect 10459 23780 10471 23783
rect 12544 23780 12572 23820
rect 14826 23808 14832 23820
rect 14884 23808 14890 23860
rect 18598 23808 18604 23860
rect 18656 23848 18662 23860
rect 21726 23848 21732 23860
rect 18656 23820 21732 23848
rect 18656 23808 18662 23820
rect 21726 23808 21732 23820
rect 21784 23848 21790 23860
rect 22005 23851 22063 23857
rect 22005 23848 22017 23851
rect 21784 23820 22017 23848
rect 21784 23808 21790 23820
rect 22005 23817 22017 23820
rect 22051 23817 22063 23851
rect 26234 23848 26240 23860
rect 26195 23820 26240 23848
rect 22005 23811 22063 23817
rect 26234 23808 26240 23820
rect 26292 23808 26298 23860
rect 27246 23848 27252 23860
rect 27207 23820 27252 23848
rect 27246 23808 27252 23820
rect 27304 23808 27310 23860
rect 30006 23848 30012 23860
rect 29967 23820 30012 23848
rect 30006 23808 30012 23820
rect 30064 23808 30070 23860
rect 12710 23780 12716 23792
rect 10459 23752 12572 23780
rect 12671 23752 12716 23780
rect 10459 23749 10471 23752
rect 10413 23743 10471 23749
rect 12710 23740 12716 23752
rect 12768 23740 12774 23792
rect 13265 23783 13323 23789
rect 13265 23749 13277 23783
rect 13311 23780 13323 23783
rect 13446 23780 13452 23792
rect 13311 23752 13452 23780
rect 13311 23749 13323 23752
rect 13265 23743 13323 23749
rect 13446 23740 13452 23752
rect 13504 23740 13510 23792
rect 13538 23740 13544 23792
rect 13596 23780 13602 23792
rect 13909 23783 13967 23789
rect 13909 23780 13921 23783
rect 13596 23752 13921 23780
rect 13596 23740 13602 23752
rect 13909 23749 13921 23752
rect 13955 23749 13967 23783
rect 13909 23743 13967 23749
rect 15381 23783 15439 23789
rect 15381 23749 15393 23783
rect 15427 23780 15439 23783
rect 15470 23780 15476 23792
rect 15427 23752 15476 23780
rect 15427 23749 15439 23752
rect 15381 23743 15439 23749
rect 15470 23740 15476 23752
rect 15528 23740 15534 23792
rect 16301 23783 16359 23789
rect 16301 23749 16313 23783
rect 16347 23780 16359 23783
rect 16390 23780 16396 23792
rect 16347 23752 16396 23780
rect 16347 23749 16359 23752
rect 16301 23743 16359 23749
rect 16390 23740 16396 23752
rect 16448 23740 16454 23792
rect 17310 23780 17316 23792
rect 17271 23752 17316 23780
rect 17310 23740 17316 23752
rect 17368 23740 17374 23792
rect 17405 23783 17463 23789
rect 17405 23749 17417 23783
rect 17451 23780 17463 23783
rect 18046 23780 18052 23792
rect 17451 23752 18052 23780
rect 17451 23749 17463 23752
rect 17405 23743 17463 23749
rect 18046 23740 18052 23752
rect 18104 23740 18110 23792
rect 18969 23783 19027 23789
rect 18969 23749 18981 23783
rect 19015 23780 19027 23783
rect 19705 23783 19763 23789
rect 19705 23780 19717 23783
rect 19015 23752 19717 23780
rect 19015 23749 19027 23752
rect 18969 23743 19027 23749
rect 19705 23749 19717 23752
rect 19751 23749 19763 23783
rect 19705 23743 19763 23749
rect 20346 23740 20352 23792
rect 20404 23780 20410 23792
rect 21177 23783 21235 23789
rect 21177 23780 21189 23783
rect 20404 23752 21189 23780
rect 20404 23740 20410 23752
rect 21177 23749 21189 23752
rect 21223 23749 21235 23783
rect 21177 23743 21235 23749
rect 10321 23715 10379 23721
rect 10321 23681 10333 23715
rect 10367 23681 10379 23715
rect 10321 23675 10379 23681
rect 10870 23672 10876 23724
rect 10928 23712 10934 23724
rect 10965 23715 11023 23721
rect 10965 23712 10977 23715
rect 10928 23684 10977 23712
rect 10928 23672 10934 23684
rect 10965 23681 10977 23684
rect 11011 23681 11023 23715
rect 10965 23675 11023 23681
rect 11054 23672 11060 23724
rect 11112 23712 11118 23724
rect 11885 23715 11943 23721
rect 11885 23712 11897 23715
rect 11112 23684 11897 23712
rect 11112 23672 11118 23684
rect 11885 23681 11897 23684
rect 11931 23712 11943 23715
rect 11974 23712 11980 23724
rect 11931 23684 11980 23712
rect 11931 23681 11943 23684
rect 11885 23675 11943 23681
rect 11974 23672 11980 23684
rect 12032 23672 12038 23724
rect 19797 23715 19855 23721
rect 19797 23681 19809 23715
rect 19843 23712 19855 23715
rect 20622 23712 20628 23724
rect 19843 23684 20628 23712
rect 19843 23681 19855 23684
rect 19797 23675 19855 23681
rect 20622 23672 20628 23684
rect 20680 23672 20686 23724
rect 26329 23715 26387 23721
rect 26329 23681 26341 23715
rect 26375 23712 26387 23715
rect 27264 23712 27292 23808
rect 26375 23684 27292 23712
rect 30101 23715 30159 23721
rect 26375 23681 26387 23684
rect 26329 23675 26387 23681
rect 30101 23681 30113 23715
rect 30147 23712 30159 23715
rect 30653 23715 30711 23721
rect 30653 23712 30665 23715
rect 30147 23684 30665 23712
rect 30147 23681 30159 23684
rect 30101 23675 30159 23681
rect 30653 23681 30665 23684
rect 30699 23712 30711 23715
rect 37826 23712 37832 23724
rect 30699 23684 37832 23712
rect 30699 23681 30711 23684
rect 30653 23675 30711 23681
rect 37826 23672 37832 23684
rect 37884 23672 37890 23724
rect 38010 23712 38016 23724
rect 37971 23684 38016 23712
rect 38010 23672 38016 23684
rect 38068 23672 38074 23724
rect 5074 23604 5080 23656
rect 5132 23644 5138 23656
rect 7193 23647 7251 23653
rect 7193 23644 7205 23647
rect 5132 23616 7205 23644
rect 5132 23604 5138 23616
rect 7193 23613 7205 23616
rect 7239 23644 7251 23647
rect 8386 23644 8392 23656
rect 7239 23616 8392 23644
rect 7239 23613 7251 23616
rect 7193 23607 7251 23613
rect 8386 23604 8392 23616
rect 8444 23604 8450 23656
rect 8573 23647 8631 23653
rect 8573 23613 8585 23647
rect 8619 23644 8631 23647
rect 9398 23644 9404 23656
rect 8619 23616 9404 23644
rect 8619 23613 8631 23616
rect 8573 23607 8631 23613
rect 9398 23604 9404 23616
rect 9456 23604 9462 23656
rect 9769 23647 9827 23653
rect 9769 23613 9781 23647
rect 9815 23644 9827 23647
rect 12250 23644 12256 23656
rect 9815 23616 12256 23644
rect 9815 23613 9827 23616
rect 9769 23607 9827 23613
rect 12250 23604 12256 23616
rect 12308 23604 12314 23656
rect 12434 23604 12440 23656
rect 12492 23644 12498 23656
rect 12621 23647 12679 23653
rect 12621 23644 12633 23647
rect 12492 23616 12633 23644
rect 12492 23604 12498 23616
rect 12621 23613 12633 23616
rect 12667 23644 12679 23647
rect 13814 23644 13820 23656
rect 12667 23616 13820 23644
rect 12667 23613 12679 23616
rect 12621 23607 12679 23613
rect 13814 23604 13820 23616
rect 13872 23604 13878 23656
rect 15010 23604 15016 23656
rect 15068 23644 15074 23656
rect 15289 23647 15347 23653
rect 15289 23644 15301 23647
rect 15068 23616 15301 23644
rect 15068 23604 15074 23616
rect 15289 23613 15301 23616
rect 15335 23613 15347 23647
rect 15289 23607 15347 23613
rect 16482 23604 16488 23656
rect 16540 23644 16546 23656
rect 19061 23647 19119 23653
rect 19061 23644 19073 23647
rect 16540 23616 19073 23644
rect 16540 23604 16546 23616
rect 19061 23613 19073 23616
rect 19107 23613 19119 23647
rect 19061 23607 19119 23613
rect 5810 23536 5816 23588
rect 5868 23576 5874 23588
rect 6733 23579 6791 23585
rect 6733 23576 6745 23579
rect 5868 23548 6745 23576
rect 5868 23536 5874 23548
rect 6733 23545 6745 23548
rect 6779 23576 6791 23579
rect 10870 23576 10876 23588
rect 6779 23548 10876 23576
rect 6779 23545 6791 23548
rect 6733 23539 6791 23545
rect 10870 23536 10876 23548
rect 10928 23576 10934 23588
rect 11882 23576 11888 23588
rect 10928 23548 11888 23576
rect 10928 23536 10934 23548
rect 11882 23536 11888 23548
rect 11940 23536 11946 23588
rect 14366 23576 14372 23588
rect 14327 23548 14372 23576
rect 14366 23536 14372 23548
rect 14424 23536 14430 23588
rect 17034 23536 17040 23588
rect 17092 23576 17098 23588
rect 17494 23576 17500 23588
rect 17092 23548 17500 23576
rect 17092 23536 17098 23548
rect 17494 23536 17500 23548
rect 17552 23576 17558 23588
rect 17865 23579 17923 23585
rect 17865 23576 17877 23579
rect 17552 23548 17877 23576
rect 17552 23536 17558 23548
rect 17865 23545 17877 23548
rect 17911 23576 17923 23579
rect 18509 23579 18567 23585
rect 18509 23576 18521 23579
rect 17911 23548 18521 23576
rect 17911 23545 17923 23548
rect 17865 23539 17923 23545
rect 18509 23545 18521 23548
rect 18555 23545 18567 23579
rect 21266 23576 21272 23588
rect 18509 23539 18567 23545
rect 19306 23548 21272 23576
rect 1765 23511 1823 23517
rect 1765 23477 1777 23511
rect 1811 23508 1823 23511
rect 1854 23508 1860 23520
rect 1811 23480 1860 23508
rect 1811 23477 1823 23480
rect 1765 23471 1823 23477
rect 1854 23468 1860 23480
rect 1912 23468 1918 23520
rect 4614 23508 4620 23520
rect 4575 23480 4620 23508
rect 4614 23468 4620 23480
rect 4672 23468 4678 23520
rect 9125 23511 9183 23517
rect 9125 23477 9137 23511
rect 9171 23508 9183 23511
rect 11606 23508 11612 23520
rect 9171 23480 11612 23508
rect 9171 23477 9183 23480
rect 9125 23471 9183 23477
rect 11606 23468 11612 23480
rect 11664 23468 11670 23520
rect 11974 23508 11980 23520
rect 11935 23480 11980 23508
rect 11974 23468 11980 23480
rect 12032 23468 12038 23520
rect 12618 23468 12624 23520
rect 12676 23508 12682 23520
rect 15746 23508 15752 23520
rect 12676 23480 15752 23508
rect 12676 23468 12682 23480
rect 15746 23468 15752 23480
rect 15804 23468 15810 23520
rect 17126 23468 17132 23520
rect 17184 23508 17190 23520
rect 19306 23508 19334 23548
rect 21266 23536 21272 23548
rect 21324 23536 21330 23588
rect 20714 23508 20720 23520
rect 17184 23480 19334 23508
rect 20675 23480 20720 23508
rect 17184 23468 17190 23480
rect 20714 23468 20720 23480
rect 20772 23468 20778 23520
rect 38194 23508 38200 23520
rect 38155 23480 38200 23508
rect 38194 23468 38200 23480
rect 38252 23468 38258 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 1670 23304 1676 23316
rect 1631 23276 1676 23304
rect 1670 23264 1676 23276
rect 1728 23304 1734 23316
rect 2406 23304 2412 23316
rect 1728 23276 2412 23304
rect 1728 23264 1734 23276
rect 2406 23264 2412 23276
rect 2464 23304 2470 23316
rect 2685 23307 2743 23313
rect 2685 23304 2697 23307
rect 2464 23276 2697 23304
rect 2464 23264 2470 23276
rect 2685 23273 2697 23276
rect 2731 23273 2743 23307
rect 3234 23304 3240 23316
rect 3195 23276 3240 23304
rect 2685 23267 2743 23273
rect 2700 23236 2728 23267
rect 3234 23264 3240 23276
rect 3292 23264 3298 23316
rect 7009 23307 7067 23313
rect 7009 23273 7021 23307
rect 7055 23304 7067 23307
rect 8294 23304 8300 23316
rect 7055 23276 8300 23304
rect 7055 23273 7067 23276
rect 7009 23267 7067 23273
rect 8294 23264 8300 23276
rect 8352 23264 8358 23316
rect 8478 23304 8484 23316
rect 8439 23276 8484 23304
rect 8478 23264 8484 23276
rect 8536 23264 8542 23316
rect 11238 23304 11244 23316
rect 9968 23276 11244 23304
rect 9968 23245 9996 23276
rect 11238 23264 11244 23276
rect 11296 23264 11302 23316
rect 13633 23307 13691 23313
rect 13633 23273 13645 23307
rect 13679 23304 13691 23307
rect 14734 23304 14740 23316
rect 13679 23276 14740 23304
rect 13679 23273 13691 23276
rect 13633 23267 13691 23273
rect 14734 23264 14740 23276
rect 14792 23264 14798 23316
rect 15286 23264 15292 23316
rect 15344 23304 15350 23316
rect 16209 23307 16267 23313
rect 16209 23304 16221 23307
rect 15344 23276 16221 23304
rect 15344 23264 15350 23276
rect 16209 23273 16221 23276
rect 16255 23273 16267 23307
rect 16209 23267 16267 23273
rect 16850 23264 16856 23316
rect 16908 23304 16914 23316
rect 17770 23304 17776 23316
rect 16908 23276 17776 23304
rect 16908 23264 16914 23276
rect 17770 23264 17776 23276
rect 17828 23264 17834 23316
rect 18046 23304 18052 23316
rect 18007 23276 18052 23304
rect 18046 23264 18052 23276
rect 18104 23264 18110 23316
rect 19150 23264 19156 23316
rect 19208 23304 19214 23316
rect 19978 23304 19984 23316
rect 19208 23276 19984 23304
rect 19208 23264 19214 23276
rect 19978 23264 19984 23276
rect 20036 23264 20042 23316
rect 9953 23239 10011 23245
rect 2700 23208 4384 23236
rect 2225 23035 2283 23041
rect 2225 23001 2237 23035
rect 2271 23032 2283 23035
rect 3786 23032 3792 23044
rect 2271 23004 3792 23032
rect 2271 23001 2283 23004
rect 2225 22995 2283 23001
rect 3786 22992 3792 23004
rect 3844 22992 3850 23044
rect 4356 23041 4384 23208
rect 9953 23205 9965 23239
rect 9999 23205 10011 23239
rect 9953 23199 10011 23205
rect 10870 23196 10876 23248
rect 10928 23236 10934 23248
rect 12802 23236 12808 23248
rect 10928 23208 12808 23236
rect 10928 23196 10934 23208
rect 12802 23196 12808 23208
rect 12860 23196 12866 23248
rect 12989 23239 13047 23245
rect 12989 23205 13001 23239
rect 13035 23236 13047 23239
rect 13035 23208 14504 23236
rect 13035 23205 13047 23208
rect 12989 23199 13047 23205
rect 8846 23168 8852 23180
rect 7668 23140 8852 23168
rect 7668 23109 7696 23140
rect 8846 23128 8852 23140
rect 8904 23128 8910 23180
rect 9398 23168 9404 23180
rect 9359 23140 9404 23168
rect 9398 23128 9404 23140
rect 9456 23128 9462 23180
rect 10042 23128 10048 23180
rect 10100 23168 10106 23180
rect 10597 23171 10655 23177
rect 10597 23168 10609 23171
rect 10100 23140 10609 23168
rect 10100 23128 10106 23140
rect 10597 23137 10609 23140
rect 10643 23137 10655 23171
rect 10597 23131 10655 23137
rect 11241 23171 11299 23177
rect 11241 23137 11253 23171
rect 11287 23168 11299 23171
rect 11514 23168 11520 23180
rect 11287 23140 11520 23168
rect 11287 23137 11299 23140
rect 11241 23131 11299 23137
rect 11514 23128 11520 23140
rect 11572 23168 11578 23180
rect 11882 23168 11888 23180
rect 11572 23140 11888 23168
rect 11572 23128 11578 23140
rect 11882 23128 11888 23140
rect 11940 23128 11946 23180
rect 13814 23128 13820 23180
rect 13872 23168 13878 23180
rect 14369 23171 14427 23177
rect 14369 23168 14381 23171
rect 13872 23140 14381 23168
rect 13872 23128 13878 23140
rect 14369 23137 14381 23140
rect 14415 23137 14427 23171
rect 14476 23168 14504 23208
rect 14550 23196 14556 23248
rect 14608 23236 14614 23248
rect 15565 23239 15623 23245
rect 15565 23236 15577 23239
rect 14608 23208 15577 23236
rect 14608 23196 14614 23208
rect 15565 23205 15577 23208
rect 15611 23205 15623 23239
rect 15565 23199 15623 23205
rect 17862 23196 17868 23248
rect 17920 23236 17926 23248
rect 18693 23239 18751 23245
rect 18693 23236 18705 23239
rect 17920 23208 18705 23236
rect 17920 23196 17926 23208
rect 18693 23205 18705 23208
rect 18739 23205 18751 23239
rect 18693 23199 18751 23205
rect 16022 23168 16028 23180
rect 14476 23140 16028 23168
rect 14369 23131 14427 23137
rect 16022 23128 16028 23140
rect 16080 23128 16086 23180
rect 17129 23171 17187 23177
rect 17129 23168 17141 23171
rect 16132 23140 17141 23168
rect 7653 23103 7711 23109
rect 7653 23069 7665 23103
rect 7699 23069 7711 23103
rect 7653 23063 7711 23069
rect 8389 23103 8447 23109
rect 8389 23069 8401 23103
rect 8435 23069 8447 23103
rect 13446 23100 13452 23112
rect 13407 23072 13452 23100
rect 8389 23063 8447 23069
rect 4341 23035 4399 23041
rect 4341 23001 4353 23035
rect 4387 23032 4399 23035
rect 6089 23035 6147 23041
rect 6089 23032 6101 23035
rect 4387 23004 6101 23032
rect 4387 23001 4399 23004
rect 4341 22995 4399 23001
rect 6089 23001 6101 23004
rect 6135 23001 6147 23035
rect 6089 22995 6147 23001
rect 6362 22992 6368 23044
rect 6420 23032 6426 23044
rect 8404 23032 8432 23063
rect 13446 23060 13452 23072
rect 13504 23060 13510 23112
rect 15562 23060 15568 23112
rect 15620 23100 15626 23112
rect 15657 23103 15715 23109
rect 15657 23100 15669 23103
rect 15620 23072 15669 23100
rect 15620 23060 15626 23072
rect 15657 23069 15669 23072
rect 15703 23069 15715 23103
rect 16132 23100 16160 23140
rect 17129 23137 17141 23140
rect 17175 23168 17187 23171
rect 17218 23168 17224 23180
rect 17175 23140 17224 23168
rect 17175 23137 17187 23140
rect 17129 23131 17187 23137
rect 17218 23128 17224 23140
rect 17276 23128 17282 23180
rect 21545 23171 21603 23177
rect 21545 23168 21557 23171
rect 18248 23140 21557 23168
rect 18248 23112 18276 23140
rect 21545 23137 21557 23140
rect 21591 23137 21603 23171
rect 31754 23168 31760 23180
rect 21545 23131 21603 23137
rect 22066 23140 31760 23168
rect 15657 23063 15715 23069
rect 15764 23072 16160 23100
rect 16301 23103 16359 23109
rect 6420 23004 8432 23032
rect 6420 22992 6426 23004
rect 8662 22992 8668 23044
rect 8720 23032 8726 23044
rect 9493 23035 9551 23041
rect 9493 23032 9505 23035
rect 8720 23004 9505 23032
rect 8720 22992 8726 23004
rect 9493 23001 9505 23004
rect 9539 23001 9551 23035
rect 9493 22995 9551 23001
rect 10689 23035 10747 23041
rect 10689 23001 10701 23035
rect 10735 23001 10747 23035
rect 11790 23032 11796 23044
rect 11751 23004 11796 23032
rect 10689 22995 10747 23001
rect 3418 22924 3424 22976
rect 3476 22964 3482 22976
rect 4614 22964 4620 22976
rect 3476 22936 4620 22964
rect 3476 22924 3482 22936
rect 4614 22924 4620 22936
rect 4672 22964 4678 22976
rect 4893 22967 4951 22973
rect 4893 22964 4905 22967
rect 4672 22936 4905 22964
rect 4672 22924 4678 22936
rect 4893 22933 4905 22936
rect 4939 22933 4951 22967
rect 5534 22964 5540 22976
rect 5495 22936 5540 22964
rect 4893 22927 4951 22933
rect 5534 22924 5540 22936
rect 5592 22924 5598 22976
rect 7558 22964 7564 22976
rect 7519 22936 7564 22964
rect 7558 22924 7564 22936
rect 7616 22924 7622 22976
rect 9858 22924 9864 22976
rect 9916 22964 9922 22976
rect 10704 22964 10732 22995
rect 11790 22992 11796 23004
rect 11848 22992 11854 23044
rect 11885 23035 11943 23041
rect 11885 23001 11897 23035
rect 11931 23001 11943 23035
rect 11885 22995 11943 23001
rect 12437 23035 12495 23041
rect 12437 23001 12449 23035
rect 12483 23032 12495 23035
rect 13906 23032 13912 23044
rect 12483 23004 13912 23032
rect 12483 23001 12495 23004
rect 12437 22995 12495 23001
rect 9916 22936 10732 22964
rect 9916 22924 9922 22936
rect 10778 22924 10784 22976
rect 10836 22964 10842 22976
rect 11900 22964 11928 22995
rect 13906 22992 13912 23004
rect 13964 22992 13970 23044
rect 14461 23035 14519 23041
rect 14461 23001 14473 23035
rect 14507 23001 14519 23035
rect 15010 23032 15016 23044
rect 14971 23004 15016 23032
rect 14461 22995 14519 23001
rect 10836 22936 11928 22964
rect 10836 22924 10842 22936
rect 12618 22924 12624 22976
rect 12676 22964 12682 22976
rect 14469 22964 14497 22995
rect 15010 22992 15016 23004
rect 15068 22992 15074 23044
rect 12676 22936 14497 22964
rect 12676 22924 12682 22936
rect 14550 22924 14556 22976
rect 14608 22964 14614 22976
rect 15764 22964 15792 23072
rect 16301 23069 16313 23103
rect 16347 23100 16359 23103
rect 16758 23100 16764 23112
rect 16347 23072 16764 23100
rect 16347 23069 16359 23072
rect 16301 23063 16359 23069
rect 16758 23060 16764 23072
rect 16816 23060 16822 23112
rect 17770 23060 17776 23112
rect 17828 23100 17834 23112
rect 18141 23103 18199 23109
rect 18141 23100 18153 23103
rect 17828 23072 18153 23100
rect 17828 23060 17834 23072
rect 18141 23069 18153 23072
rect 18187 23100 18199 23103
rect 18230 23100 18236 23112
rect 18187 23072 18236 23100
rect 18187 23069 18199 23072
rect 18141 23063 18199 23069
rect 18230 23060 18236 23072
rect 18288 23060 18294 23112
rect 18785 23103 18843 23109
rect 18785 23069 18797 23103
rect 18831 23100 18843 23103
rect 18966 23100 18972 23112
rect 18831 23072 18972 23100
rect 18831 23069 18843 23072
rect 18785 23063 18843 23069
rect 18966 23060 18972 23072
rect 19024 23060 19030 23112
rect 19334 23060 19340 23112
rect 19392 23100 19398 23112
rect 19613 23103 19671 23109
rect 19613 23100 19625 23103
rect 19392 23072 19625 23100
rect 19392 23060 19398 23072
rect 19613 23069 19625 23072
rect 19659 23069 19671 23103
rect 19613 23063 19671 23069
rect 20714 23060 20720 23112
rect 20772 23100 20778 23112
rect 20898 23100 20904 23112
rect 20772 23072 20904 23100
rect 20772 23060 20778 23072
rect 20898 23060 20904 23072
rect 20956 23060 20962 23112
rect 16114 22992 16120 23044
rect 16172 23032 16178 23044
rect 17313 23035 17371 23041
rect 16172 23004 16344 23032
rect 16172 22992 16178 23004
rect 14608 22936 15792 22964
rect 16316 22964 16344 23004
rect 17313 23001 17325 23035
rect 17359 23001 17371 23035
rect 17313 22995 17371 23001
rect 17405 23035 17463 23041
rect 17405 23001 17417 23035
rect 17451 23001 17463 23035
rect 17405 22995 17463 23001
rect 17328 22964 17356 22995
rect 16316 22936 17356 22964
rect 17420 22964 17448 22995
rect 17678 22992 17684 23044
rect 17736 23032 17742 23044
rect 19521 23035 19579 23041
rect 19521 23032 19533 23035
rect 17736 23004 19533 23032
rect 17736 22992 17742 23004
rect 19521 23001 19533 23004
rect 19567 23001 19579 23035
rect 19521 22995 19579 23001
rect 21085 23035 21143 23041
rect 21085 23001 21097 23035
rect 21131 23032 21143 23035
rect 22066 23032 22094 23140
rect 31754 23128 31760 23140
rect 31812 23128 31818 23180
rect 22922 23060 22928 23112
rect 22980 23100 22986 23112
rect 29917 23103 29975 23109
rect 29917 23100 29929 23103
rect 22980 23072 29929 23100
rect 22980 23060 22986 23072
rect 29917 23069 29929 23072
rect 29963 23100 29975 23103
rect 30561 23103 30619 23109
rect 30561 23100 30573 23103
rect 29963 23072 30573 23100
rect 29963 23069 29975 23072
rect 29917 23063 29975 23069
rect 30561 23069 30573 23072
rect 30607 23069 30619 23103
rect 30561 23063 30619 23069
rect 21131 23004 22094 23032
rect 30116 23004 35894 23032
rect 21131 23001 21143 23004
rect 21085 22995 21143 23001
rect 18414 22964 18420 22976
rect 17420 22936 18420 22964
rect 14608 22924 14614 22936
rect 18414 22924 18420 22936
rect 18472 22964 18478 22976
rect 18598 22964 18604 22976
rect 18472 22936 18604 22964
rect 18472 22924 18478 22936
rect 18598 22924 18604 22936
rect 18656 22924 18662 22976
rect 20070 22964 20076 22976
rect 20031 22936 20076 22964
rect 20070 22924 20076 22936
rect 20128 22924 20134 22976
rect 30116 22973 30144 23004
rect 30101 22967 30159 22973
rect 30101 22933 30113 22967
rect 30147 22933 30159 22967
rect 35866 22964 35894 23004
rect 38010 22964 38016 22976
rect 35866 22936 38016 22964
rect 30101 22927 30159 22933
rect 38010 22924 38016 22936
rect 38068 22924 38074 22976
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 2317 22763 2375 22769
rect 2317 22729 2329 22763
rect 2363 22729 2375 22763
rect 3786 22760 3792 22772
rect 3747 22732 3792 22760
rect 2317 22723 2375 22729
rect 1857 22627 1915 22633
rect 1857 22593 1869 22627
rect 1903 22624 1915 22627
rect 2332 22624 2360 22723
rect 3786 22720 3792 22732
rect 3844 22760 3850 22772
rect 4062 22760 4068 22772
rect 3844 22732 4068 22760
rect 3844 22720 3850 22732
rect 4062 22720 4068 22732
rect 4120 22720 4126 22772
rect 5442 22760 5448 22772
rect 5403 22732 5448 22760
rect 5442 22720 5448 22732
rect 5500 22720 5506 22772
rect 8662 22760 8668 22772
rect 8623 22732 8668 22760
rect 8662 22720 8668 22732
rect 8720 22720 8726 22772
rect 9953 22763 10011 22769
rect 9953 22729 9965 22763
rect 9999 22760 10011 22763
rect 12526 22760 12532 22772
rect 9999 22732 12532 22760
rect 9999 22729 10011 22732
rect 9953 22723 10011 22729
rect 12526 22720 12532 22732
rect 12584 22720 12590 22772
rect 12710 22720 12716 22772
rect 12768 22760 12774 22772
rect 13081 22763 13139 22769
rect 13081 22760 13093 22763
rect 12768 22732 13093 22760
rect 12768 22720 12774 22732
rect 13081 22729 13093 22732
rect 13127 22729 13139 22763
rect 13081 22723 13139 22729
rect 13262 22720 13268 22772
rect 13320 22760 13326 22772
rect 13446 22760 13452 22772
rect 13320 22732 13452 22760
rect 13320 22720 13326 22732
rect 13446 22720 13452 22732
rect 13504 22720 13510 22772
rect 15194 22760 15200 22772
rect 14200 22732 15200 22760
rect 4893 22695 4951 22701
rect 4893 22661 4905 22695
rect 4939 22692 4951 22695
rect 5994 22692 6000 22704
rect 4939 22664 6000 22692
rect 4939 22661 4951 22664
rect 4893 22655 4951 22661
rect 5994 22652 6000 22664
rect 6052 22652 6058 22704
rect 7561 22695 7619 22701
rect 7561 22661 7573 22695
rect 7607 22692 7619 22695
rect 7607 22664 9444 22692
rect 7607 22661 7619 22664
rect 7561 22655 7619 22661
rect 9416 22636 9444 22664
rect 11606 22652 11612 22704
rect 11664 22692 11670 22704
rect 11885 22695 11943 22701
rect 11885 22692 11897 22695
rect 11664 22664 11897 22692
rect 11664 22652 11670 22664
rect 11885 22661 11897 22664
rect 11931 22661 11943 22695
rect 11885 22655 11943 22661
rect 12158 22652 12164 22704
rect 12216 22692 12222 22704
rect 14200 22701 14228 22732
rect 15194 22720 15200 22732
rect 15252 22720 15258 22772
rect 18046 22760 18052 22772
rect 18007 22732 18052 22760
rect 18046 22720 18052 22732
rect 18104 22720 18110 22772
rect 22186 22760 22192 22772
rect 19536 22732 22192 22760
rect 14185 22695 14243 22701
rect 12216 22664 13124 22692
rect 12216 22652 12222 22664
rect 1903 22596 2360 22624
rect 2501 22627 2559 22633
rect 1903 22593 1915 22596
rect 1857 22587 1915 22593
rect 2501 22593 2513 22627
rect 2547 22624 2559 22627
rect 8570 22624 8576 22636
rect 2547 22596 2581 22624
rect 8531 22596 8576 22624
rect 2547 22593 2559 22596
rect 2501 22587 2559 22593
rect 1946 22516 1952 22568
rect 2004 22556 2010 22568
rect 2516 22556 2544 22587
rect 8570 22584 8576 22596
rect 8628 22584 8634 22636
rect 9398 22624 9404 22636
rect 9311 22596 9404 22624
rect 9398 22584 9404 22596
rect 9456 22584 9462 22636
rect 9861 22627 9919 22633
rect 9861 22624 9873 22627
rect 9600 22596 9873 22624
rect 2961 22559 3019 22565
rect 2961 22556 2973 22559
rect 2004 22528 2973 22556
rect 2004 22516 2010 22528
rect 2961 22525 2973 22528
rect 3007 22525 3019 22559
rect 2961 22519 3019 22525
rect 8113 22559 8171 22565
rect 8113 22525 8125 22559
rect 8159 22556 8171 22559
rect 9600 22556 9628 22596
rect 9861 22593 9873 22596
rect 9907 22624 9919 22627
rect 10870 22624 10876 22636
rect 9907 22596 10876 22624
rect 9907 22593 9919 22596
rect 9861 22587 9919 22593
rect 10870 22584 10876 22596
rect 10928 22584 10934 22636
rect 12989 22627 13047 22633
rect 12989 22593 13001 22627
rect 13035 22593 13047 22627
rect 12989 22587 13047 22593
rect 8159 22528 9628 22556
rect 8159 22525 8171 22528
rect 8113 22519 8171 22525
rect 9674 22516 9680 22568
rect 9732 22556 9738 22568
rect 10505 22559 10563 22565
rect 10505 22556 10517 22559
rect 9732 22528 10517 22556
rect 9732 22516 9738 22528
rect 10505 22525 10517 22528
rect 10551 22525 10563 22559
rect 10686 22556 10692 22568
rect 10647 22528 10692 22556
rect 10505 22519 10563 22525
rect 1670 22488 1676 22500
rect 1631 22460 1676 22488
rect 1670 22448 1676 22460
rect 1728 22448 1734 22500
rect 2038 22448 2044 22500
rect 2096 22488 2102 22500
rect 9217 22491 9275 22497
rect 9217 22488 9229 22491
rect 2096 22460 9229 22488
rect 2096 22448 2102 22460
rect 9217 22457 9229 22460
rect 9263 22457 9275 22491
rect 10520 22488 10548 22519
rect 10686 22516 10692 22528
rect 10744 22516 10750 22568
rect 11793 22559 11851 22565
rect 11793 22525 11805 22559
rect 11839 22525 11851 22559
rect 11793 22519 11851 22525
rect 11808 22488 11836 22519
rect 11882 22516 11888 22568
rect 11940 22556 11946 22568
rect 12069 22559 12127 22565
rect 12069 22556 12081 22559
rect 11940 22528 12081 22556
rect 11940 22516 11946 22528
rect 12069 22525 12081 22528
rect 12115 22525 12127 22559
rect 12069 22519 12127 22525
rect 10520 22460 12112 22488
rect 9217 22451 9275 22457
rect 5534 22380 5540 22432
rect 5592 22420 5598 22432
rect 5997 22423 6055 22429
rect 5997 22420 6009 22423
rect 5592 22392 6009 22420
rect 5592 22380 5598 22392
rect 5997 22389 6009 22392
rect 6043 22420 6055 22423
rect 6454 22420 6460 22432
rect 6043 22392 6460 22420
rect 6043 22389 6055 22392
rect 5997 22383 6055 22389
rect 6454 22380 6460 22392
rect 6512 22420 6518 22432
rect 6825 22423 6883 22429
rect 6825 22420 6837 22423
rect 6512 22392 6837 22420
rect 6512 22380 6518 22392
rect 6825 22389 6837 22392
rect 6871 22389 6883 22423
rect 11054 22420 11060 22432
rect 11015 22392 11060 22420
rect 6825 22383 6883 22389
rect 11054 22380 11060 22392
rect 11112 22380 11118 22432
rect 12084 22420 12112 22460
rect 12250 22448 12256 22500
rect 12308 22488 12314 22500
rect 13004 22488 13032 22587
rect 13096 22556 13124 22664
rect 14185 22661 14197 22695
rect 14231 22661 14243 22695
rect 14918 22692 14924 22704
rect 14879 22664 14924 22692
rect 14185 22655 14243 22661
rect 14918 22652 14924 22664
rect 14976 22652 14982 22704
rect 15013 22695 15071 22701
rect 15013 22661 15025 22695
rect 15059 22692 15071 22695
rect 16117 22695 16175 22701
rect 16117 22692 16129 22695
rect 15059 22664 16129 22692
rect 15059 22661 15071 22664
rect 15013 22655 15071 22661
rect 16117 22661 16129 22664
rect 16163 22661 16175 22695
rect 16117 22655 16175 22661
rect 16298 22652 16304 22704
rect 16356 22692 16362 22704
rect 19536 22701 19564 22732
rect 22186 22720 22192 22732
rect 22244 22720 22250 22772
rect 18969 22695 19027 22701
rect 18969 22692 18981 22695
rect 16356 22664 18981 22692
rect 16356 22652 16362 22664
rect 18969 22661 18981 22664
rect 19015 22661 19027 22695
rect 18969 22655 19027 22661
rect 19521 22695 19579 22701
rect 19521 22661 19533 22695
rect 19567 22661 19579 22695
rect 20162 22692 20168 22704
rect 20123 22664 20168 22692
rect 19521 22655 19579 22661
rect 20162 22652 20168 22664
rect 20220 22652 20226 22704
rect 20717 22695 20775 22701
rect 20717 22661 20729 22695
rect 20763 22692 20775 22695
rect 20806 22692 20812 22704
rect 20763 22664 20812 22692
rect 20763 22661 20775 22664
rect 20717 22655 20775 22661
rect 16022 22584 16028 22636
rect 16080 22624 16086 22636
rect 16209 22627 16267 22633
rect 16209 22624 16221 22627
rect 16080 22596 16221 22624
rect 16080 22584 16086 22596
rect 16209 22593 16221 22596
rect 16255 22593 16267 22627
rect 17586 22624 17592 22636
rect 17547 22596 17592 22624
rect 16209 22587 16267 22593
rect 17586 22584 17592 22596
rect 17644 22584 17650 22636
rect 18233 22627 18291 22633
rect 18233 22593 18245 22627
rect 18279 22593 18291 22627
rect 18233 22587 18291 22593
rect 14001 22559 14059 22565
rect 14001 22556 14013 22559
rect 13096 22528 14013 22556
rect 14001 22525 14013 22528
rect 14047 22525 14059 22559
rect 14001 22519 14059 22525
rect 14277 22559 14335 22565
rect 14277 22525 14289 22559
rect 14323 22556 14335 22559
rect 15378 22556 15384 22568
rect 14323 22528 15384 22556
rect 14323 22525 14335 22528
rect 14277 22519 14335 22525
rect 12308 22460 13032 22488
rect 14016 22488 14044 22519
rect 15378 22516 15384 22528
rect 15436 22516 15442 22568
rect 16850 22516 16856 22568
rect 16908 22556 16914 22568
rect 16945 22559 17003 22565
rect 16945 22556 16957 22559
rect 16908 22528 16957 22556
rect 16908 22516 16914 22528
rect 16945 22525 16957 22528
rect 16991 22556 17003 22559
rect 18248 22556 18276 22587
rect 16991 22528 18276 22556
rect 16991 22525 17003 22528
rect 16945 22519 17003 22525
rect 18322 22516 18328 22568
rect 18380 22556 18386 22568
rect 18877 22559 18935 22565
rect 18877 22556 18889 22559
rect 18380 22528 18889 22556
rect 18380 22516 18386 22528
rect 18877 22525 18889 22528
rect 18923 22525 18935 22559
rect 20070 22556 20076 22568
rect 20031 22528 20076 22556
rect 18877 22519 18935 22525
rect 20070 22516 20076 22528
rect 20128 22516 20134 22568
rect 20346 22516 20352 22568
rect 20404 22556 20410 22568
rect 20732 22556 20760 22655
rect 20806 22652 20812 22664
rect 20864 22652 20870 22704
rect 20404 22528 20760 22556
rect 20404 22516 20410 22528
rect 14550 22488 14556 22500
rect 14016 22460 14556 22488
rect 12308 22448 12314 22460
rect 14550 22448 14556 22460
rect 14608 22448 14614 22500
rect 15473 22491 15531 22497
rect 15473 22457 15485 22491
rect 15519 22488 15531 22491
rect 15519 22460 19380 22488
rect 15519 22457 15531 22460
rect 15473 22451 15531 22457
rect 12894 22420 12900 22432
rect 12084 22392 12900 22420
rect 12894 22380 12900 22392
rect 12952 22380 12958 22432
rect 15286 22380 15292 22432
rect 15344 22420 15350 22432
rect 17497 22423 17555 22429
rect 17497 22420 17509 22423
rect 15344 22392 17509 22420
rect 15344 22380 15350 22392
rect 17497 22389 17509 22392
rect 17543 22389 17555 22423
rect 19352 22420 19380 22460
rect 23566 22420 23572 22432
rect 19352 22392 23572 22420
rect 17497 22383 17555 22389
rect 23566 22380 23572 22392
rect 23624 22380 23630 22432
rect 37826 22380 37832 22432
rect 37884 22420 37890 22432
rect 38105 22423 38163 22429
rect 38105 22420 38117 22423
rect 37884 22392 38117 22420
rect 37884 22380 37890 22392
rect 38105 22389 38117 22392
rect 38151 22389 38163 22423
rect 38105 22383 38163 22389
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 2406 22216 2412 22228
rect 2367 22188 2412 22216
rect 2406 22176 2412 22188
rect 2464 22176 2470 22228
rect 8481 22219 8539 22225
rect 8481 22185 8493 22219
rect 8527 22216 8539 22219
rect 12434 22216 12440 22228
rect 8527 22188 12440 22216
rect 8527 22185 8539 22188
rect 8481 22179 8539 22185
rect 12434 22176 12440 22188
rect 12492 22176 12498 22228
rect 15562 22176 15568 22228
rect 15620 22216 15626 22228
rect 20438 22216 20444 22228
rect 15620 22188 20444 22216
rect 15620 22176 15626 22188
rect 20438 22176 20444 22188
rect 20496 22176 20502 22228
rect 6454 22148 6460 22160
rect 6415 22120 6460 22148
rect 6454 22108 6460 22120
rect 6512 22108 6518 22160
rect 11238 22108 11244 22160
rect 11296 22148 11302 22160
rect 11609 22151 11667 22157
rect 11609 22148 11621 22151
rect 11296 22120 11621 22148
rect 11296 22108 11302 22120
rect 11609 22117 11621 22120
rect 11655 22117 11667 22151
rect 11609 22111 11667 22117
rect 12345 22151 12403 22157
rect 12345 22117 12357 22151
rect 12391 22148 12403 22151
rect 12618 22148 12624 22160
rect 12391 22120 12624 22148
rect 12391 22117 12403 22120
rect 12345 22111 12403 22117
rect 12618 22108 12624 22120
rect 12676 22108 12682 22160
rect 20456 22148 20484 22176
rect 13464 22120 13768 22148
rect 20456 22120 20576 22148
rect 1673 22083 1731 22089
rect 1673 22049 1685 22083
rect 1719 22080 1731 22083
rect 1762 22080 1768 22092
rect 1719 22052 1768 22080
rect 1719 22049 1731 22052
rect 1673 22043 1731 22049
rect 1762 22040 1768 22052
rect 1820 22040 1826 22092
rect 9217 22083 9275 22089
rect 7300 22052 8432 22080
rect 2958 21972 2964 22024
rect 3016 22012 3022 22024
rect 7300 22021 7328 22052
rect 8404 22021 8432 22052
rect 9217 22049 9229 22083
rect 9263 22080 9275 22083
rect 13464 22080 13492 22120
rect 13630 22080 13636 22092
rect 9263 22052 12296 22080
rect 9263 22049 9275 22052
rect 9217 22043 9275 22049
rect 5445 22015 5503 22021
rect 5445 22012 5457 22015
rect 3016 21984 5457 22012
rect 3016 21972 3022 21984
rect 5445 21981 5457 21984
rect 5491 22012 5503 22015
rect 5905 22015 5963 22021
rect 5905 22012 5917 22015
rect 5491 21984 5917 22012
rect 5491 21981 5503 21984
rect 5445 21975 5503 21981
rect 5905 21981 5917 21984
rect 5951 22012 5963 22015
rect 7285 22015 7343 22021
rect 7285 22012 7297 22015
rect 5951 21984 7297 22012
rect 5951 21981 5963 21984
rect 5905 21975 5963 21981
rect 7285 21981 7297 21984
rect 7331 21981 7343 22015
rect 7285 21975 7343 21981
rect 8389 22015 8447 22021
rect 8389 21981 8401 22015
rect 8435 21981 8447 22015
rect 9766 22012 9772 22024
rect 9727 21984 9772 22012
rect 8389 21975 8447 21981
rect 9766 21972 9772 21984
rect 9824 21972 9830 22024
rect 9861 22015 9919 22021
rect 9861 21981 9873 22015
rect 9907 22012 9919 22015
rect 10134 22012 10140 22024
rect 9907 21984 10140 22012
rect 9907 21981 9919 21984
rect 9861 21975 9919 21981
rect 10134 21972 10140 21984
rect 10192 21972 10198 22024
rect 10318 22012 10324 22024
rect 10244 21984 10324 22012
rect 4798 21904 4804 21956
rect 4856 21944 4862 21956
rect 7837 21947 7895 21953
rect 7837 21944 7849 21947
rect 4856 21916 7849 21944
rect 4856 21904 4862 21916
rect 7837 21913 7849 21916
rect 7883 21944 7895 21947
rect 10244 21944 10272 21984
rect 10318 21972 10324 21984
rect 10376 22012 10382 22024
rect 12268 22021 12296 22052
rect 12728 22052 13492 22080
rect 13591 22052 13636 22080
rect 12253 22015 12311 22021
rect 10376 21984 10469 22012
rect 10376 21972 10382 21984
rect 12253 21981 12265 22015
rect 12299 22012 12311 22015
rect 12728 22012 12756 22052
rect 13630 22040 13636 22052
rect 13688 22040 13694 22092
rect 13740 22080 13768 22120
rect 17865 22083 17923 22089
rect 13740 22052 16574 22080
rect 14550 22012 14556 22024
rect 12299 21984 12756 22012
rect 14511 21984 14556 22012
rect 12299 21981 12311 21984
rect 12253 21975 12311 21981
rect 14550 21972 14556 21984
rect 14608 21972 14614 22024
rect 15378 21972 15384 22024
rect 15436 22012 15442 22024
rect 16206 22012 16212 22024
rect 15436 21984 16212 22012
rect 15436 21972 15442 21984
rect 16206 21972 16212 21984
rect 16264 21972 16270 22024
rect 7883 21916 10272 21944
rect 10413 21947 10471 21953
rect 7883 21913 7895 21916
rect 7837 21907 7895 21913
rect 10413 21913 10425 21947
rect 10459 21944 10471 21947
rect 11057 21947 11115 21953
rect 11057 21944 11069 21947
rect 10459 21916 11069 21944
rect 10459 21913 10471 21916
rect 10413 21907 10471 21913
rect 11057 21913 11069 21916
rect 11103 21913 11115 21947
rect 11057 21907 11115 21913
rect 3421 21879 3479 21885
rect 3421 21845 3433 21879
rect 3467 21876 3479 21879
rect 4062 21876 4068 21888
rect 3467 21848 4068 21876
rect 3467 21845 3479 21848
rect 3421 21839 3479 21845
rect 4062 21836 4068 21848
rect 4120 21876 4126 21888
rect 4617 21879 4675 21885
rect 4617 21876 4629 21879
rect 4120 21848 4629 21876
rect 4120 21836 4126 21848
rect 4617 21845 4629 21848
rect 4663 21845 4675 21879
rect 5258 21876 5264 21888
rect 5219 21848 5264 21876
rect 4617 21839 4675 21845
rect 5258 21836 5264 21848
rect 5316 21836 5322 21888
rect 8202 21836 8208 21888
rect 8260 21876 8266 21888
rect 10962 21876 10968 21888
rect 8260 21848 10968 21876
rect 8260 21836 8266 21848
rect 10962 21836 10968 21848
rect 11020 21836 11026 21888
rect 11072 21876 11100 21907
rect 11146 21904 11152 21956
rect 11204 21944 11210 21956
rect 12986 21944 12992 21956
rect 11204 21916 11249 21944
rect 12947 21916 12992 21944
rect 11204 21904 11210 21916
rect 12986 21904 12992 21916
rect 13044 21904 13050 21956
rect 13081 21947 13139 21953
rect 13081 21913 13093 21947
rect 13127 21913 13139 21947
rect 13081 21907 13139 21913
rect 15105 21947 15163 21953
rect 15105 21913 15117 21947
rect 15151 21913 15163 21947
rect 15105 21907 15163 21913
rect 15197 21947 15255 21953
rect 15197 21913 15209 21947
rect 15243 21944 15255 21947
rect 15396 21944 15424 21972
rect 15930 21944 15936 21956
rect 15243 21916 15424 21944
rect 15891 21916 15936 21944
rect 15243 21913 15255 21916
rect 15197 21907 15255 21913
rect 11790 21876 11796 21888
rect 11072 21848 11796 21876
rect 11790 21836 11796 21848
rect 11848 21836 11854 21888
rect 11974 21836 11980 21888
rect 12032 21876 12038 21888
rect 13096 21876 13124 21907
rect 12032 21848 13124 21876
rect 15120 21876 15148 21907
rect 15930 21904 15936 21916
rect 15988 21904 15994 21956
rect 16546 21944 16574 22052
rect 17865 22049 17877 22083
rect 17911 22080 17923 22083
rect 18322 22080 18328 22092
rect 17911 22052 18328 22080
rect 17911 22049 17923 22052
rect 17865 22043 17923 22049
rect 18322 22040 18328 22052
rect 18380 22040 18386 22092
rect 18509 22083 18567 22089
rect 18509 22049 18521 22083
rect 18555 22080 18567 22083
rect 20346 22080 20352 22092
rect 18555 22052 20352 22080
rect 18555 22049 18567 22052
rect 18509 22043 18567 22049
rect 20346 22040 20352 22052
rect 20404 22040 20410 22092
rect 20548 22089 20576 22120
rect 20533 22083 20591 22089
rect 20533 22049 20545 22083
rect 20579 22049 20591 22083
rect 21174 22080 21180 22092
rect 21135 22052 21180 22080
rect 20533 22043 20591 22049
rect 21174 22040 21180 22052
rect 21232 22040 21238 22092
rect 17126 22012 17132 22024
rect 17087 21984 17132 22012
rect 17126 21972 17132 21984
rect 17184 21972 17190 22024
rect 18966 21972 18972 22024
rect 19024 22012 19030 22024
rect 21085 22015 21143 22021
rect 21085 22012 21097 22015
rect 19024 21984 21097 22012
rect 19024 21972 19030 21984
rect 21085 21981 21097 21984
rect 21131 22012 21143 22015
rect 21821 22015 21879 22021
rect 21821 22012 21833 22015
rect 21131 21984 21833 22012
rect 21131 21981 21143 21984
rect 21085 21975 21143 21981
rect 21821 21981 21833 21984
rect 21867 21981 21879 22015
rect 21821 21975 21879 21981
rect 37826 21972 37832 22024
rect 37884 22012 37890 22024
rect 38013 22015 38071 22021
rect 38013 22012 38025 22015
rect 37884 21984 38025 22012
rect 37884 21972 37890 21984
rect 38013 21981 38025 21984
rect 38059 21981 38071 22015
rect 38013 21975 38071 21981
rect 16546 21916 17172 21944
rect 15378 21876 15384 21888
rect 15120 21848 15384 21876
rect 12032 21836 12038 21848
rect 15378 21836 15384 21848
rect 15436 21836 15442 21888
rect 16022 21876 16028 21888
rect 15983 21848 16028 21876
rect 16022 21836 16028 21848
rect 16080 21836 16086 21888
rect 17034 21876 17040 21888
rect 16995 21848 17040 21876
rect 17034 21836 17040 21848
rect 17092 21836 17098 21888
rect 17144 21876 17172 21916
rect 17218 21904 17224 21956
rect 17276 21944 17282 21956
rect 17957 21947 18015 21953
rect 17957 21944 17969 21947
rect 17276 21916 17969 21944
rect 17276 21904 17282 21916
rect 17957 21913 17969 21916
rect 18003 21913 18015 21947
rect 17957 21907 18015 21913
rect 19426 21876 19432 21888
rect 17144 21848 19432 21876
rect 19426 21836 19432 21848
rect 19484 21836 19490 21888
rect 19978 21876 19984 21888
rect 19939 21848 19984 21876
rect 19978 21836 19984 21848
rect 20036 21836 20042 21888
rect 37366 21836 37372 21888
rect 37424 21876 37430 21888
rect 37829 21879 37887 21885
rect 37829 21876 37841 21879
rect 37424 21848 37841 21876
rect 37424 21836 37430 21848
rect 37829 21845 37841 21848
rect 37875 21845 37887 21879
rect 37829 21839 37887 21845
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 2498 21672 2504 21684
rect 2459 21644 2504 21672
rect 2498 21632 2504 21644
rect 2556 21632 2562 21684
rect 3053 21675 3111 21681
rect 3053 21641 3065 21675
rect 3099 21672 3111 21675
rect 3418 21672 3424 21684
rect 3099 21644 3424 21672
rect 3099 21641 3111 21644
rect 3053 21635 3111 21641
rect 3418 21632 3424 21644
rect 3476 21632 3482 21684
rect 3602 21672 3608 21684
rect 3563 21644 3608 21672
rect 3602 21632 3608 21644
rect 3660 21632 3666 21684
rect 4062 21632 4068 21684
rect 4120 21672 4126 21684
rect 4157 21675 4215 21681
rect 4157 21672 4169 21675
rect 4120 21644 4169 21672
rect 4120 21632 4126 21644
rect 4157 21641 4169 21644
rect 4203 21672 4215 21675
rect 4709 21675 4767 21681
rect 4709 21672 4721 21675
rect 4203 21644 4721 21672
rect 4203 21641 4215 21644
rect 4157 21635 4215 21641
rect 4709 21641 4721 21644
rect 4755 21672 4767 21675
rect 6454 21672 6460 21684
rect 4755 21644 6460 21672
rect 4755 21641 4767 21644
rect 4709 21635 4767 21641
rect 6454 21632 6460 21644
rect 6512 21672 6518 21684
rect 6549 21675 6607 21681
rect 6549 21672 6561 21675
rect 6512 21644 6561 21672
rect 6512 21632 6518 21644
rect 6549 21641 6561 21644
rect 6595 21641 6607 21675
rect 6549 21635 6607 21641
rect 9493 21675 9551 21681
rect 9493 21641 9505 21675
rect 9539 21672 9551 21675
rect 9674 21672 9680 21684
rect 9539 21644 9680 21672
rect 9539 21641 9551 21644
rect 9493 21635 9551 21641
rect 9674 21632 9680 21644
rect 9732 21632 9738 21684
rect 9766 21632 9772 21684
rect 9824 21672 9830 21684
rect 17034 21672 17040 21684
rect 9824 21644 12388 21672
rect 9824 21632 9830 21644
rect 5166 21604 5172 21616
rect 5127 21576 5172 21604
rect 5166 21564 5172 21576
rect 5224 21564 5230 21616
rect 8849 21607 8907 21613
rect 8849 21573 8861 21607
rect 8895 21604 8907 21607
rect 10686 21604 10692 21616
rect 8895 21576 10692 21604
rect 8895 21573 8907 21576
rect 8849 21567 8907 21573
rect 10686 21564 10692 21576
rect 10744 21564 10750 21616
rect 10962 21604 10968 21616
rect 10923 21576 10968 21604
rect 10962 21564 10968 21576
rect 11020 21564 11026 21616
rect 12360 21613 12388 21644
rect 14292 21644 17040 21672
rect 14292 21613 14320 21644
rect 17034 21632 17040 21644
rect 17092 21632 17098 21684
rect 18322 21672 18328 21684
rect 18283 21644 18328 21672
rect 18322 21632 18328 21644
rect 18380 21632 18386 21684
rect 19889 21675 19947 21681
rect 19889 21641 19901 21675
rect 19935 21672 19947 21675
rect 20162 21672 20168 21684
rect 19935 21644 20168 21672
rect 19935 21641 19947 21644
rect 19889 21635 19947 21641
rect 20162 21632 20168 21644
rect 20220 21632 20226 21684
rect 12345 21607 12403 21613
rect 12345 21573 12357 21607
rect 12391 21573 12403 21607
rect 12345 21567 12403 21573
rect 14277 21607 14335 21613
rect 14277 21573 14289 21607
rect 14323 21573 14335 21607
rect 14277 21567 14335 21573
rect 14369 21607 14427 21613
rect 14369 21573 14381 21607
rect 14415 21604 14427 21607
rect 15470 21604 15476 21616
rect 14415 21576 15476 21604
rect 14415 21573 14427 21576
rect 14369 21567 14427 21573
rect 15470 21564 15476 21576
rect 15528 21564 15534 21616
rect 15565 21607 15623 21613
rect 15565 21573 15577 21607
rect 15611 21604 15623 21607
rect 17129 21607 17187 21613
rect 17129 21604 17141 21607
rect 15611 21576 17141 21604
rect 15611 21573 15623 21576
rect 15565 21567 15623 21573
rect 17129 21573 17141 21576
rect 17175 21573 17187 21607
rect 17954 21604 17960 21616
rect 17129 21567 17187 21573
rect 17236 21576 17960 21604
rect 1854 21536 1860 21548
rect 1815 21508 1860 21536
rect 1854 21496 1860 21508
rect 1912 21496 1918 21548
rect 8113 21539 8171 21545
rect 8113 21536 8125 21539
rect 7576 21508 8125 21536
rect 1946 21428 1952 21480
rect 2004 21468 2010 21480
rect 7576 21477 7604 21508
rect 8113 21505 8125 21508
rect 8159 21505 8171 21539
rect 8113 21499 8171 21505
rect 8570 21496 8576 21548
rect 8628 21536 8634 21548
rect 8757 21539 8815 21545
rect 8757 21536 8769 21539
rect 8628 21508 8769 21536
rect 8628 21496 8634 21508
rect 8757 21505 8769 21508
rect 8803 21505 8815 21539
rect 9398 21536 9404 21548
rect 9359 21508 9404 21536
rect 8757 21499 8815 21505
rect 9398 21496 9404 21508
rect 9456 21496 9462 21548
rect 17236 21545 17264 21576
rect 17954 21564 17960 21576
rect 18012 21564 18018 21616
rect 21450 21604 21456 21616
rect 18432 21576 21456 21604
rect 17221 21539 17279 21545
rect 17221 21536 17233 21539
rect 15856 21508 17233 21536
rect 7561 21471 7619 21477
rect 7561 21468 7573 21471
rect 2004 21440 7573 21468
rect 2004 21428 2010 21440
rect 7561 21437 7573 21440
rect 7607 21437 7619 21471
rect 7561 21431 7619 21437
rect 9674 21428 9680 21480
rect 9732 21468 9738 21480
rect 10045 21471 10103 21477
rect 10045 21468 10057 21471
rect 9732 21440 10057 21468
rect 9732 21428 9738 21440
rect 10045 21437 10057 21440
rect 10091 21468 10103 21471
rect 10226 21468 10232 21480
rect 10091 21440 10232 21468
rect 10091 21437 10103 21440
rect 10045 21431 10103 21437
rect 10226 21428 10232 21440
rect 10284 21428 10290 21480
rect 11054 21468 11060 21480
rect 10967 21440 11060 21468
rect 11054 21428 11060 21440
rect 11112 21468 11118 21480
rect 11974 21468 11980 21480
rect 11112 21440 11980 21468
rect 11112 21428 11118 21440
rect 11974 21428 11980 21440
rect 12032 21428 12038 21480
rect 12253 21471 12311 21477
rect 12253 21437 12265 21471
rect 12299 21437 12311 21471
rect 12253 21431 12311 21437
rect 8205 21403 8263 21409
rect 8205 21369 8217 21403
rect 8251 21400 8263 21403
rect 11238 21400 11244 21412
rect 8251 21372 11244 21400
rect 8251 21369 8263 21372
rect 8205 21363 8263 21369
rect 11238 21360 11244 21372
rect 11296 21400 11302 21412
rect 12268 21400 12296 21431
rect 12434 21428 12440 21480
rect 12492 21468 12498 21480
rect 14093 21471 14151 21477
rect 12492 21440 12940 21468
rect 12492 21428 12498 21440
rect 12802 21400 12808 21412
rect 11296 21372 12296 21400
rect 12763 21372 12808 21400
rect 11296 21360 11302 21372
rect 12802 21360 12808 21372
rect 12860 21360 12866 21412
rect 12912 21400 12940 21440
rect 14093 21437 14105 21471
rect 14139 21468 14151 21471
rect 14274 21468 14280 21480
rect 14139 21440 14280 21468
rect 14139 21437 14151 21440
rect 14093 21431 14151 21437
rect 14274 21428 14280 21440
rect 14332 21428 14338 21480
rect 15010 21468 15016 21480
rect 14971 21440 15016 21468
rect 15010 21428 15016 21440
rect 15068 21428 15074 21480
rect 15654 21468 15660 21480
rect 15615 21440 15660 21468
rect 15654 21428 15660 21440
rect 15712 21428 15718 21480
rect 15856 21400 15884 21508
rect 17221 21505 17233 21508
rect 17267 21505 17279 21539
rect 17221 21499 17279 21505
rect 17678 21496 17684 21548
rect 17736 21536 17742 21548
rect 18432 21545 18460 21576
rect 21450 21564 21456 21576
rect 21508 21564 21514 21616
rect 18417 21539 18475 21545
rect 18417 21536 18429 21539
rect 17736 21508 18429 21536
rect 17736 21496 17742 21508
rect 18417 21505 18429 21508
rect 18463 21505 18475 21539
rect 18417 21499 18475 21505
rect 19058 21496 19064 21548
rect 19116 21536 19122 21548
rect 19797 21539 19855 21545
rect 19797 21536 19809 21539
rect 19116 21508 19809 21536
rect 19116 21496 19122 21508
rect 19797 21505 19809 21508
rect 19843 21536 19855 21539
rect 20441 21539 20499 21545
rect 20441 21536 20453 21539
rect 19843 21508 20453 21536
rect 19843 21505 19855 21508
rect 19797 21499 19855 21505
rect 20441 21505 20453 21508
rect 20487 21505 20499 21539
rect 38010 21536 38016 21548
rect 37971 21508 38016 21536
rect 20441 21499 20499 21505
rect 38010 21496 38016 21508
rect 38068 21496 38074 21548
rect 16022 21428 16028 21480
rect 16080 21468 16086 21480
rect 26510 21468 26516 21480
rect 16080 21440 26516 21468
rect 16080 21428 16086 21440
rect 26510 21428 26516 21440
rect 26568 21428 26574 21480
rect 12912 21372 15884 21400
rect 16301 21403 16359 21409
rect 16301 21369 16313 21403
rect 16347 21400 16359 21403
rect 17586 21400 17592 21412
rect 16347 21372 17592 21400
rect 16347 21369 16359 21372
rect 16301 21363 16359 21369
rect 17586 21360 17592 21372
rect 17644 21360 17650 21412
rect 17954 21360 17960 21412
rect 18012 21400 18018 21412
rect 18877 21403 18935 21409
rect 18877 21400 18889 21403
rect 18012 21372 18889 21400
rect 18012 21360 18018 21372
rect 18877 21369 18889 21372
rect 18923 21400 18935 21403
rect 18966 21400 18972 21412
rect 18923 21372 18972 21400
rect 18923 21369 18935 21372
rect 18877 21363 18935 21369
rect 18966 21360 18972 21372
rect 19024 21360 19030 21412
rect 1670 21332 1676 21344
rect 1631 21304 1676 21332
rect 1670 21292 1676 21304
rect 1728 21292 1734 21344
rect 10318 21292 10324 21344
rect 10376 21332 10382 21344
rect 15930 21332 15936 21344
rect 10376 21304 15936 21332
rect 10376 21292 10382 21304
rect 15930 21292 15936 21304
rect 15988 21292 15994 21344
rect 17678 21332 17684 21344
rect 17639 21304 17684 21332
rect 17678 21292 17684 21304
rect 17736 21292 17742 21344
rect 38194 21332 38200 21344
rect 38155 21304 38200 21332
rect 38194 21292 38200 21304
rect 38252 21292 38258 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 2222 21128 2228 21140
rect 2183 21100 2228 21128
rect 2222 21088 2228 21100
rect 2280 21088 2286 21140
rect 2777 21131 2835 21137
rect 2777 21097 2789 21131
rect 2823 21128 2835 21131
rect 3050 21128 3056 21140
rect 2823 21100 3056 21128
rect 2823 21097 2835 21100
rect 2777 21091 2835 21097
rect 3050 21088 3056 21100
rect 3108 21088 3114 21140
rect 4062 21128 4068 21140
rect 4023 21100 4068 21128
rect 4062 21088 4068 21100
rect 4120 21128 4126 21140
rect 4525 21131 4583 21137
rect 4525 21128 4537 21131
rect 4120 21100 4537 21128
rect 4120 21088 4126 21100
rect 4525 21097 4537 21100
rect 4571 21097 4583 21131
rect 4525 21091 4583 21097
rect 8110 21088 8116 21140
rect 8168 21128 8174 21140
rect 8481 21131 8539 21137
rect 8481 21128 8493 21131
rect 8168 21100 8493 21128
rect 8168 21088 8174 21100
rect 8481 21097 8493 21100
rect 8527 21128 8539 21131
rect 9490 21128 9496 21140
rect 8527 21100 9496 21128
rect 8527 21097 8539 21100
rect 8481 21091 8539 21097
rect 9490 21088 9496 21100
rect 9548 21088 9554 21140
rect 9585 21131 9643 21137
rect 9585 21097 9597 21131
rect 9631 21128 9643 21131
rect 10778 21128 10784 21140
rect 9631 21100 10784 21128
rect 9631 21097 9643 21100
rect 9585 21091 9643 21097
rect 10778 21088 10784 21100
rect 10836 21088 10842 21140
rect 11425 21131 11483 21137
rect 11425 21097 11437 21131
rect 11471 21128 11483 21131
rect 13262 21128 13268 21140
rect 11471 21100 13268 21128
rect 11471 21097 11483 21100
rect 11425 21091 11483 21097
rect 13262 21088 13268 21100
rect 13320 21128 13326 21140
rect 15562 21128 15568 21140
rect 13320 21100 15568 21128
rect 13320 21088 13326 21100
rect 15562 21088 15568 21100
rect 15620 21088 15626 21140
rect 15930 21088 15936 21140
rect 15988 21128 15994 21140
rect 19978 21128 19984 21140
rect 15988 21100 19984 21128
rect 15988 21088 15994 21100
rect 19978 21088 19984 21100
rect 20036 21088 20042 21140
rect 10226 21060 10232 21072
rect 10187 21032 10232 21060
rect 10226 21020 10232 21032
rect 10284 21020 10290 21072
rect 12802 21020 12808 21072
rect 12860 21060 12866 21072
rect 17494 21060 17500 21072
rect 12860 21032 17500 21060
rect 12860 21020 12866 21032
rect 17494 21020 17500 21032
rect 17552 21020 17558 21072
rect 18049 21063 18107 21069
rect 18049 21029 18061 21063
rect 18095 21060 18107 21063
rect 18230 21060 18236 21072
rect 18095 21032 18236 21060
rect 18095 21029 18107 21032
rect 18049 21023 18107 21029
rect 18230 21020 18236 21032
rect 18288 21020 18294 21072
rect 3421 20995 3479 21001
rect 3421 20961 3433 20995
rect 3467 20992 3479 20995
rect 6914 20992 6920 21004
rect 3467 20964 6920 20992
rect 3467 20961 3479 20964
rect 3421 20955 3479 20961
rect 6914 20952 6920 20964
rect 6972 20992 6978 21004
rect 12434 20992 12440 21004
rect 6972 20964 12440 20992
rect 6972 20952 6978 20964
rect 12434 20952 12440 20964
rect 12492 20952 12498 21004
rect 12529 20995 12587 21001
rect 12529 20961 12541 20995
rect 12575 20992 12587 20995
rect 13078 20992 13084 21004
rect 12575 20964 13084 20992
rect 12575 20961 12587 20964
rect 12529 20955 12587 20961
rect 13078 20952 13084 20964
rect 13136 20952 13142 21004
rect 13722 20992 13728 21004
rect 13683 20964 13728 20992
rect 13722 20952 13728 20964
rect 13780 20952 13786 21004
rect 14366 20952 14372 21004
rect 14424 20992 14430 21004
rect 14737 20995 14795 21001
rect 14737 20992 14749 20995
rect 14424 20964 14749 20992
rect 14424 20952 14430 20964
rect 14737 20961 14749 20964
rect 14783 20961 14795 20995
rect 14737 20955 14795 20961
rect 15381 20995 15439 21001
rect 15381 20961 15393 20995
rect 15427 20992 15439 20995
rect 15654 20992 15660 21004
rect 15427 20964 15660 20992
rect 15427 20961 15439 20964
rect 15381 20955 15439 20961
rect 15654 20952 15660 20964
rect 15712 20992 15718 21004
rect 16761 20995 16819 21001
rect 16761 20992 16773 20995
rect 15712 20964 16773 20992
rect 15712 20952 15718 20964
rect 16761 20961 16773 20964
rect 16807 20961 16819 20995
rect 16761 20955 16819 20961
rect 9490 20924 9496 20936
rect 9451 20896 9496 20924
rect 9490 20884 9496 20896
rect 9548 20884 9554 20936
rect 12345 20927 12403 20933
rect 12345 20893 12357 20927
rect 12391 20924 12403 20927
rect 12894 20924 12900 20936
rect 12391 20896 12900 20924
rect 12391 20893 12403 20896
rect 12345 20887 12403 20893
rect 12894 20884 12900 20896
rect 12952 20884 12958 20936
rect 16217 20927 16275 20933
rect 16217 20893 16229 20927
rect 16263 20924 16275 20927
rect 16850 20924 16856 20936
rect 16263 20896 16344 20924
rect 16811 20896 16856 20924
rect 16263 20893 16275 20896
rect 16217 20887 16275 20893
rect 10689 20859 10747 20865
rect 10689 20825 10701 20859
rect 10735 20825 10747 20859
rect 10689 20819 10747 20825
rect 9950 20748 9956 20800
rect 10008 20788 10014 20800
rect 10704 20788 10732 20819
rect 10778 20816 10784 20868
rect 10836 20856 10842 20868
rect 10836 20828 10881 20856
rect 10836 20816 10842 20828
rect 12618 20816 12624 20868
rect 12676 20856 12682 20868
rect 13081 20859 13139 20865
rect 13081 20856 13093 20859
rect 12676 20828 13093 20856
rect 12676 20816 12682 20828
rect 13081 20825 13093 20828
rect 13127 20825 13139 20859
rect 13081 20819 13139 20825
rect 13170 20816 13176 20868
rect 13228 20856 13234 20868
rect 15289 20859 15347 20865
rect 13228 20828 13273 20856
rect 13228 20816 13234 20828
rect 15289 20825 15301 20859
rect 15335 20825 15347 20859
rect 15289 20819 15347 20825
rect 16316 20856 16344 20896
rect 16850 20884 16856 20896
rect 16908 20884 16914 20936
rect 17494 20924 17500 20936
rect 17455 20896 17500 20924
rect 17494 20884 17500 20896
rect 17552 20884 17558 20936
rect 18785 20927 18843 20933
rect 18785 20893 18797 20927
rect 18831 20924 18843 20927
rect 18874 20924 18880 20936
rect 18831 20896 18880 20924
rect 18831 20893 18843 20896
rect 18785 20887 18843 20893
rect 18874 20884 18880 20896
rect 18932 20924 18938 20936
rect 19429 20927 19487 20933
rect 19429 20924 19441 20927
rect 18932 20896 19441 20924
rect 18932 20884 18938 20896
rect 19429 20893 19441 20896
rect 19475 20893 19487 20927
rect 19429 20887 19487 20893
rect 16942 20856 16948 20868
rect 16316 20828 16948 20856
rect 10008 20760 10732 20788
rect 11885 20791 11943 20797
rect 10008 20748 10014 20760
rect 11885 20757 11897 20791
rect 11931 20788 11943 20791
rect 11974 20788 11980 20800
rect 11931 20760 11980 20788
rect 11931 20757 11943 20760
rect 11885 20751 11943 20757
rect 11974 20748 11980 20760
rect 12032 20748 12038 20800
rect 15304 20788 15332 20819
rect 16117 20791 16175 20797
rect 16117 20788 16129 20791
rect 15304 20760 16129 20788
rect 16117 20757 16129 20760
rect 16163 20757 16175 20791
rect 16117 20751 16175 20757
rect 16206 20748 16212 20800
rect 16264 20788 16270 20800
rect 16316 20788 16344 20828
rect 16942 20816 16948 20828
rect 17000 20856 17006 20868
rect 19058 20856 19064 20868
rect 17000 20828 19064 20856
rect 17000 20816 17006 20828
rect 19058 20816 19064 20828
rect 19116 20816 19122 20868
rect 17310 20788 17316 20800
rect 16264 20760 16344 20788
rect 17271 20760 17316 20788
rect 16264 20748 16270 20760
rect 17310 20748 17316 20760
rect 17368 20748 17374 20800
rect 18690 20788 18696 20800
rect 18651 20760 18696 20788
rect 18690 20748 18696 20760
rect 18748 20748 18754 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 3605 20587 3663 20593
rect 3605 20553 3617 20587
rect 3651 20584 3663 20587
rect 5074 20584 5080 20596
rect 3651 20556 5080 20584
rect 3651 20553 3663 20556
rect 3605 20547 3663 20553
rect 5074 20544 5080 20556
rect 5132 20544 5138 20596
rect 9858 20584 9864 20596
rect 9819 20556 9864 20584
rect 9858 20544 9864 20556
rect 9916 20544 9922 20596
rect 11793 20587 11851 20593
rect 11793 20553 11805 20587
rect 11839 20584 11851 20587
rect 12342 20584 12348 20596
rect 11839 20556 12348 20584
rect 11839 20553 11851 20556
rect 11793 20547 11851 20553
rect 12342 20544 12348 20556
rect 12400 20584 12406 20596
rect 13538 20584 13544 20596
rect 12400 20556 13124 20584
rect 13499 20556 13544 20584
rect 12400 20544 12406 20556
rect 10870 20516 10876 20528
rect 9784 20488 10876 20516
rect 9784 20460 9812 20488
rect 10870 20476 10876 20488
rect 10928 20476 10934 20528
rect 10965 20519 11023 20525
rect 10965 20485 10977 20519
rect 11011 20516 11023 20519
rect 11054 20516 11060 20528
rect 11011 20488 11060 20516
rect 11011 20485 11023 20488
rect 10965 20479 11023 20485
rect 11054 20476 11060 20488
rect 11112 20476 11118 20528
rect 12066 20476 12072 20528
rect 12124 20516 12130 20528
rect 12253 20519 12311 20525
rect 12253 20516 12265 20519
rect 12124 20488 12265 20516
rect 12124 20476 12130 20488
rect 12253 20485 12265 20488
rect 12299 20485 12311 20519
rect 12802 20516 12808 20528
rect 12763 20488 12808 20516
rect 12253 20479 12311 20485
rect 12802 20476 12808 20488
rect 12860 20476 12866 20528
rect 9766 20448 9772 20460
rect 9679 20420 9772 20448
rect 9766 20408 9772 20420
rect 9824 20408 9830 20460
rect 13096 20448 13124 20556
rect 13538 20544 13544 20556
rect 13596 20544 13602 20596
rect 15378 20584 15384 20596
rect 13740 20556 15240 20584
rect 15339 20556 15384 20584
rect 13740 20528 13768 20556
rect 13262 20476 13268 20528
rect 13320 20516 13326 20528
rect 13722 20516 13728 20528
rect 13320 20488 13728 20516
rect 13320 20476 13326 20488
rect 13722 20476 13728 20488
rect 13780 20476 13786 20528
rect 14274 20516 14280 20528
rect 14235 20488 14280 20516
rect 14274 20476 14280 20488
rect 14332 20476 14338 20528
rect 15212 20516 15240 20556
rect 15378 20544 15384 20556
rect 15436 20544 15442 20596
rect 15470 20544 15476 20596
rect 15528 20584 15534 20596
rect 16945 20587 17003 20593
rect 16945 20584 16957 20587
rect 15528 20556 16957 20584
rect 15528 20544 15534 20556
rect 16945 20553 16957 20556
rect 16991 20553 17003 20587
rect 16945 20547 17003 20553
rect 17126 20544 17132 20596
rect 17184 20584 17190 20596
rect 17497 20587 17555 20593
rect 17497 20584 17509 20587
rect 17184 20556 17509 20584
rect 17184 20544 17190 20556
rect 17497 20553 17509 20556
rect 17543 20553 17555 20587
rect 17497 20547 17555 20553
rect 18693 20587 18751 20593
rect 18693 20553 18705 20587
rect 18739 20584 18751 20587
rect 19150 20584 19156 20596
rect 18739 20556 19156 20584
rect 18739 20553 18751 20556
rect 18693 20547 18751 20553
rect 16025 20519 16083 20525
rect 15212 20488 15976 20516
rect 13449 20451 13507 20457
rect 13449 20448 13461 20451
rect 13096 20420 13461 20448
rect 13449 20417 13461 20420
rect 13495 20417 13507 20451
rect 13449 20411 13507 20417
rect 15473 20451 15531 20457
rect 15473 20417 15485 20451
rect 15519 20448 15531 20451
rect 15838 20448 15844 20460
rect 15519 20420 15844 20448
rect 15519 20417 15531 20420
rect 15473 20411 15531 20417
rect 15838 20408 15844 20420
rect 15896 20408 15902 20460
rect 15948 20457 15976 20488
rect 16025 20485 16037 20519
rect 16071 20516 16083 20519
rect 16114 20516 16120 20528
rect 16071 20488 16120 20516
rect 16071 20485 16083 20488
rect 16025 20479 16083 20485
rect 16114 20476 16120 20488
rect 16172 20476 16178 20528
rect 15933 20451 15991 20457
rect 15933 20417 15945 20451
rect 15979 20417 15991 20451
rect 15933 20411 15991 20417
rect 17037 20451 17095 20457
rect 17037 20417 17049 20451
rect 17083 20448 17095 20451
rect 17494 20448 17500 20460
rect 17083 20420 17500 20448
rect 17083 20417 17095 20420
rect 17037 20411 17095 20417
rect 17494 20408 17500 20420
rect 17552 20448 17558 20460
rect 17862 20448 17868 20460
rect 17552 20420 17868 20448
rect 17552 20408 17558 20420
rect 17862 20408 17868 20420
rect 17920 20408 17926 20460
rect 10778 20380 10784 20392
rect 10691 20352 10784 20380
rect 10778 20340 10784 20352
rect 10836 20340 10842 20392
rect 11057 20383 11115 20389
rect 11057 20349 11069 20383
rect 11103 20380 11115 20383
rect 11238 20380 11244 20392
rect 11103 20352 11244 20380
rect 11103 20349 11115 20352
rect 11057 20343 11115 20349
rect 11238 20340 11244 20352
rect 11296 20340 11302 20392
rect 12897 20383 12955 20389
rect 12897 20349 12909 20383
rect 12943 20349 12955 20383
rect 14182 20380 14188 20392
rect 14143 20352 14188 20380
rect 12897 20343 12955 20349
rect 10796 20312 10824 20340
rect 12912 20312 12940 20343
rect 14182 20340 14188 20352
rect 14240 20340 14246 20392
rect 14366 20340 14372 20392
rect 14424 20380 14430 20392
rect 14461 20383 14519 20389
rect 14461 20380 14473 20383
rect 14424 20352 14473 20380
rect 14424 20340 14430 20352
rect 14461 20349 14473 20352
rect 14507 20349 14519 20383
rect 15856 20380 15884 20408
rect 18708 20380 18736 20547
rect 19150 20544 19156 20556
rect 19208 20544 19214 20596
rect 37829 20451 37887 20457
rect 37829 20417 37841 20451
rect 37875 20448 37887 20451
rect 37918 20448 37924 20460
rect 37875 20420 37924 20448
rect 37875 20417 37887 20420
rect 37829 20411 37887 20417
rect 37918 20408 37924 20420
rect 37976 20408 37982 20460
rect 15856 20352 18736 20380
rect 14461 20343 14519 20349
rect 13262 20312 13268 20324
rect 10796 20284 12434 20312
rect 12912 20284 13268 20312
rect 9309 20247 9367 20253
rect 9309 20213 9321 20247
rect 9355 20244 9367 20247
rect 9398 20244 9404 20256
rect 9355 20216 9404 20244
rect 9355 20213 9367 20216
rect 9309 20207 9367 20213
rect 9398 20204 9404 20216
rect 9456 20204 9462 20256
rect 12406 20244 12434 20284
rect 13262 20272 13268 20284
rect 13320 20312 13326 20324
rect 14918 20312 14924 20324
rect 13320 20284 14924 20312
rect 13320 20272 13326 20284
rect 14918 20272 14924 20284
rect 14976 20272 14982 20324
rect 14826 20244 14832 20256
rect 12406 20216 14832 20244
rect 14826 20204 14832 20216
rect 14884 20204 14890 20256
rect 17862 20204 17868 20256
rect 17920 20244 17926 20256
rect 18049 20247 18107 20253
rect 18049 20244 18061 20247
rect 17920 20216 18061 20244
rect 17920 20204 17926 20216
rect 18049 20213 18061 20216
rect 18095 20213 18107 20247
rect 18049 20207 18107 20213
rect 38013 20247 38071 20253
rect 38013 20213 38025 20247
rect 38059 20244 38071 20247
rect 38102 20244 38108 20256
rect 38059 20216 38108 20244
rect 38059 20213 38071 20216
rect 38013 20207 38071 20213
rect 38102 20204 38108 20216
rect 38160 20204 38166 20256
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 9309 20043 9367 20049
rect 9309 20009 9321 20043
rect 9355 20040 9367 20043
rect 9766 20040 9772 20052
rect 9355 20012 9772 20040
rect 9355 20009 9367 20012
rect 9309 20003 9367 20009
rect 9766 20000 9772 20012
rect 9824 20000 9830 20052
rect 9861 20043 9919 20049
rect 9861 20009 9873 20043
rect 9907 20040 9919 20043
rect 11146 20040 11152 20052
rect 9907 20012 11152 20040
rect 9907 20009 9919 20012
rect 9861 20003 9919 20009
rect 11146 20000 11152 20012
rect 11204 20000 11210 20052
rect 11256 20012 13492 20040
rect 9398 19932 9404 19984
rect 9456 19972 9462 19984
rect 11256 19972 11284 20012
rect 9456 19944 11284 19972
rect 12345 19975 12403 19981
rect 9456 19932 9462 19944
rect 12345 19941 12357 19975
rect 12391 19972 12403 19975
rect 13354 19972 13360 19984
rect 12391 19944 13360 19972
rect 12391 19941 12403 19944
rect 12345 19935 12403 19941
rect 13354 19932 13360 19944
rect 13412 19932 13418 19984
rect 13464 19972 13492 20012
rect 13722 20000 13728 20052
rect 13780 20040 13786 20052
rect 14277 20043 14335 20049
rect 14277 20040 14289 20043
rect 13780 20012 14289 20040
rect 13780 20000 13786 20012
rect 14277 20009 14289 20012
rect 14323 20009 14335 20043
rect 14277 20003 14335 20009
rect 16117 20043 16175 20049
rect 16117 20009 16129 20043
rect 16163 20040 16175 20043
rect 16298 20040 16304 20052
rect 16163 20012 16304 20040
rect 16163 20009 16175 20012
rect 16117 20003 16175 20009
rect 16298 20000 16304 20012
rect 16356 20000 16362 20052
rect 16945 20043 17003 20049
rect 16945 20009 16957 20043
rect 16991 20040 17003 20043
rect 17954 20040 17960 20052
rect 16991 20012 17960 20040
rect 16991 20009 17003 20012
rect 16945 20003 17003 20009
rect 17954 20000 17960 20012
rect 18012 20000 18018 20052
rect 21450 20040 21456 20052
rect 21411 20012 21456 20040
rect 21450 20000 21456 20012
rect 21508 20000 21514 20052
rect 23290 19972 23296 19984
rect 13464 19944 23296 19972
rect 23290 19932 23296 19944
rect 23348 19932 23354 19984
rect 11422 19904 11428 19916
rect 7300 19876 11428 19904
rect 7300 19845 7328 19876
rect 11422 19864 11428 19876
rect 11480 19864 11486 19916
rect 11793 19907 11851 19913
rect 11793 19873 11805 19907
rect 11839 19904 11851 19907
rect 12618 19904 12624 19916
rect 11839 19876 12624 19904
rect 11839 19873 11851 19876
rect 11793 19867 11851 19873
rect 12618 19864 12624 19876
rect 12676 19864 12682 19916
rect 13725 19907 13783 19913
rect 13725 19873 13737 19907
rect 13771 19904 13783 19907
rect 14550 19904 14556 19916
rect 13771 19876 14556 19904
rect 13771 19873 13783 19876
rect 13725 19867 13783 19873
rect 14550 19864 14556 19876
rect 14608 19864 14614 19916
rect 15473 19907 15531 19913
rect 15473 19873 15485 19907
rect 15519 19904 15531 19907
rect 16482 19904 16488 19916
rect 15519 19876 16488 19904
rect 15519 19873 15531 19876
rect 15473 19867 15531 19873
rect 16482 19864 16488 19876
rect 16540 19864 16546 19916
rect 16850 19864 16856 19916
rect 16908 19904 16914 19916
rect 17497 19907 17555 19913
rect 17497 19904 17509 19907
rect 16908 19876 17509 19904
rect 16908 19864 16914 19876
rect 17497 19873 17509 19876
rect 17543 19904 17555 19907
rect 22281 19907 22339 19913
rect 17543 19876 22232 19904
rect 17543 19873 17555 19876
rect 17497 19867 17555 19873
rect 7285 19839 7343 19845
rect 7285 19805 7297 19839
rect 7331 19805 7343 19839
rect 7285 19799 7343 19805
rect 7834 19796 7840 19848
rect 7892 19836 7898 19848
rect 9769 19839 9827 19845
rect 9769 19836 9781 19839
rect 7892 19808 9781 19836
rect 7892 19796 7898 19808
rect 9769 19805 9781 19808
rect 9815 19836 9827 19839
rect 10134 19836 10140 19848
rect 9815 19808 10140 19836
rect 9815 19805 9827 19808
rect 9769 19799 9827 19805
rect 10134 19796 10140 19808
rect 10192 19836 10198 19848
rect 10413 19839 10471 19845
rect 10413 19836 10425 19839
rect 10192 19808 10425 19836
rect 10192 19796 10198 19808
rect 10413 19805 10425 19808
rect 10459 19805 10471 19839
rect 10413 19799 10471 19805
rect 10870 19796 10876 19848
rect 10928 19836 10934 19848
rect 11057 19839 11115 19845
rect 11057 19836 11069 19839
rect 10928 19808 11069 19836
rect 10928 19796 10934 19808
rect 11057 19805 11069 19808
rect 11103 19805 11115 19839
rect 11057 19799 11115 19805
rect 15746 19796 15752 19848
rect 15804 19836 15810 19848
rect 16025 19839 16083 19845
rect 16025 19836 16037 19839
rect 15804 19808 16037 19836
rect 15804 19796 15810 19808
rect 16025 19805 16037 19808
rect 16071 19805 16083 19839
rect 16025 19799 16083 19805
rect 21450 19796 21456 19848
rect 21508 19836 21514 19848
rect 22097 19839 22155 19845
rect 22097 19836 22109 19839
rect 21508 19808 22109 19836
rect 21508 19796 21514 19808
rect 22097 19805 22109 19808
rect 22143 19805 22155 19839
rect 22097 19799 22155 19805
rect 10505 19771 10563 19777
rect 10505 19737 10517 19771
rect 10551 19768 10563 19771
rect 11422 19768 11428 19780
rect 10551 19740 11428 19768
rect 10551 19737 10563 19740
rect 10505 19731 10563 19737
rect 11422 19728 11428 19740
rect 11480 19728 11486 19780
rect 11885 19771 11943 19777
rect 11885 19737 11897 19771
rect 11931 19737 11943 19771
rect 13078 19768 13084 19780
rect 13039 19740 13084 19768
rect 11885 19731 11943 19737
rect 1854 19660 1860 19712
rect 1912 19700 1918 19712
rect 7193 19703 7251 19709
rect 7193 19700 7205 19703
rect 1912 19672 7205 19700
rect 1912 19660 1918 19672
rect 7193 19669 7205 19672
rect 7239 19669 7251 19703
rect 7193 19663 7251 19669
rect 11149 19703 11207 19709
rect 11149 19669 11161 19703
rect 11195 19700 11207 19703
rect 11900 19700 11928 19731
rect 13078 19728 13084 19740
rect 13136 19728 13142 19780
rect 13173 19771 13231 19777
rect 13173 19737 13185 19771
rect 13219 19768 13231 19771
rect 13538 19768 13544 19780
rect 13219 19740 13544 19768
rect 13219 19737 13231 19740
rect 13173 19731 13231 19737
rect 13538 19728 13544 19740
rect 13596 19728 13602 19780
rect 14826 19768 14832 19780
rect 13832 19740 14412 19768
rect 14787 19740 14832 19768
rect 11195 19672 11928 19700
rect 11195 19669 11207 19672
rect 11149 19663 11207 19669
rect 13630 19660 13636 19712
rect 13688 19700 13694 19712
rect 13832 19700 13860 19740
rect 13688 19672 13860 19700
rect 14384 19700 14412 19740
rect 14826 19728 14832 19740
rect 14884 19728 14890 19780
rect 15286 19728 15292 19780
rect 15344 19768 15350 19780
rect 15381 19771 15439 19777
rect 15381 19768 15393 19771
rect 15344 19740 15393 19768
rect 15344 19728 15350 19740
rect 15381 19737 15393 19740
rect 15427 19737 15439 19771
rect 15381 19731 15439 19737
rect 17862 19728 17868 19780
rect 17920 19768 17926 19780
rect 18049 19771 18107 19777
rect 18049 19768 18061 19771
rect 17920 19740 18061 19768
rect 17920 19728 17926 19740
rect 18049 19737 18061 19740
rect 18095 19768 18107 19771
rect 22204 19768 22232 19876
rect 22281 19873 22293 19907
rect 22327 19904 22339 19907
rect 37458 19904 37464 19916
rect 22327 19876 37464 19904
rect 22327 19873 22339 19876
rect 22281 19867 22339 19873
rect 37458 19864 37464 19876
rect 37516 19864 37522 19916
rect 36538 19796 36544 19848
rect 36596 19836 36602 19848
rect 38013 19839 38071 19845
rect 38013 19836 38025 19839
rect 36596 19808 38025 19836
rect 36596 19796 36602 19808
rect 38013 19805 38025 19808
rect 38059 19805 38071 19839
rect 38013 19799 38071 19805
rect 33686 19768 33692 19780
rect 18095 19740 21588 19768
rect 22204 19740 33692 19768
rect 18095 19737 18107 19740
rect 18049 19731 18107 19737
rect 16298 19700 16304 19712
rect 14384 19672 16304 19700
rect 13688 19660 13694 19672
rect 16298 19660 16304 19672
rect 16356 19660 16362 19712
rect 21560 19700 21588 19740
rect 33686 19728 33692 19740
rect 33744 19728 33750 19780
rect 36722 19700 36728 19712
rect 21560 19672 36728 19700
rect 36722 19660 36728 19672
rect 36780 19660 36786 19712
rect 38194 19700 38200 19712
rect 38155 19672 38200 19700
rect 38194 19660 38200 19672
rect 38252 19660 38258 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 10505 19499 10563 19505
rect 10505 19465 10517 19499
rect 10551 19496 10563 19499
rect 10870 19496 10876 19508
rect 10551 19468 10876 19496
rect 10551 19465 10563 19468
rect 10505 19459 10563 19465
rect 10870 19456 10876 19468
rect 10928 19456 10934 19508
rect 11054 19496 11060 19508
rect 11015 19468 11060 19496
rect 11054 19456 11060 19468
rect 11112 19456 11118 19508
rect 11974 19496 11980 19508
rect 11935 19468 11980 19496
rect 11974 19456 11980 19468
rect 12032 19456 12038 19508
rect 13538 19496 13544 19508
rect 13499 19468 13544 19496
rect 13538 19456 13544 19468
rect 13596 19456 13602 19508
rect 16209 19499 16267 19505
rect 16209 19496 16221 19499
rect 14292 19468 16221 19496
rect 13722 19428 13728 19440
rect 12406 19400 13728 19428
rect 1854 19360 1860 19372
rect 1815 19332 1860 19360
rect 1854 19320 1860 19332
rect 1912 19320 1918 19372
rect 11149 19363 11207 19369
rect 11149 19329 11161 19363
rect 11195 19360 11207 19363
rect 12406 19360 12434 19400
rect 13722 19388 13728 19400
rect 13780 19388 13786 19440
rect 14182 19428 14188 19440
rect 14143 19400 14188 19428
rect 14182 19388 14188 19400
rect 14240 19388 14246 19440
rect 14292 19437 14320 19468
rect 16209 19465 16221 19468
rect 16255 19465 16267 19499
rect 16209 19459 16267 19465
rect 16298 19456 16304 19508
rect 16356 19496 16362 19508
rect 22738 19496 22744 19508
rect 16356 19468 22744 19496
rect 16356 19456 16362 19468
rect 22738 19456 22744 19468
rect 22796 19456 22802 19508
rect 14277 19431 14335 19437
rect 14277 19397 14289 19431
rect 14323 19397 14335 19431
rect 14277 19391 14335 19397
rect 15565 19431 15623 19437
rect 15565 19397 15577 19431
rect 15611 19428 15623 19431
rect 15611 19400 16574 19428
rect 15611 19397 15623 19400
rect 15565 19391 15623 19397
rect 12618 19360 12624 19372
rect 11195 19332 12434 19360
rect 12579 19332 12624 19360
rect 11195 19329 11207 19332
rect 11149 19323 11207 19329
rect 9953 19295 10011 19301
rect 9953 19261 9965 19295
rect 9999 19292 10011 19295
rect 11164 19292 11192 19323
rect 12618 19320 12624 19332
rect 12676 19320 12682 19372
rect 13630 19360 13636 19372
rect 13591 19332 13636 19360
rect 13630 19320 13636 19332
rect 13688 19320 13694 19372
rect 15473 19363 15531 19369
rect 15473 19360 15485 19363
rect 15212 19332 15485 19360
rect 9999 19264 11192 19292
rect 9999 19261 10011 19264
rect 9953 19255 10011 19261
rect 11422 19252 11428 19304
rect 11480 19292 11486 19304
rect 12437 19295 12495 19301
rect 12437 19292 12449 19295
rect 11480 19264 12449 19292
rect 11480 19252 11486 19264
rect 12437 19261 12449 19264
rect 12483 19261 12495 19295
rect 12437 19255 12495 19261
rect 14829 19295 14887 19301
rect 14829 19261 14841 19295
rect 14875 19292 14887 19295
rect 15010 19292 15016 19304
rect 14875 19264 15016 19292
rect 14875 19261 14887 19264
rect 14829 19255 14887 19261
rect 15010 19252 15016 19264
rect 15068 19252 15074 19304
rect 12986 19184 12992 19236
rect 13044 19224 13050 19236
rect 15212 19224 15240 19332
rect 15473 19329 15485 19332
rect 15519 19329 15531 19363
rect 15473 19323 15531 19329
rect 15746 19320 15752 19372
rect 15804 19360 15810 19372
rect 16301 19363 16359 19369
rect 16301 19360 16313 19363
rect 15804 19332 16313 19360
rect 15804 19320 15810 19332
rect 16301 19329 16313 19332
rect 16347 19329 16359 19363
rect 16546 19360 16574 19400
rect 17218 19360 17224 19372
rect 16546 19332 17224 19360
rect 16301 19323 16359 19329
rect 15286 19224 15292 19236
rect 13044 19196 15292 19224
rect 13044 19184 13050 19196
rect 15286 19184 15292 19196
rect 15344 19184 15350 19236
rect 16316 19224 16344 19323
rect 17218 19320 17224 19332
rect 17276 19320 17282 19372
rect 16945 19227 17003 19233
rect 16945 19224 16957 19227
rect 16316 19196 16957 19224
rect 16945 19193 16957 19196
rect 16991 19224 17003 19227
rect 17405 19227 17463 19233
rect 17405 19224 17417 19227
rect 16991 19196 17417 19224
rect 16991 19193 17003 19196
rect 16945 19187 17003 19193
rect 17405 19193 17417 19196
rect 17451 19193 17463 19227
rect 17405 19187 17463 19193
rect 1670 19156 1676 19168
rect 1631 19128 1676 19156
rect 1670 19116 1676 19128
rect 1728 19116 1734 19168
rect 11330 19116 11336 19168
rect 11388 19156 11394 19168
rect 14642 19156 14648 19168
rect 11388 19128 14648 19156
rect 11388 19116 11394 19128
rect 14642 19116 14648 19128
rect 14700 19116 14706 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 4709 18955 4767 18961
rect 4709 18921 4721 18955
rect 4755 18952 4767 18955
rect 7098 18952 7104 18964
rect 4755 18924 7104 18952
rect 4755 18921 4767 18924
rect 4709 18915 4767 18921
rect 4157 18751 4215 18757
rect 4157 18717 4169 18751
rect 4203 18748 4215 18751
rect 4724 18748 4752 18915
rect 7098 18912 7104 18924
rect 7156 18912 7162 18964
rect 10134 18952 10140 18964
rect 10095 18924 10140 18952
rect 10134 18912 10140 18924
rect 10192 18952 10198 18964
rect 10689 18955 10747 18961
rect 10689 18952 10701 18955
rect 10192 18924 10701 18952
rect 10192 18912 10198 18924
rect 10689 18921 10701 18924
rect 10735 18921 10747 18955
rect 10689 18915 10747 18921
rect 12618 18912 12624 18964
rect 12676 18952 12682 18964
rect 12713 18955 12771 18961
rect 12713 18952 12725 18955
rect 12676 18924 12725 18952
rect 12676 18912 12682 18924
rect 12713 18921 12725 18924
rect 12759 18921 12771 18955
rect 12713 18915 12771 18921
rect 12894 18912 12900 18964
rect 12952 18952 12958 18964
rect 13449 18955 13507 18961
rect 13449 18952 13461 18955
rect 12952 18924 13461 18952
rect 12952 18912 12958 18924
rect 13449 18921 13461 18924
rect 13495 18921 13507 18955
rect 13449 18915 13507 18921
rect 14182 18912 14188 18964
rect 14240 18952 14246 18964
rect 14553 18955 14611 18961
rect 14553 18952 14565 18955
rect 14240 18924 14565 18952
rect 14240 18912 14246 18924
rect 14553 18921 14565 18924
rect 14599 18921 14611 18955
rect 15194 18952 15200 18964
rect 15155 18924 15200 18952
rect 14553 18915 14611 18921
rect 15194 18912 15200 18924
rect 15252 18912 15258 18964
rect 15933 18955 15991 18961
rect 15933 18921 15945 18955
rect 15979 18952 15991 18955
rect 16206 18952 16212 18964
rect 15979 18924 16212 18952
rect 15979 18921 15991 18924
rect 15933 18915 15991 18921
rect 16206 18912 16212 18924
rect 16264 18912 16270 18964
rect 16482 18952 16488 18964
rect 16443 18924 16488 18952
rect 16482 18912 16488 18924
rect 16540 18912 16546 18964
rect 12161 18887 12219 18893
rect 12161 18853 12173 18887
rect 12207 18884 12219 18887
rect 13630 18884 13636 18896
rect 12207 18856 13636 18884
rect 12207 18853 12219 18856
rect 12161 18847 12219 18853
rect 13630 18844 13636 18856
rect 13688 18844 13694 18896
rect 13740 18856 16574 18884
rect 9490 18776 9496 18828
rect 9548 18816 9554 18828
rect 11606 18816 11612 18828
rect 9548 18788 11612 18816
rect 9548 18776 9554 18788
rect 11606 18776 11612 18788
rect 11664 18776 11670 18828
rect 13740 18816 13768 18856
rect 12820 18788 13768 18816
rect 4203 18720 4752 18748
rect 4203 18717 4215 18720
rect 4157 18711 4215 18717
rect 11514 18708 11520 18760
rect 11572 18748 11578 18760
rect 12820 18757 12848 18788
rect 13906 18776 13912 18828
rect 13964 18816 13970 18828
rect 15102 18816 15108 18828
rect 13964 18788 15108 18816
rect 13964 18776 13970 18788
rect 15102 18776 15108 18788
rect 15160 18816 15166 18828
rect 16546 18816 16574 18856
rect 20898 18816 20904 18828
rect 15160 18788 15332 18816
rect 16546 18788 20904 18816
rect 15160 18776 15166 18788
rect 12805 18751 12863 18757
rect 12805 18748 12817 18751
rect 11572 18720 12817 18748
rect 11572 18708 11578 18720
rect 12805 18717 12817 18720
rect 12851 18717 12863 18751
rect 13538 18748 13544 18760
rect 13499 18720 13544 18748
rect 12805 18711 12863 18717
rect 13538 18708 13544 18720
rect 13596 18708 13602 18760
rect 14642 18748 14648 18760
rect 14603 18720 14648 18748
rect 14642 18708 14648 18720
rect 14700 18748 14706 18760
rect 15194 18748 15200 18760
rect 14700 18720 15200 18748
rect 14700 18708 14706 18720
rect 15194 18708 15200 18720
rect 15252 18708 15258 18760
rect 15304 18757 15332 18788
rect 20898 18776 20904 18788
rect 20956 18776 20962 18828
rect 15289 18751 15347 18757
rect 15289 18717 15301 18751
rect 15335 18717 15347 18751
rect 15289 18711 15347 18717
rect 7466 18640 7472 18692
rect 7524 18680 7530 18692
rect 17310 18680 17316 18692
rect 7524 18652 17316 18680
rect 7524 18640 7530 18652
rect 17310 18640 17316 18652
rect 17368 18640 17374 18692
rect 3970 18612 3976 18624
rect 3931 18584 3976 18612
rect 3970 18572 3976 18584
rect 4028 18572 4034 18624
rect 11514 18612 11520 18624
rect 11475 18584 11520 18612
rect 11514 18572 11520 18584
rect 11572 18572 11578 18624
rect 11606 18572 11612 18624
rect 11664 18612 11670 18624
rect 12986 18612 12992 18624
rect 11664 18584 12992 18612
rect 11664 18572 11670 18584
rect 12986 18572 12992 18584
rect 13044 18612 13050 18624
rect 13722 18612 13728 18624
rect 13044 18584 13728 18612
rect 13044 18572 13050 18584
rect 13722 18572 13728 18584
rect 13780 18572 13786 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 2409 18411 2467 18417
rect 2409 18377 2421 18411
rect 2455 18408 2467 18411
rect 7466 18408 7472 18420
rect 2455 18380 7472 18408
rect 2455 18377 2467 18380
rect 2409 18371 2467 18377
rect 1857 18275 1915 18281
rect 1857 18241 1869 18275
rect 1903 18272 1915 18275
rect 2424 18272 2452 18371
rect 7466 18368 7472 18380
rect 7524 18368 7530 18420
rect 12802 18368 12808 18420
rect 12860 18408 12866 18420
rect 12989 18411 13047 18417
rect 12989 18408 13001 18411
rect 12860 18380 13001 18408
rect 12860 18368 12866 18380
rect 12989 18377 13001 18380
rect 13035 18377 13047 18411
rect 12989 18371 13047 18377
rect 13170 18368 13176 18420
rect 13228 18408 13234 18420
rect 13633 18411 13691 18417
rect 13633 18408 13645 18411
rect 13228 18380 13645 18408
rect 13228 18368 13234 18380
rect 13633 18377 13645 18380
rect 13679 18377 13691 18411
rect 13633 18371 13691 18377
rect 14274 18368 14280 18420
rect 14332 18408 14338 18420
rect 14553 18411 14611 18417
rect 14553 18408 14565 18411
rect 14332 18380 14565 18408
rect 14332 18368 14338 18380
rect 14553 18377 14565 18380
rect 14599 18377 14611 18411
rect 14553 18371 14611 18377
rect 15102 18368 15108 18420
rect 15160 18408 15166 18420
rect 15841 18411 15899 18417
rect 15841 18408 15853 18411
rect 15160 18380 15853 18408
rect 15160 18368 15166 18380
rect 15841 18377 15853 18380
rect 15887 18377 15899 18411
rect 15841 18371 15899 18377
rect 9214 18300 9220 18352
rect 9272 18340 9278 18352
rect 12437 18343 12495 18349
rect 12437 18340 12449 18343
rect 9272 18312 12449 18340
rect 9272 18300 9278 18312
rect 12437 18309 12449 18312
rect 12483 18340 12495 18343
rect 13538 18340 13544 18352
rect 12483 18312 13544 18340
rect 12483 18309 12495 18312
rect 12437 18303 12495 18309
rect 13538 18300 13544 18312
rect 13596 18300 13602 18352
rect 15286 18340 15292 18352
rect 15247 18312 15292 18340
rect 15286 18300 15292 18312
rect 15344 18300 15350 18352
rect 1903 18244 2452 18272
rect 4709 18275 4767 18281
rect 1903 18241 1915 18244
rect 1857 18235 1915 18241
rect 4709 18241 4721 18275
rect 4755 18272 4767 18275
rect 10226 18272 10232 18284
rect 4755 18244 10232 18272
rect 4755 18241 4767 18244
rect 4709 18235 4767 18241
rect 10226 18232 10232 18244
rect 10284 18232 10290 18284
rect 13081 18275 13139 18281
rect 13081 18272 13093 18275
rect 12406 18244 13093 18272
rect 5442 18164 5448 18216
rect 5500 18204 5506 18216
rect 11793 18207 11851 18213
rect 11793 18204 11805 18207
rect 5500 18176 11805 18204
rect 5500 18164 5506 18176
rect 11793 18173 11805 18176
rect 11839 18204 11851 18207
rect 12406 18204 12434 18244
rect 13081 18241 13093 18244
rect 13127 18241 13139 18275
rect 13722 18272 13728 18284
rect 13683 18244 13728 18272
rect 13081 18235 13139 18241
rect 11839 18176 12434 18204
rect 13096 18204 13124 18235
rect 13722 18232 13728 18244
rect 13780 18232 13786 18284
rect 14645 18275 14703 18281
rect 14645 18241 14657 18275
rect 14691 18272 14703 18275
rect 15304 18272 15332 18300
rect 14691 18244 15332 18272
rect 14691 18241 14703 18244
rect 14645 18235 14703 18241
rect 13906 18204 13912 18216
rect 13096 18176 13912 18204
rect 11839 18173 11851 18176
rect 11793 18167 11851 18173
rect 13906 18164 13912 18176
rect 13964 18164 13970 18216
rect 1670 18068 1676 18080
rect 1631 18040 1676 18068
rect 1670 18028 1676 18040
rect 1728 18028 1734 18080
rect 3326 18028 3332 18080
rect 3384 18068 3390 18080
rect 4617 18071 4675 18077
rect 4617 18068 4629 18071
rect 3384 18040 4629 18068
rect 3384 18028 3390 18040
rect 4617 18037 4629 18040
rect 4663 18037 4675 18071
rect 4617 18031 4675 18037
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 12986 17864 12992 17876
rect 12947 17836 12992 17864
rect 12986 17824 12992 17836
rect 13044 17824 13050 17876
rect 15194 17824 15200 17876
rect 15252 17864 15258 17876
rect 15473 17867 15531 17873
rect 15473 17864 15485 17867
rect 15252 17836 15485 17864
rect 15252 17824 15258 17836
rect 15473 17833 15485 17836
rect 15519 17833 15531 17867
rect 15473 17827 15531 17833
rect 14826 17728 14832 17740
rect 14787 17700 14832 17728
rect 14826 17688 14832 17700
rect 14884 17688 14890 17740
rect 30285 17663 30343 17669
rect 30285 17629 30297 17663
rect 30331 17660 30343 17663
rect 38010 17660 38016 17672
rect 30331 17632 38016 17660
rect 30331 17629 30343 17632
rect 30285 17623 30343 17629
rect 38010 17620 38016 17632
rect 38068 17620 38074 17672
rect 13725 17595 13783 17601
rect 13725 17561 13737 17595
rect 13771 17592 13783 17595
rect 14369 17595 14427 17601
rect 14369 17592 14381 17595
rect 13771 17564 14381 17592
rect 13771 17561 13783 17564
rect 13725 17555 13783 17561
rect 14369 17561 14381 17564
rect 14415 17561 14427 17595
rect 14369 17555 14427 17561
rect 14461 17595 14519 17601
rect 14461 17561 14473 17595
rect 14507 17592 14519 17595
rect 14550 17592 14556 17604
rect 14507 17564 14556 17592
rect 14507 17561 14519 17564
rect 14461 17555 14519 17561
rect 14550 17552 14556 17564
rect 14608 17552 14614 17604
rect 16482 17484 16488 17536
rect 16540 17524 16546 17536
rect 30193 17527 30251 17533
rect 30193 17524 30205 17527
rect 16540 17496 30205 17524
rect 16540 17484 16546 17496
rect 30193 17493 30205 17496
rect 30239 17493 30251 17527
rect 30193 17487 30251 17493
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 13906 17320 13912 17332
rect 13867 17292 13912 17320
rect 13906 17280 13912 17292
rect 13964 17280 13970 17332
rect 14550 17320 14556 17332
rect 14511 17292 14556 17320
rect 14550 17280 14556 17292
rect 14608 17280 14614 17332
rect 15197 17323 15255 17329
rect 15197 17289 15209 17323
rect 15243 17320 15255 17323
rect 15286 17320 15292 17332
rect 15243 17292 15292 17320
rect 15243 17289 15255 17292
rect 15197 17283 15255 17289
rect 15286 17280 15292 17292
rect 15344 17280 15350 17332
rect 13924 17184 13952 17280
rect 14645 17187 14703 17193
rect 14645 17184 14657 17187
rect 13924 17156 14657 17184
rect 14645 17153 14657 17156
rect 14691 17153 14703 17187
rect 14645 17147 14703 17153
rect 15010 17144 15016 17196
rect 15068 17184 15074 17196
rect 25041 17187 25099 17193
rect 25041 17184 25053 17187
rect 15068 17156 25053 17184
rect 15068 17144 15074 17156
rect 25041 17153 25053 17156
rect 25087 17184 25099 17187
rect 25685 17187 25743 17193
rect 25685 17184 25697 17187
rect 25087 17156 25697 17184
rect 25087 17153 25099 17156
rect 25041 17147 25099 17153
rect 25685 17153 25697 17156
rect 25731 17153 25743 17187
rect 25685 17147 25743 17153
rect 25777 16983 25835 16989
rect 25777 16949 25789 16983
rect 25823 16980 25835 16983
rect 34790 16980 34796 16992
rect 25823 16952 34796 16980
rect 25823 16949 25835 16952
rect 25777 16943 25835 16949
rect 34790 16940 34796 16952
rect 34848 16940 34854 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 21821 16643 21879 16649
rect 21821 16640 21833 16643
rect 21284 16612 21833 16640
rect 18598 16532 18604 16584
rect 18656 16572 18662 16584
rect 21284 16581 21312 16612
rect 21821 16609 21833 16612
rect 21867 16640 21879 16643
rect 24578 16640 24584 16652
rect 21867 16612 24584 16640
rect 21867 16609 21879 16612
rect 21821 16603 21879 16609
rect 24578 16600 24584 16612
rect 24636 16600 24642 16652
rect 21177 16575 21235 16581
rect 21177 16572 21189 16575
rect 18656 16544 21189 16572
rect 18656 16532 18662 16544
rect 21177 16541 21189 16544
rect 21223 16541 21235 16575
rect 21177 16535 21235 16541
rect 21269 16575 21327 16581
rect 21269 16541 21281 16575
rect 21315 16574 21327 16575
rect 21315 16546 21349 16574
rect 21315 16541 21327 16546
rect 21269 16535 21327 16541
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 1857 16099 1915 16105
rect 1857 16065 1869 16099
rect 1903 16096 1915 16099
rect 3970 16096 3976 16108
rect 1903 16068 3976 16096
rect 1903 16065 1915 16068
rect 1857 16059 1915 16065
rect 3970 16056 3976 16068
rect 4028 16056 4034 16108
rect 38013 16099 38071 16105
rect 38013 16065 38025 16099
rect 38059 16096 38071 16099
rect 38102 16096 38108 16108
rect 38059 16068 38108 16096
rect 38059 16065 38071 16068
rect 38013 16059 38071 16065
rect 38102 16056 38108 16068
rect 38160 16056 38166 16108
rect 1670 15892 1676 15904
rect 1631 15864 1676 15892
rect 1670 15852 1676 15864
rect 1728 15852 1734 15904
rect 38194 15892 38200 15904
rect 38155 15864 38200 15892
rect 38194 15852 38200 15864
rect 38252 15852 38258 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 38010 14464 38016 14476
rect 37971 14436 38016 14464
rect 38010 14424 38016 14436
rect 38068 14424 38074 14476
rect 38286 14396 38292 14408
rect 38247 14368 38292 14396
rect 38286 14356 38292 14368
rect 38344 14356 38350 14408
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 38286 14056 38292 14068
rect 38247 14028 38292 14056
rect 38286 14016 38292 14028
rect 38344 14016 38350 14068
rect 1857 13923 1915 13929
rect 1857 13889 1869 13923
rect 1903 13920 1915 13923
rect 5258 13920 5264 13932
rect 1903 13892 5264 13920
rect 1903 13889 1915 13892
rect 1857 13883 1915 13889
rect 5258 13880 5264 13892
rect 5316 13880 5322 13932
rect 1670 13716 1676 13728
rect 1631 13688 1676 13716
rect 1670 13676 1676 13688
rect 1728 13676 1734 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 13262 13512 13268 13524
rect 13223 13484 13268 13512
rect 13262 13472 13268 13484
rect 13320 13472 13326 13524
rect 20438 13512 20444 13524
rect 20399 13484 20444 13512
rect 20438 13472 20444 13484
rect 20496 13472 20502 13524
rect 13357 13311 13415 13317
rect 13357 13277 13369 13311
rect 13403 13308 13415 13311
rect 13446 13308 13452 13320
rect 13403 13280 13452 13308
rect 13403 13277 13415 13280
rect 13357 13271 13415 13277
rect 13446 13268 13452 13280
rect 13504 13268 13510 13320
rect 19705 13311 19763 13317
rect 19705 13277 19717 13311
rect 19751 13308 19763 13311
rect 20438 13308 20444 13320
rect 19751 13280 20444 13308
rect 19751 13277 19763 13280
rect 19705 13271 19763 13277
rect 20438 13268 20444 13280
rect 20496 13268 20502 13320
rect 19889 13175 19947 13181
rect 19889 13141 19901 13175
rect 19935 13172 19947 13175
rect 20070 13172 20076 13184
rect 19935 13144 20076 13172
rect 19935 13141 19947 13144
rect 19889 13135 19947 13141
rect 20070 13132 20076 13144
rect 20128 13132 20134 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 16945 12971 17003 12977
rect 16945 12968 16957 12971
rect 16546 12940 16957 12968
rect 1857 12835 1915 12841
rect 1857 12801 1869 12835
rect 1903 12832 1915 12835
rect 3326 12832 3332 12844
rect 1903 12804 3332 12832
rect 1903 12801 1915 12804
rect 1857 12795 1915 12801
rect 3326 12792 3332 12804
rect 3384 12792 3390 12844
rect 16301 12835 16359 12841
rect 16301 12801 16313 12835
rect 16347 12832 16359 12835
rect 16546 12832 16574 12940
rect 16945 12937 16957 12940
rect 16991 12968 17003 12971
rect 21818 12968 21824 12980
rect 16991 12940 21824 12968
rect 16991 12937 17003 12940
rect 16945 12931 17003 12937
rect 21818 12928 21824 12940
rect 21876 12928 21882 12980
rect 16347 12804 16574 12832
rect 38013 12835 38071 12841
rect 16347 12801 16359 12804
rect 16301 12795 16359 12801
rect 38013 12801 38025 12835
rect 38059 12801 38071 12835
rect 38013 12795 38071 12801
rect 37458 12764 37464 12776
rect 37419 12736 37464 12764
rect 37458 12724 37464 12736
rect 37516 12764 37522 12776
rect 38028 12764 38056 12795
rect 37516 12736 38056 12764
rect 37516 12724 37522 12736
rect 1670 12628 1676 12640
rect 1631 12600 1676 12628
rect 1670 12588 1676 12600
rect 1728 12588 1734 12640
rect 16114 12628 16120 12640
rect 16075 12600 16120 12628
rect 16114 12588 16120 12600
rect 16172 12588 16178 12640
rect 38194 12628 38200 12640
rect 38155 12600 38200 12628
rect 38194 12588 38200 12600
rect 38252 12588 38258 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 15657 12359 15715 12365
rect 15657 12325 15669 12359
rect 15703 12356 15715 12359
rect 16850 12356 16856 12368
rect 15703 12328 16856 12356
rect 15703 12325 15715 12328
rect 15657 12319 15715 12325
rect 16850 12316 16856 12328
rect 16908 12316 16914 12368
rect 15473 12223 15531 12229
rect 15473 12189 15485 12223
rect 15519 12220 15531 12223
rect 15562 12220 15568 12232
rect 15519 12192 15568 12220
rect 15519 12189 15531 12192
rect 15473 12183 15531 12189
rect 15562 12180 15568 12192
rect 15620 12220 15626 12232
rect 16117 12223 16175 12229
rect 16117 12220 16129 12223
rect 15620 12192 16129 12220
rect 15620 12180 15626 12192
rect 16117 12189 16129 12192
rect 16163 12189 16175 12223
rect 16117 12183 16175 12189
rect 37829 12223 37887 12229
rect 37829 12189 37841 12223
rect 37875 12220 37887 12223
rect 38010 12220 38016 12232
rect 37875 12192 38016 12220
rect 37875 12189 37887 12192
rect 37829 12183 37887 12189
rect 38010 12180 38016 12192
rect 38068 12180 38074 12232
rect 38010 12084 38016 12096
rect 37971 12056 38016 12084
rect 38010 12044 38016 12056
rect 38068 12044 38074 12096
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 18782 11840 18788 11892
rect 18840 11880 18846 11892
rect 24397 11883 24455 11889
rect 24397 11880 24409 11883
rect 18840 11852 24409 11880
rect 18840 11840 18846 11852
rect 24397 11849 24409 11852
rect 24443 11849 24455 11883
rect 24397 11843 24455 11849
rect 24489 11747 24547 11753
rect 24489 11713 24501 11747
rect 24535 11744 24547 11747
rect 24946 11744 24952 11756
rect 24535 11716 24952 11744
rect 24535 11713 24547 11716
rect 24489 11707 24547 11713
rect 24946 11704 24952 11716
rect 25004 11704 25010 11756
rect 24946 11540 24952 11552
rect 24907 11512 24952 11540
rect 24946 11500 24952 11512
rect 25004 11500 25010 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 37553 11135 37611 11141
rect 37553 11101 37565 11135
rect 37599 11132 37611 11135
rect 37599 11104 38240 11132
rect 37599 11101 37611 11104
rect 37553 11095 37611 11101
rect 38212 11076 38240 11104
rect 38013 11067 38071 11073
rect 38013 11033 38025 11067
rect 38059 11064 38071 11067
rect 38102 11064 38108 11076
rect 38059 11036 38108 11064
rect 38059 11033 38071 11036
rect 38013 11027 38071 11033
rect 38102 11024 38108 11036
rect 38160 11024 38166 11076
rect 38194 11024 38200 11076
rect 38252 11064 38258 11076
rect 38252 11036 38297 11064
rect 38252 11024 38258 11036
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 13078 10752 13084 10804
rect 13136 10792 13142 10804
rect 13173 10795 13231 10801
rect 13173 10792 13185 10795
rect 13136 10764 13185 10792
rect 13136 10752 13142 10764
rect 13173 10761 13185 10764
rect 13219 10761 13231 10795
rect 13173 10755 13231 10761
rect 2409 10727 2467 10733
rect 2409 10724 2421 10727
rect 1872 10696 2421 10724
rect 1872 10665 1900 10696
rect 2409 10693 2421 10696
rect 2455 10724 2467 10727
rect 18506 10724 18512 10736
rect 2455 10696 18512 10724
rect 2455 10693 2467 10696
rect 2409 10687 2467 10693
rect 18506 10684 18512 10696
rect 18564 10684 18570 10736
rect 1857 10659 1915 10665
rect 1857 10625 1869 10659
rect 1903 10625 1915 10659
rect 1857 10619 1915 10625
rect 13265 10659 13323 10665
rect 13265 10625 13277 10659
rect 13311 10656 13323 10659
rect 13311 10628 13860 10656
rect 13311 10625 13323 10628
rect 13265 10619 13323 10625
rect 13832 10464 13860 10628
rect 1670 10452 1676 10464
rect 1631 10424 1676 10452
rect 1670 10412 1676 10424
rect 1728 10412 1734 10464
rect 13814 10452 13820 10464
rect 13775 10424 13820 10452
rect 13814 10412 13820 10424
rect 13872 10412 13878 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 9861 10251 9919 10257
rect 9861 10217 9873 10251
rect 9907 10248 9919 10251
rect 10042 10248 10048 10260
rect 9907 10220 10048 10248
rect 9907 10217 9919 10220
rect 9861 10211 9919 10217
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 12710 10248 12716 10260
rect 12671 10220 12716 10248
rect 12710 10208 12716 10220
rect 12768 10208 12774 10260
rect 8570 10004 8576 10056
rect 8628 10044 8634 10056
rect 9769 10047 9827 10053
rect 9769 10044 9781 10047
rect 8628 10016 9781 10044
rect 8628 10004 8634 10016
rect 9769 10013 9781 10016
rect 9815 10013 9827 10047
rect 9769 10007 9827 10013
rect 12710 10004 12716 10056
rect 12768 10044 12774 10056
rect 13449 10047 13507 10053
rect 13449 10044 13461 10047
rect 12768 10016 13461 10044
rect 12768 10004 12774 10016
rect 13449 10013 13461 10016
rect 13495 10013 13507 10047
rect 13449 10007 13507 10013
rect 13262 9908 13268 9920
rect 13223 9880 13268 9908
rect 13262 9868 13268 9880
rect 13320 9868 13326 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 13814 9664 13820 9716
rect 13872 9704 13878 9716
rect 19978 9704 19984 9716
rect 13872 9676 19984 9704
rect 13872 9664 13878 9676
rect 19978 9664 19984 9676
rect 20036 9664 20042 9716
rect 20254 9596 20260 9648
rect 20312 9636 20318 9648
rect 20717 9639 20775 9645
rect 20717 9636 20729 9639
rect 20312 9608 20729 9636
rect 20312 9596 20318 9608
rect 20717 9605 20729 9608
rect 20763 9636 20775 9639
rect 20763 9608 21312 9636
rect 20763 9605 20775 9608
rect 20717 9599 20775 9605
rect 21284 9577 21312 9608
rect 21269 9571 21327 9577
rect 21269 9537 21281 9571
rect 21315 9537 21327 9571
rect 21269 9531 21327 9537
rect 21361 9367 21419 9373
rect 21361 9333 21373 9367
rect 21407 9364 21419 9367
rect 24762 9364 24768 9376
rect 21407 9336 24768 9364
rect 21407 9333 21419 9336
rect 21361 9327 21419 9333
rect 24762 9324 24768 9336
rect 24820 9324 24826 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 38010 8956 38016 8968
rect 37971 8928 38016 8956
rect 38010 8916 38016 8928
rect 38068 8916 38074 8968
rect 1670 8888 1676 8900
rect 1631 8860 1676 8888
rect 1670 8848 1676 8860
rect 1728 8848 1734 8900
rect 1765 8823 1823 8829
rect 1765 8789 1777 8823
rect 1811 8820 1823 8823
rect 17678 8820 17684 8832
rect 1811 8792 17684 8820
rect 1811 8789 1823 8792
rect 1765 8783 1823 8789
rect 17678 8780 17684 8792
rect 17736 8780 17742 8832
rect 38194 8820 38200 8832
rect 38155 8792 38200 8820
rect 38194 8780 38200 8792
rect 38252 8780 38258 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 1670 8616 1676 8628
rect 1631 8588 1676 8616
rect 1670 8576 1676 8588
rect 1728 8576 1734 8628
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 1857 7463 1915 7469
rect 1857 7429 1869 7463
rect 1903 7460 1915 7463
rect 4798 7460 4804 7472
rect 1903 7432 4804 7460
rect 1903 7429 1915 7432
rect 1857 7423 1915 7429
rect 4798 7420 4804 7432
rect 4856 7420 4862 7472
rect 37734 7420 37740 7472
rect 37792 7460 37798 7472
rect 38013 7463 38071 7469
rect 38013 7460 38025 7463
rect 37792 7432 38025 7460
rect 37792 7420 37798 7432
rect 38013 7429 38025 7432
rect 38059 7429 38071 7463
rect 38013 7423 38071 7429
rect 1578 7352 1584 7404
rect 1636 7392 1642 7404
rect 1673 7395 1731 7401
rect 1673 7392 1685 7395
rect 1636 7364 1685 7392
rect 1636 7352 1642 7364
rect 1673 7361 1685 7364
rect 1719 7361 1731 7395
rect 1673 7355 1731 7361
rect 37553 7395 37611 7401
rect 37553 7361 37565 7395
rect 37599 7392 37611 7395
rect 38194 7392 38200 7404
rect 37599 7364 38200 7392
rect 37599 7361 37611 7364
rect 37553 7355 37611 7361
rect 38194 7352 38200 7364
rect 38252 7352 38258 7404
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 1578 6984 1584 6996
rect 1539 6956 1584 6984
rect 1578 6944 1584 6956
rect 1636 6944 1642 6996
rect 7285 6851 7343 6857
rect 7285 6848 7297 6851
rect 6886 6820 7297 6848
rect 6733 6783 6791 6789
rect 6733 6749 6745 6783
rect 6779 6780 6791 6783
rect 6886 6780 6914 6820
rect 7285 6817 7297 6820
rect 7331 6848 7343 6851
rect 9674 6848 9680 6860
rect 7331 6820 9680 6848
rect 7331 6817 7343 6820
rect 7285 6811 7343 6817
rect 9674 6808 9680 6820
rect 9732 6808 9738 6860
rect 6779 6752 6914 6780
rect 23661 6783 23719 6789
rect 6779 6749 6791 6752
rect 6733 6743 6791 6749
rect 23661 6749 23673 6783
rect 23707 6780 23719 6783
rect 24670 6780 24676 6792
rect 23707 6752 24676 6780
rect 23707 6749 23719 6752
rect 23661 6743 23719 6749
rect 24670 6740 24676 6752
rect 24728 6740 24734 6792
rect 25222 6712 25228 6724
rect 23860 6684 25228 6712
rect 2774 6604 2780 6656
rect 2832 6644 2838 6656
rect 23860 6653 23888 6684
rect 25222 6672 25228 6684
rect 25280 6672 25286 6724
rect 6641 6647 6699 6653
rect 6641 6644 6653 6647
rect 2832 6616 6653 6644
rect 2832 6604 2838 6616
rect 6641 6613 6653 6616
rect 6687 6613 6699 6647
rect 6641 6607 6699 6613
rect 23845 6647 23903 6653
rect 23845 6613 23857 6647
rect 23891 6613 23903 6647
rect 24670 6644 24676 6656
rect 24583 6616 24676 6644
rect 23845 6607 23903 6613
rect 24670 6604 24676 6616
rect 24728 6644 24734 6656
rect 38102 6644 38108 6656
rect 24728 6616 38108 6644
rect 24728 6604 24734 6616
rect 38102 6604 38108 6616
rect 38160 6604 38166 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 32950 6440 32956 6452
rect 32911 6412 32956 6440
rect 32950 6400 32956 6412
rect 33008 6400 33014 6452
rect 32309 6307 32367 6313
rect 32309 6273 32321 6307
rect 32355 6304 32367 6307
rect 32968 6304 32996 6400
rect 32355 6276 32996 6304
rect 32355 6273 32367 6276
rect 32309 6267 32367 6273
rect 32401 6171 32459 6177
rect 32401 6137 32413 6171
rect 32447 6168 32459 6171
rect 34514 6168 34520 6180
rect 32447 6140 34520 6168
rect 32447 6137 32459 6140
rect 32401 6131 32459 6137
rect 34514 6128 34520 6140
rect 34572 6128 34578 6180
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 37918 5788 37924 5840
rect 37976 5828 37982 5840
rect 38013 5831 38071 5837
rect 38013 5828 38025 5831
rect 37976 5800 38025 5828
rect 37976 5788 37982 5800
rect 38013 5797 38025 5800
rect 38059 5797 38071 5831
rect 38013 5791 38071 5797
rect 37553 5627 37611 5633
rect 37553 5593 37565 5627
rect 37599 5624 37611 5627
rect 38194 5624 38200 5636
rect 37599 5596 38200 5624
rect 37599 5593 37611 5596
rect 37553 5587 37611 5593
rect 38194 5584 38200 5596
rect 38252 5584 38258 5636
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 1762 5352 1768 5364
rect 1723 5324 1768 5352
rect 1762 5312 1768 5324
rect 1820 5312 1826 5364
rect 1578 5176 1584 5228
rect 1636 5216 1642 5228
rect 1673 5219 1731 5225
rect 1673 5216 1685 5219
rect 1636 5188 1685 5216
rect 1636 5176 1642 5188
rect 1673 5185 1685 5188
rect 1719 5185 1731 5219
rect 1673 5179 1731 5185
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 1578 4808 1584 4820
rect 1539 4780 1584 4808
rect 1578 4768 1584 4780
rect 1636 4768 1642 4820
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 1857 3519 1915 3525
rect 1857 3485 1869 3519
rect 1903 3516 1915 3519
rect 2774 3516 2780 3528
rect 1903 3488 2780 3516
rect 1903 3485 1915 3488
rect 1857 3479 1915 3485
rect 2774 3476 2780 3488
rect 2832 3476 2838 3528
rect 38013 3519 38071 3525
rect 38013 3516 38025 3519
rect 37476 3488 38025 3516
rect 1946 3408 1952 3460
rect 2004 3448 2010 3460
rect 2409 3451 2467 3457
rect 2409 3448 2421 3451
rect 2004 3420 2421 3448
rect 2004 3408 2010 3420
rect 2409 3417 2421 3420
rect 2455 3448 2467 3451
rect 18690 3448 18696 3460
rect 2455 3420 18696 3448
rect 2455 3417 2467 3420
rect 2409 3411 2467 3417
rect 18690 3408 18696 3420
rect 18748 3408 18754 3460
rect 37476 3392 37504 3488
rect 38013 3485 38025 3488
rect 38059 3485 38071 3519
rect 38013 3479 38071 3485
rect 1670 3380 1676 3392
rect 1631 3352 1676 3380
rect 1670 3340 1676 3352
rect 1728 3340 1734 3392
rect 37458 3380 37464 3392
rect 37419 3352 37464 3380
rect 37458 3340 37464 3352
rect 37516 3340 37522 3392
rect 38194 3380 38200 3392
rect 38155 3352 38200 3380
rect 38194 3340 38200 3352
rect 38252 3340 38258 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 5534 3136 5540 3188
rect 5592 3176 5598 3188
rect 5721 3179 5779 3185
rect 5721 3176 5733 3179
rect 5592 3148 5733 3176
rect 5592 3136 5598 3148
rect 5721 3145 5733 3148
rect 5767 3176 5779 3179
rect 7558 3176 7564 3188
rect 5767 3148 7564 3176
rect 5767 3145 5779 3148
rect 5721 3139 5779 3145
rect 7558 3136 7564 3148
rect 7616 3136 7622 3188
rect 34790 3136 34796 3188
rect 34848 3176 34854 3188
rect 35069 3179 35127 3185
rect 35069 3176 35081 3179
rect 34848 3148 35081 3176
rect 34848 3136 34854 3148
rect 35069 3145 35081 3148
rect 35115 3145 35127 3179
rect 35069 3139 35127 3145
rect 34609 3111 34667 3117
rect 34609 3108 34621 3111
rect 33888 3080 34621 3108
rect 33888 3052 33916 3080
rect 34609 3077 34621 3080
rect 34655 3077 34667 3111
rect 34609 3071 34667 3077
rect 1670 3040 1676 3052
rect 1631 3012 1676 3040
rect 1670 3000 1676 3012
rect 1728 3040 1734 3052
rect 2869 3043 2927 3049
rect 2869 3040 2881 3043
rect 1728 3012 2881 3040
rect 1728 3000 1734 3012
rect 2869 3009 2881 3012
rect 2915 3009 2927 3043
rect 8570 3040 8576 3052
rect 8531 3012 8576 3040
rect 2869 3003 2927 3009
rect 8570 3000 8576 3012
rect 8628 3000 8634 3052
rect 12710 3000 12716 3052
rect 12768 3040 12774 3052
rect 13446 3040 13452 3052
rect 12768 3012 13452 3040
rect 12768 3000 12774 3012
rect 13446 3000 13452 3012
rect 13504 3000 13510 3052
rect 19978 3040 19984 3052
rect 19939 3012 19984 3040
rect 19978 3000 19984 3012
rect 20036 3040 20042 3052
rect 20625 3043 20683 3049
rect 20625 3040 20637 3043
rect 20036 3012 20637 3040
rect 20036 3000 20042 3012
rect 20625 3009 20637 3012
rect 20671 3009 20683 3043
rect 33870 3040 33876 3052
rect 33831 3012 33876 3040
rect 20625 3003 20683 3009
rect 33870 3000 33876 3012
rect 33928 3000 33934 3052
rect 34514 3000 34520 3052
rect 34572 3040 34578 3052
rect 38013 3043 38071 3049
rect 38013 3040 38025 3043
rect 34572 3012 38025 3040
rect 34572 3000 34578 3012
rect 38013 3009 38025 3012
rect 38059 3009 38071 3043
rect 38013 3003 38071 3009
rect 13633 2975 13691 2981
rect 13633 2941 13645 2975
rect 13679 2972 13691 2975
rect 37458 2972 37464 2984
rect 13679 2944 37464 2972
rect 13679 2941 13691 2944
rect 13633 2935 13691 2941
rect 37458 2932 37464 2944
rect 37516 2932 37522 2984
rect 1857 2907 1915 2913
rect 1857 2873 1869 2907
rect 1903 2904 1915 2907
rect 11514 2904 11520 2916
rect 1903 2876 11520 2904
rect 1903 2873 1915 2876
rect 1857 2867 1915 2873
rect 11514 2864 11520 2876
rect 11572 2864 11578 2916
rect 20165 2907 20223 2913
rect 20165 2873 20177 2907
rect 20211 2904 20223 2907
rect 27338 2904 27344 2916
rect 20211 2876 27344 2904
rect 20211 2873 20223 2876
rect 20165 2867 20223 2873
rect 27338 2864 27344 2876
rect 27396 2864 27402 2916
rect 34057 2907 34115 2913
rect 34057 2873 34069 2907
rect 34103 2904 34115 2907
rect 35894 2904 35900 2916
rect 34103 2876 35900 2904
rect 34103 2873 34115 2876
rect 34057 2867 34115 2873
rect 35894 2864 35900 2876
rect 35952 2864 35958 2916
rect 2406 2836 2412 2848
rect 2367 2808 2412 2836
rect 2406 2796 2412 2808
rect 2464 2796 2470 2848
rect 8294 2796 8300 2848
rect 8352 2836 8358 2848
rect 8389 2839 8447 2845
rect 8389 2836 8401 2839
rect 8352 2808 8401 2836
rect 8352 2796 8358 2808
rect 8389 2805 8401 2808
rect 8435 2805 8447 2839
rect 29638 2836 29644 2848
rect 29599 2808 29644 2836
rect 8389 2799 8447 2805
rect 29638 2796 29644 2808
rect 29696 2796 29702 2848
rect 36814 2796 36820 2848
rect 36872 2836 36878 2848
rect 37553 2839 37611 2845
rect 37553 2836 37565 2839
rect 36872 2808 37565 2836
rect 36872 2796 36878 2808
rect 37553 2805 37565 2808
rect 37599 2836 37611 2839
rect 37642 2836 37648 2848
rect 37599 2808 37648 2836
rect 37599 2805 37611 2808
rect 37553 2799 37611 2805
rect 37642 2796 37648 2808
rect 37700 2796 37706 2848
rect 38010 2796 38016 2848
rect 38068 2836 38074 2848
rect 38197 2839 38255 2845
rect 38197 2836 38209 2839
rect 38068 2808 38209 2836
rect 38068 2796 38074 2808
rect 38197 2805 38209 2808
rect 38243 2805 38255 2839
rect 38197 2799 38255 2805
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 11882 2632 11888 2644
rect 11843 2604 11888 2632
rect 11882 2592 11888 2604
rect 11940 2592 11946 2644
rect 14458 2592 14464 2644
rect 14516 2632 14522 2644
rect 14516 2604 15516 2632
rect 14516 2592 14522 2604
rect 2593 2567 2651 2573
rect 2593 2533 2605 2567
rect 2639 2564 2651 2567
rect 15194 2564 15200 2576
rect 2639 2536 8892 2564
rect 15155 2536 15200 2564
rect 2639 2533 2651 2536
rect 2593 2527 2651 2533
rect 4249 2499 4307 2505
rect 4249 2465 4261 2499
rect 4295 2496 4307 2499
rect 8570 2496 8576 2508
rect 4295 2468 8576 2496
rect 4295 2465 4307 2468
rect 4249 2459 4307 2465
rect 8570 2456 8576 2468
rect 8628 2456 8634 2508
rect 8864 2496 8892 2536
rect 15194 2524 15200 2536
rect 15252 2524 15258 2576
rect 15488 2564 15516 2604
rect 16482 2592 16488 2644
rect 16540 2632 16546 2644
rect 18325 2635 18383 2641
rect 18325 2632 18337 2635
rect 16540 2604 18337 2632
rect 16540 2592 16546 2604
rect 18325 2601 18337 2604
rect 18371 2601 18383 2635
rect 32398 2632 32404 2644
rect 32359 2604 32404 2632
rect 18325 2595 18383 2601
rect 32398 2592 32404 2604
rect 32456 2592 32462 2644
rect 33686 2632 33692 2644
rect 33647 2604 33692 2632
rect 33686 2592 33692 2604
rect 33744 2592 33750 2644
rect 36722 2632 36728 2644
rect 36683 2604 36728 2632
rect 36722 2592 36728 2604
rect 36780 2592 36786 2644
rect 37550 2632 37556 2644
rect 37511 2604 37556 2632
rect 37550 2592 37556 2604
rect 37608 2592 37614 2644
rect 21361 2567 21419 2573
rect 21361 2564 21373 2567
rect 15488 2536 21373 2564
rect 21361 2533 21373 2536
rect 21407 2533 21419 2567
rect 23290 2564 23296 2576
rect 23251 2536 23296 2564
rect 21361 2527 21419 2533
rect 19978 2496 19984 2508
rect 8864 2468 19984 2496
rect 19978 2456 19984 2468
rect 20036 2456 20042 2508
rect 1857 2431 1915 2437
rect 1857 2397 1869 2431
rect 1903 2428 1915 2431
rect 1946 2428 1952 2440
rect 1903 2400 1952 2428
rect 1903 2397 1915 2400
rect 1857 2391 1915 2397
rect 1946 2388 1952 2400
rect 2004 2388 2010 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3344 2400 3985 2428
rect 2406 2360 2412 2372
rect 2367 2332 2412 2360
rect 2406 2320 2412 2332
rect 2464 2320 2470 2372
rect 1302 2252 1308 2304
rect 1360 2292 1366 2304
rect 1673 2295 1731 2301
rect 1673 2292 1685 2295
rect 1360 2264 1685 2292
rect 1360 2252 1366 2264
rect 1673 2261 1685 2264
rect 1719 2261 1731 2295
rect 1673 2255 1731 2261
rect 3234 2252 3240 2304
rect 3292 2292 3298 2304
rect 3344 2301 3372 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 5534 2428 5540 2440
rect 5495 2400 5540 2428
rect 3973 2391 4031 2397
rect 5534 2388 5540 2400
rect 5592 2388 5598 2440
rect 6825 2431 6883 2437
rect 6825 2397 6837 2431
rect 6871 2428 6883 2431
rect 8294 2428 8300 2440
rect 6871 2400 7420 2428
rect 8255 2400 8300 2428
rect 6871 2397 6883 2400
rect 6825 2391 6883 2397
rect 7392 2369 7420 2400
rect 8294 2388 8300 2400
rect 8352 2388 8358 2440
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2428 9367 2431
rect 9674 2428 9680 2440
rect 9355 2400 9680 2428
rect 9355 2397 9367 2400
rect 9309 2391 9367 2397
rect 9674 2388 9680 2400
rect 9732 2428 9738 2440
rect 9769 2431 9827 2437
rect 9769 2428 9781 2431
rect 9732 2400 9781 2428
rect 9732 2388 9738 2400
rect 9769 2397 9781 2400
rect 9815 2397 9827 2431
rect 9769 2391 9827 2397
rect 10045 2431 10103 2437
rect 10045 2397 10057 2431
rect 10091 2428 10103 2431
rect 12710 2428 12716 2440
rect 10091 2400 12716 2428
rect 10091 2397 10103 2400
rect 10045 2391 10103 2397
rect 12710 2388 12716 2400
rect 12768 2388 12774 2440
rect 13262 2428 13268 2440
rect 13223 2400 13268 2428
rect 13262 2388 13268 2400
rect 13320 2388 13326 2440
rect 16114 2428 16120 2440
rect 13372 2400 16120 2428
rect 7377 2363 7435 2369
rect 7377 2329 7389 2363
rect 7423 2360 7435 2363
rect 11149 2363 11207 2369
rect 7423 2332 10088 2360
rect 7423 2329 7435 2332
rect 7377 2323 7435 2329
rect 3329 2295 3387 2301
rect 3329 2292 3341 2295
rect 3292 2264 3341 2292
rect 3292 2252 3298 2264
rect 3329 2261 3341 2264
rect 3375 2261 3387 2295
rect 3329 2255 3387 2261
rect 4522 2252 4528 2304
rect 4580 2292 4586 2304
rect 5353 2295 5411 2301
rect 5353 2292 5365 2295
rect 4580 2264 5365 2292
rect 4580 2252 4586 2264
rect 5353 2261 5365 2264
rect 5399 2261 5411 2295
rect 5353 2255 5411 2261
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 6641 2295 6699 2301
rect 6641 2292 6653 2295
rect 6512 2264 6653 2292
rect 6512 2252 6518 2264
rect 6641 2261 6653 2264
rect 6687 2261 6699 2295
rect 6641 2255 6699 2261
rect 8386 2252 8392 2304
rect 8444 2292 8450 2304
rect 8481 2295 8539 2301
rect 8481 2292 8493 2295
rect 8444 2264 8493 2292
rect 8444 2252 8450 2264
rect 8481 2261 8493 2264
rect 8527 2261 8539 2295
rect 10060 2292 10088 2332
rect 11149 2329 11161 2363
rect 11195 2360 11207 2363
rect 11606 2360 11612 2372
rect 11195 2332 11612 2360
rect 11195 2329 11207 2332
rect 11149 2323 11207 2329
rect 11606 2320 11612 2332
rect 11664 2360 11670 2372
rect 11793 2363 11851 2369
rect 11793 2360 11805 2363
rect 11664 2332 11805 2360
rect 11664 2320 11670 2332
rect 11793 2329 11805 2332
rect 11839 2329 11851 2363
rect 13372 2360 13400 2400
rect 16114 2388 16120 2400
rect 16172 2388 16178 2440
rect 16850 2428 16856 2440
rect 16811 2400 16856 2428
rect 16850 2388 16856 2400
rect 16908 2388 16914 2440
rect 20070 2428 20076 2440
rect 20031 2400 20076 2428
rect 20070 2388 20076 2400
rect 20128 2388 20134 2440
rect 21376 2428 21404 2527
rect 23290 2524 23296 2536
rect 23348 2524 23354 2576
rect 24946 2456 24952 2508
rect 25004 2496 25010 2508
rect 30009 2499 30067 2505
rect 30009 2496 30021 2499
rect 25004 2468 30021 2496
rect 25004 2456 25010 2468
rect 30009 2465 30021 2468
rect 30055 2496 30067 2499
rect 33870 2496 33876 2508
rect 30055 2468 33876 2496
rect 30055 2465 30067 2468
rect 30009 2459 30067 2465
rect 33870 2456 33876 2468
rect 33928 2456 33934 2508
rect 22005 2431 22063 2437
rect 22005 2428 22017 2431
rect 21376 2400 22017 2428
rect 22005 2397 22017 2400
rect 22051 2397 22063 2431
rect 25222 2428 25228 2440
rect 25183 2400 25228 2428
rect 22005 2391 22063 2397
rect 25222 2388 25228 2400
rect 25280 2388 25286 2440
rect 27157 2431 27215 2437
rect 27157 2428 27169 2431
rect 26206 2400 27169 2428
rect 11793 2323 11851 2329
rect 11900 2332 13400 2360
rect 14461 2363 14519 2369
rect 11900 2292 11928 2332
rect 14461 2329 14473 2363
rect 14507 2360 14519 2363
rect 14826 2360 14832 2372
rect 14507 2332 14832 2360
rect 14507 2329 14519 2332
rect 14461 2323 14519 2329
rect 14826 2320 14832 2332
rect 14884 2360 14890 2372
rect 15013 2363 15071 2369
rect 15013 2360 15025 2363
rect 14884 2332 15025 2360
rect 14884 2320 14890 2332
rect 15013 2329 15025 2332
rect 15059 2329 15071 2363
rect 15013 2323 15071 2329
rect 17681 2363 17739 2369
rect 17681 2329 17693 2363
rect 17727 2360 17739 2363
rect 18046 2360 18052 2372
rect 17727 2332 18052 2360
rect 17727 2329 17739 2332
rect 17681 2323 17739 2329
rect 18046 2320 18052 2332
rect 18104 2360 18110 2372
rect 18233 2363 18291 2369
rect 18233 2360 18245 2363
rect 18104 2332 18245 2360
rect 18104 2320 18110 2332
rect 18233 2329 18245 2332
rect 18279 2329 18291 2363
rect 18233 2323 18291 2329
rect 22833 2363 22891 2369
rect 22833 2329 22845 2363
rect 22879 2360 22891 2363
rect 23198 2360 23204 2372
rect 22879 2332 23204 2360
rect 22879 2329 22891 2332
rect 22833 2323 22891 2329
rect 23198 2320 23204 2332
rect 23256 2360 23262 2372
rect 23477 2363 23535 2369
rect 23477 2360 23489 2363
rect 23256 2332 23489 2360
rect 23256 2320 23262 2332
rect 23477 2329 23489 2332
rect 23523 2329 23535 2363
rect 23477 2323 23535 2329
rect 24762 2320 24768 2372
rect 24820 2360 24826 2372
rect 26206 2360 26234 2400
rect 27157 2397 27169 2400
rect 27203 2397 27215 2431
rect 27157 2391 27215 2397
rect 27338 2388 27344 2440
rect 27396 2428 27402 2440
rect 28445 2431 28503 2437
rect 28445 2428 28457 2431
rect 27396 2400 28457 2428
rect 27396 2388 27402 2400
rect 28445 2397 28457 2400
rect 28491 2397 28503 2431
rect 28445 2391 28503 2397
rect 29638 2388 29644 2440
rect 29696 2428 29702 2440
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29696 2400 29745 2428
rect 29696 2388 29702 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 34790 2388 34796 2440
rect 34848 2428 34854 2440
rect 35161 2431 35219 2437
rect 35161 2428 35173 2431
rect 34848 2400 35173 2428
rect 34848 2388 34854 2400
rect 35161 2397 35173 2400
rect 35207 2397 35219 2431
rect 35161 2391 35219 2397
rect 35894 2388 35900 2440
rect 35952 2428 35958 2440
rect 35952 2400 35997 2428
rect 35952 2388 35958 2400
rect 37274 2388 37280 2440
rect 37332 2428 37338 2440
rect 37645 2431 37703 2437
rect 37645 2428 37657 2431
rect 37332 2400 37657 2428
rect 37332 2388 37338 2400
rect 37645 2397 37657 2400
rect 37691 2428 37703 2431
rect 38197 2431 38255 2437
rect 38197 2428 38209 2431
rect 37691 2400 38209 2428
rect 37691 2397 37703 2400
rect 37645 2391 37703 2397
rect 38197 2397 38209 2400
rect 38243 2397 38255 2431
rect 38197 2391 38255 2397
rect 32493 2363 32551 2369
rect 32493 2360 32505 2363
rect 24820 2332 26234 2360
rect 31772 2332 32505 2360
rect 24820 2320 24826 2332
rect 31772 2304 31800 2332
rect 32493 2329 32505 2332
rect 32539 2329 32551 2363
rect 32493 2323 32551 2329
rect 33137 2363 33195 2369
rect 33137 2329 33149 2363
rect 33183 2360 33195 2363
rect 33502 2360 33508 2372
rect 33183 2332 33508 2360
rect 33183 2329 33195 2332
rect 33137 2323 33195 2329
rect 33502 2320 33508 2332
rect 33560 2360 33566 2372
rect 33781 2363 33839 2369
rect 33781 2360 33793 2363
rect 33560 2332 33793 2360
rect 33560 2320 33566 2332
rect 33781 2329 33793 2332
rect 33827 2329 33839 2363
rect 36814 2360 36820 2372
rect 36775 2332 36820 2360
rect 33781 2323 33839 2329
rect 36814 2320 36820 2332
rect 36872 2320 36878 2372
rect 10060 2264 11928 2292
rect 8481 2255 8539 2261
rect 12894 2252 12900 2304
rect 12952 2292 12958 2304
rect 13081 2295 13139 2301
rect 13081 2292 13093 2295
rect 12952 2264 13093 2292
rect 12952 2252 12958 2264
rect 13081 2261 13093 2264
rect 13127 2261 13139 2295
rect 13081 2255 13139 2261
rect 16758 2252 16764 2304
rect 16816 2292 16822 2304
rect 17037 2295 17095 2301
rect 17037 2292 17049 2295
rect 16816 2264 17049 2292
rect 16816 2252 16822 2264
rect 17037 2261 17049 2264
rect 17083 2261 17095 2295
rect 17037 2255 17095 2261
rect 19978 2252 19984 2304
rect 20036 2292 20042 2304
rect 20257 2295 20315 2301
rect 20257 2292 20269 2295
rect 20036 2264 20269 2292
rect 20036 2252 20042 2264
rect 20257 2261 20269 2264
rect 20303 2261 20315 2295
rect 20257 2255 20315 2261
rect 21634 2252 21640 2304
rect 21692 2292 21698 2304
rect 22189 2295 22247 2301
rect 22189 2292 22201 2295
rect 21692 2264 22201 2292
rect 21692 2252 21698 2264
rect 22189 2261 22201 2264
rect 22235 2261 22247 2295
rect 22189 2255 22247 2261
rect 25130 2252 25136 2304
rect 25188 2292 25194 2304
rect 25409 2295 25467 2301
rect 25409 2292 25421 2295
rect 25188 2264 25421 2292
rect 25188 2252 25194 2264
rect 25409 2261 25421 2264
rect 25455 2261 25467 2295
rect 25409 2255 25467 2261
rect 26418 2252 26424 2304
rect 26476 2292 26482 2304
rect 27341 2295 27399 2301
rect 27341 2292 27353 2295
rect 26476 2264 27353 2292
rect 26476 2252 26482 2264
rect 27341 2261 27353 2264
rect 27387 2261 27399 2295
rect 27341 2255 27399 2261
rect 28350 2252 28356 2304
rect 28408 2292 28414 2304
rect 28629 2295 28687 2301
rect 28629 2292 28641 2295
rect 28408 2264 28641 2292
rect 28408 2252 28414 2264
rect 28629 2261 28641 2264
rect 28675 2261 28687 2295
rect 31754 2292 31760 2304
rect 31715 2264 31760 2292
rect 28629 2255 28687 2261
rect 31754 2252 31760 2264
rect 31812 2252 31818 2304
rect 34790 2252 34796 2304
rect 34848 2292 34854 2304
rect 34977 2295 35035 2301
rect 34977 2292 34989 2295
rect 34848 2264 34989 2292
rect 34848 2252 34854 2264
rect 34977 2261 34989 2264
rect 35023 2261 35035 2295
rect 34977 2255 35035 2261
rect 35802 2252 35808 2304
rect 35860 2292 35866 2304
rect 36081 2295 36139 2301
rect 36081 2292 36093 2295
rect 35860 2264 36093 2292
rect 35860 2252 35866 2264
rect 36081 2261 36093 2264
rect 36127 2261 36139 2295
rect 36081 2255 36139 2261
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 14 1300 20 1352
rect 72 1340 78 1352
rect 2406 1340 2412 1352
rect 72 1312 2412 1340
rect 72 1300 78 1312
rect 2406 1300 2412 1312
rect 2464 1300 2470 1352
<< via1 >>
rect 4804 37748 4856 37800
rect 16672 37748 16724 37800
rect 10600 37680 10652 37732
rect 22744 37680 22796 37732
rect 20 37612 72 37664
rect 4896 37612 4948 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 3148 37315 3200 37324
rect 3148 37281 3157 37315
rect 3157 37281 3191 37315
rect 3191 37281 3200 37315
rect 3148 37272 3200 37281
rect 3884 37272 3936 37324
rect 4804 37272 4856 37324
rect 10232 37408 10284 37460
rect 10600 37408 10652 37460
rect 9864 37272 9916 37324
rect 10968 37272 11020 37324
rect 2044 37204 2096 37256
rect 5540 37204 5592 37256
rect 8944 37204 8996 37256
rect 11520 37204 11572 37256
rect 12624 37272 12676 37324
rect 20536 37408 20588 37460
rect 22744 37451 22796 37460
rect 22744 37417 22753 37451
rect 22753 37417 22787 37451
rect 22787 37417 22796 37451
rect 22744 37408 22796 37417
rect 23848 37408 23900 37460
rect 36728 37451 36780 37460
rect 36728 37417 36737 37451
rect 36737 37417 36771 37451
rect 36771 37417 36780 37451
rect 36728 37408 36780 37417
rect 13820 37272 13872 37324
rect 16856 37315 16908 37324
rect 16856 37281 16865 37315
rect 16865 37281 16899 37315
rect 16899 37281 16908 37315
rect 16856 37272 16908 37281
rect 18604 37272 18656 37324
rect 32404 37340 32456 37392
rect 30288 37272 30340 37324
rect 5724 37136 5776 37188
rect 5816 37068 5868 37120
rect 6736 37068 6788 37120
rect 6828 37111 6880 37120
rect 6828 37077 6837 37111
rect 6837 37077 6871 37111
rect 6871 37077 6880 37111
rect 7840 37136 7892 37188
rect 6828 37068 6880 37077
rect 9128 37111 9180 37120
rect 9128 37077 9137 37111
rect 9137 37077 9171 37111
rect 9171 37077 9180 37111
rect 10692 37136 10744 37188
rect 13728 37204 13780 37256
rect 15844 37247 15896 37256
rect 11704 37136 11756 37188
rect 14648 37136 14700 37188
rect 15844 37213 15853 37247
rect 15853 37213 15887 37247
rect 15887 37213 15896 37247
rect 15844 37204 15896 37213
rect 16764 37204 16816 37256
rect 19432 37247 19484 37256
rect 19432 37213 19441 37247
rect 19441 37213 19475 37247
rect 19475 37213 19484 37247
rect 19432 37204 19484 37213
rect 20720 37204 20772 37256
rect 21456 37204 21508 37256
rect 23848 37204 23900 37256
rect 19984 37136 20036 37188
rect 23204 37136 23256 37188
rect 28908 37247 28960 37256
rect 28908 37213 28917 37247
rect 28917 37213 28951 37247
rect 28951 37213 28960 37247
rect 28908 37204 28960 37213
rect 30656 37247 30708 37256
rect 30656 37213 30665 37247
rect 30665 37213 30699 37247
rect 30699 37213 30708 37247
rect 30656 37204 30708 37213
rect 33600 37247 33652 37256
rect 33600 37213 33609 37247
rect 33609 37213 33643 37247
rect 33643 37213 33652 37247
rect 33600 37204 33652 37213
rect 35532 37247 35584 37256
rect 35532 37213 35541 37247
rect 35541 37213 35575 37247
rect 35575 37213 35584 37247
rect 35532 37204 35584 37213
rect 37372 37204 37424 37256
rect 31852 37136 31904 37188
rect 9128 37068 9180 37077
rect 12900 37068 12952 37120
rect 15200 37068 15252 37120
rect 15476 37068 15528 37120
rect 15752 37068 15804 37120
rect 18512 37068 18564 37120
rect 18788 37068 18840 37120
rect 20720 37111 20772 37120
rect 20720 37077 20729 37111
rect 20729 37077 20763 37111
rect 20763 37077 20772 37111
rect 20720 37068 20772 37077
rect 22100 37068 22152 37120
rect 23296 37111 23348 37120
rect 23296 37077 23305 37111
rect 23305 37077 23339 37111
rect 23339 37077 23348 37111
rect 23296 37068 23348 37077
rect 24676 37111 24728 37120
rect 24676 37077 24685 37111
rect 24685 37077 24719 37111
rect 24719 37077 24728 37111
rect 24676 37068 24728 37077
rect 25136 37068 25188 37120
rect 26516 37111 26568 37120
rect 26516 37077 26525 37111
rect 26525 37077 26559 37111
rect 26559 37077 26568 37111
rect 26516 37068 26568 37077
rect 27068 37068 27120 37120
rect 29000 37068 29052 37120
rect 31760 37111 31812 37120
rect 31760 37077 31769 37111
rect 31769 37077 31803 37111
rect 31803 37077 31812 37111
rect 31760 37068 31812 37077
rect 32220 37068 32272 37120
rect 33508 37068 33560 37120
rect 35440 37068 35492 37120
rect 37464 37068 37516 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 7840 36864 7892 36916
rect 12532 36864 12584 36916
rect 12624 36864 12676 36916
rect 15568 36864 15620 36916
rect 21456 36864 21508 36916
rect 1584 36796 1636 36848
rect 3700 36796 3752 36848
rect 5724 36839 5776 36848
rect 5724 36805 5733 36839
rect 5733 36805 5767 36839
rect 5767 36805 5776 36839
rect 5724 36796 5776 36805
rect 8668 36796 8720 36848
rect 9128 36796 9180 36848
rect 9588 36796 9640 36848
rect 10600 36796 10652 36848
rect 1676 36728 1728 36780
rect 1308 36660 1360 36712
rect 5356 36660 5408 36712
rect 3332 36524 3384 36576
rect 4620 36524 4672 36576
rect 8576 36728 8628 36780
rect 11336 36796 11388 36848
rect 11888 36796 11940 36848
rect 13452 36839 13504 36848
rect 13452 36805 13461 36839
rect 13461 36805 13495 36839
rect 13495 36805 13504 36839
rect 13452 36796 13504 36805
rect 6828 36660 6880 36712
rect 9036 36592 9088 36644
rect 8392 36524 8444 36576
rect 8944 36524 8996 36576
rect 9864 36660 9916 36712
rect 10876 36703 10928 36712
rect 10876 36669 10885 36703
rect 10885 36669 10919 36703
rect 10919 36669 10928 36703
rect 10876 36660 10928 36669
rect 11520 36660 11572 36712
rect 13728 36771 13780 36780
rect 13728 36737 13737 36771
rect 13737 36737 13771 36771
rect 13771 36737 13780 36771
rect 17868 36796 17920 36848
rect 30656 36864 30708 36916
rect 38200 36907 38252 36916
rect 38200 36873 38209 36907
rect 38209 36873 38243 36907
rect 38243 36873 38252 36907
rect 38200 36864 38252 36873
rect 27620 36796 27672 36848
rect 35532 36796 35584 36848
rect 13728 36728 13780 36737
rect 15016 36728 15068 36780
rect 15752 36728 15804 36780
rect 12440 36592 12492 36644
rect 11152 36524 11204 36576
rect 15292 36660 15344 36712
rect 17500 36728 17552 36780
rect 18052 36728 18104 36780
rect 19984 36728 20036 36780
rect 20720 36660 20772 36712
rect 20812 36660 20864 36712
rect 31668 36728 31720 36780
rect 34336 36771 34388 36780
rect 34336 36737 34345 36771
rect 34345 36737 34379 36771
rect 34379 36737 34388 36771
rect 34336 36728 34388 36737
rect 22192 36592 22244 36644
rect 23296 36592 23348 36644
rect 15016 36567 15068 36576
rect 15016 36533 15025 36567
rect 15025 36533 15059 36567
rect 15059 36533 15068 36567
rect 16856 36567 16908 36576
rect 15016 36524 15068 36533
rect 16856 36533 16865 36567
rect 16865 36533 16899 36567
rect 16899 36533 16908 36567
rect 16856 36524 16908 36533
rect 18788 36567 18840 36576
rect 18788 36533 18797 36567
rect 18797 36533 18831 36567
rect 18831 36533 18840 36567
rect 18788 36524 18840 36533
rect 19340 36524 19392 36576
rect 19984 36567 20036 36576
rect 19984 36533 19993 36567
rect 19993 36533 20027 36567
rect 20027 36533 20036 36567
rect 19984 36524 20036 36533
rect 20536 36567 20588 36576
rect 20536 36533 20545 36567
rect 20545 36533 20579 36567
rect 20579 36533 20588 36567
rect 20536 36524 20588 36533
rect 31852 36660 31904 36712
rect 28908 36592 28960 36644
rect 34428 36567 34480 36576
rect 34428 36533 34437 36567
rect 34437 36533 34471 36567
rect 34471 36533 34480 36567
rect 34428 36524 34480 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 4620 36320 4672 36372
rect 11152 36320 11204 36372
rect 10324 36252 10376 36304
rect 12164 36320 12216 36372
rect 12256 36320 12308 36372
rect 13268 36320 13320 36372
rect 22192 36363 22244 36372
rect 22192 36329 22201 36363
rect 22201 36329 22235 36363
rect 22235 36329 22244 36363
rect 22192 36320 22244 36329
rect 23296 36363 23348 36372
rect 23296 36329 23305 36363
rect 23305 36329 23339 36363
rect 23339 36329 23348 36363
rect 23296 36320 23348 36329
rect 38660 36320 38712 36372
rect 1676 36227 1728 36236
rect 1676 36193 1685 36227
rect 1685 36193 1719 36227
rect 1719 36193 1728 36227
rect 1676 36184 1728 36193
rect 3884 36184 3936 36236
rect 4804 36184 4856 36236
rect 8116 36227 8168 36236
rect 8116 36193 8125 36227
rect 8125 36193 8159 36227
rect 8159 36193 8168 36227
rect 8116 36184 8168 36193
rect 8576 36184 8628 36236
rect 12256 36184 12308 36236
rect 12348 36227 12400 36236
rect 12348 36193 12357 36227
rect 12357 36193 12391 36227
rect 12391 36193 12400 36227
rect 15752 36252 15804 36304
rect 15936 36252 15988 36304
rect 19156 36252 19208 36304
rect 19248 36252 19300 36304
rect 24768 36252 24820 36304
rect 12348 36184 12400 36193
rect 13728 36184 13780 36236
rect 19984 36227 20036 36236
rect 19984 36193 19993 36227
rect 19993 36193 20027 36227
rect 20027 36193 20036 36227
rect 19984 36184 20036 36193
rect 8392 36159 8444 36168
rect 8392 36125 8401 36159
rect 8401 36125 8435 36159
rect 8435 36125 8444 36159
rect 8392 36116 8444 36125
rect 8852 36116 8904 36168
rect 10324 36116 10376 36168
rect 14648 36159 14700 36168
rect 2504 36048 2556 36100
rect 3516 36048 3568 36100
rect 8760 36048 8812 36100
rect 9680 36048 9732 36100
rect 11336 36048 11388 36100
rect 1768 35980 1820 36032
rect 4712 35980 4764 36032
rect 12348 36048 12400 36100
rect 12440 36048 12492 36100
rect 13268 36048 13320 36100
rect 14648 36125 14657 36159
rect 14657 36125 14691 36159
rect 14691 36125 14700 36159
rect 14648 36116 14700 36125
rect 15292 36159 15344 36168
rect 15292 36125 15301 36159
rect 15301 36125 15335 36159
rect 15335 36125 15344 36159
rect 15292 36116 15344 36125
rect 15752 36159 15804 36168
rect 15752 36125 15761 36159
rect 15761 36125 15795 36159
rect 15795 36125 15804 36159
rect 15752 36116 15804 36125
rect 16028 36116 16080 36168
rect 16856 36048 16908 36100
rect 18880 36116 18932 36168
rect 34336 36184 34388 36236
rect 34428 36116 34480 36168
rect 12256 35980 12308 36032
rect 14464 35980 14516 36032
rect 14740 35980 14792 36032
rect 14924 35980 14976 36032
rect 15384 35980 15436 36032
rect 16396 36023 16448 36032
rect 16396 35989 16405 36023
rect 16405 35989 16439 36023
rect 16439 35989 16448 36023
rect 16396 35980 16448 35989
rect 17776 35980 17828 36032
rect 18512 36023 18564 36032
rect 18512 35989 18521 36023
rect 18521 35989 18555 36023
rect 18555 35989 18564 36023
rect 18512 35980 18564 35989
rect 19064 35980 19116 36032
rect 19340 36048 19392 36100
rect 23112 36048 23164 36100
rect 20812 35980 20864 36032
rect 21640 36023 21692 36032
rect 21640 35989 21649 36023
rect 21649 35989 21683 36023
rect 21683 35989 21692 36023
rect 21640 35980 21692 35989
rect 24584 36023 24636 36032
rect 24584 35989 24593 36023
rect 24593 35989 24627 36023
rect 24627 35989 24636 36023
rect 24584 35980 24636 35989
rect 25688 36023 25740 36032
rect 25688 35989 25697 36023
rect 25697 35989 25731 36023
rect 25731 35989 25740 36023
rect 25688 35980 25740 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 3516 35776 3568 35828
rect 8024 35776 8076 35828
rect 8484 35776 8536 35828
rect 10600 35776 10652 35828
rect 10692 35776 10744 35828
rect 2872 35708 2924 35760
rect 3792 35708 3844 35760
rect 5448 35708 5500 35760
rect 8208 35708 8260 35760
rect 8668 35751 8720 35760
rect 8668 35717 8677 35751
rect 8677 35717 8711 35751
rect 8711 35717 8720 35751
rect 8668 35708 8720 35717
rect 10784 35708 10836 35760
rect 11336 35776 11388 35828
rect 11520 35776 11572 35828
rect 13176 35751 13228 35760
rect 1952 35640 2004 35692
rect 2780 35640 2832 35692
rect 3976 35640 4028 35692
rect 5356 35683 5408 35692
rect 5356 35649 5365 35683
rect 5365 35649 5399 35683
rect 5399 35649 5408 35683
rect 5356 35640 5408 35649
rect 6644 35640 6696 35692
rect 8944 35683 8996 35692
rect 8944 35649 8953 35683
rect 8953 35649 8987 35683
rect 8987 35649 8996 35683
rect 8944 35640 8996 35649
rect 9772 35640 9824 35692
rect 13176 35717 13185 35751
rect 13185 35717 13219 35751
rect 13219 35717 13228 35751
rect 13176 35708 13228 35717
rect 14464 35776 14516 35828
rect 17960 35776 18012 35828
rect 2872 35615 2924 35624
rect 2872 35581 2881 35615
rect 2881 35581 2915 35615
rect 2915 35581 2924 35615
rect 2872 35572 2924 35581
rect 5080 35572 5132 35624
rect 1860 35547 1912 35556
rect 1860 35513 1869 35547
rect 1869 35513 1903 35547
rect 1903 35513 1912 35547
rect 1860 35504 1912 35513
rect 1952 35504 2004 35556
rect 9312 35572 9364 35624
rect 9404 35572 9456 35624
rect 10508 35572 10560 35624
rect 3608 35479 3660 35488
rect 3608 35445 3617 35479
rect 3617 35445 3651 35479
rect 3651 35445 3660 35479
rect 3608 35436 3660 35445
rect 7472 35504 7524 35556
rect 5632 35436 5684 35488
rect 5908 35479 5960 35488
rect 5908 35445 5917 35479
rect 5917 35445 5951 35479
rect 5951 35445 5960 35479
rect 5908 35436 5960 35445
rect 7196 35436 7248 35488
rect 8208 35436 8260 35488
rect 9864 35504 9916 35556
rect 11336 35572 11388 35624
rect 13728 35640 13780 35692
rect 14188 35640 14240 35692
rect 15200 35708 15252 35760
rect 15292 35640 15344 35692
rect 15476 35683 15528 35692
rect 15476 35649 15485 35683
rect 15485 35649 15519 35683
rect 15519 35649 15528 35683
rect 15476 35640 15528 35649
rect 16028 35640 16080 35692
rect 16948 35708 17000 35760
rect 19984 35776 20036 35828
rect 21088 35776 21140 35828
rect 27620 35776 27672 35828
rect 21640 35708 21692 35760
rect 17776 35683 17828 35692
rect 17776 35649 17785 35683
rect 17785 35649 17819 35683
rect 17819 35649 17828 35683
rect 17776 35640 17828 35649
rect 18420 35640 18472 35692
rect 37464 35640 37516 35692
rect 12716 35572 12768 35624
rect 12808 35572 12860 35624
rect 15660 35572 15712 35624
rect 16120 35572 16172 35624
rect 19524 35572 19576 35624
rect 25320 35615 25372 35624
rect 25320 35581 25329 35615
rect 25329 35581 25363 35615
rect 25363 35581 25372 35615
rect 25320 35572 25372 35581
rect 10876 35436 10928 35488
rect 11612 35436 11664 35488
rect 14004 35504 14056 35556
rect 12808 35436 12860 35488
rect 15476 35436 15528 35488
rect 16120 35436 16172 35488
rect 16488 35436 16540 35488
rect 16948 35479 17000 35488
rect 16948 35445 16957 35479
rect 16957 35445 16991 35479
rect 16991 35445 17000 35479
rect 16948 35436 17000 35445
rect 17776 35436 17828 35488
rect 19248 35436 19300 35488
rect 19524 35479 19576 35488
rect 19524 35445 19533 35479
rect 19533 35445 19567 35479
rect 19567 35445 19576 35479
rect 19524 35436 19576 35445
rect 20168 35436 20220 35488
rect 37464 35479 37516 35488
rect 37464 35445 37473 35479
rect 37473 35445 37507 35479
rect 37507 35445 37516 35479
rect 37464 35436 37516 35445
rect 38200 35479 38252 35488
rect 38200 35445 38209 35479
rect 38209 35445 38243 35479
rect 38243 35445 38252 35479
rect 38200 35436 38252 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 3516 35232 3568 35284
rect 1676 35139 1728 35148
rect 1676 35105 1685 35139
rect 1685 35105 1719 35139
rect 1719 35105 1728 35139
rect 1676 35096 1728 35105
rect 10692 35232 10744 35284
rect 7656 35164 7708 35216
rect 12256 35232 12308 35284
rect 15108 35232 15160 35284
rect 15200 35232 15252 35284
rect 18052 35275 18104 35284
rect 11520 35096 11572 35148
rect 11612 35096 11664 35148
rect 13176 35164 13228 35216
rect 18052 35241 18061 35275
rect 18061 35241 18095 35275
rect 18095 35241 18104 35275
rect 18052 35232 18104 35241
rect 18696 35275 18748 35284
rect 18696 35241 18705 35275
rect 18705 35241 18739 35275
rect 18739 35241 18748 35275
rect 18696 35232 18748 35241
rect 21088 35275 21140 35284
rect 21088 35241 21097 35275
rect 21097 35241 21131 35275
rect 21131 35241 21140 35275
rect 21088 35232 21140 35241
rect 12716 35096 12768 35148
rect 6276 35071 6328 35080
rect 1952 35003 2004 35012
rect 1952 34969 1961 35003
rect 1961 34969 1995 35003
rect 1995 34969 2004 35003
rect 1952 34960 2004 34969
rect 4068 34960 4120 35012
rect 5356 34960 5408 35012
rect 6276 35037 6285 35071
rect 6285 35037 6319 35071
rect 6319 35037 6328 35071
rect 6276 35028 6328 35037
rect 8116 35028 8168 35080
rect 9128 35071 9180 35080
rect 5816 34960 5868 35012
rect 6552 35003 6604 35012
rect 6552 34969 6561 35003
rect 6561 34969 6595 35003
rect 6595 34969 6604 35003
rect 6552 34960 6604 34969
rect 8024 34960 8076 35012
rect 8300 35003 8352 35012
rect 8300 34969 8309 35003
rect 8309 34969 8343 35003
rect 8343 34969 8352 35003
rect 8300 34960 8352 34969
rect 9128 35037 9137 35071
rect 9137 35037 9171 35071
rect 9171 35037 9180 35071
rect 9128 35028 9180 35037
rect 10784 35028 10836 35080
rect 13912 35028 13964 35080
rect 10876 34960 10928 35012
rect 11152 35003 11204 35012
rect 11152 34969 11161 35003
rect 11161 34969 11195 35003
rect 11195 34969 11204 35003
rect 11152 34960 11204 34969
rect 11244 34960 11296 35012
rect 12440 34960 12492 35012
rect 14004 34960 14056 35012
rect 20352 35096 20404 35148
rect 16120 35071 16172 35080
rect 16120 35037 16129 35071
rect 16129 35037 16163 35071
rect 16163 35037 16172 35071
rect 16120 35028 16172 35037
rect 16212 35071 16264 35080
rect 16212 35037 16221 35071
rect 16221 35037 16255 35071
rect 16255 35037 16264 35071
rect 16212 35028 16264 35037
rect 15568 34960 15620 35012
rect 18696 35028 18748 35080
rect 19248 35028 19300 35080
rect 17316 34960 17368 35012
rect 17868 34960 17920 35012
rect 17960 34960 18012 35012
rect 23020 34960 23072 35012
rect 3792 34892 3844 34944
rect 5632 34892 5684 34944
rect 12716 34892 12768 34944
rect 14096 34892 14148 34944
rect 15292 34892 15344 34944
rect 16856 34892 16908 34944
rect 17040 34892 17092 34944
rect 20444 34892 20496 34944
rect 21364 34892 21416 34944
rect 23388 34892 23440 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 12716 34688 12768 34740
rect 12808 34688 12860 34740
rect 18236 34688 18288 34740
rect 19156 34731 19208 34740
rect 19156 34697 19165 34731
rect 19165 34697 19199 34731
rect 19199 34697 19208 34731
rect 19156 34688 19208 34697
rect 21088 34688 21140 34740
rect 22928 34688 22980 34740
rect 23388 34688 23440 34740
rect 1676 34552 1728 34604
rect 3884 34552 3936 34604
rect 5356 34552 5408 34604
rect 7288 34620 7340 34672
rect 6276 34552 6328 34604
rect 8116 34552 8168 34604
rect 7104 34484 7156 34536
rect 9128 34620 9180 34672
rect 12256 34620 12308 34672
rect 12440 34620 12492 34672
rect 15016 34620 15068 34672
rect 17592 34620 17644 34672
rect 10508 34552 10560 34604
rect 11520 34552 11572 34604
rect 15108 34552 15160 34604
rect 15660 34552 15712 34604
rect 18052 34620 18104 34672
rect 23112 34663 23164 34672
rect 17960 34595 18012 34604
rect 17960 34561 17969 34595
rect 17969 34561 18003 34595
rect 18003 34561 18012 34595
rect 23112 34629 23121 34663
rect 23121 34629 23155 34663
rect 23155 34629 23164 34663
rect 23112 34620 23164 34629
rect 17960 34552 18012 34561
rect 18236 34552 18288 34604
rect 19248 34595 19300 34604
rect 19248 34561 19257 34595
rect 19257 34561 19291 34595
rect 19291 34561 19300 34595
rect 19248 34552 19300 34561
rect 20720 34552 20772 34604
rect 20812 34552 20864 34604
rect 8576 34484 8628 34536
rect 8944 34527 8996 34536
rect 8944 34493 8953 34527
rect 8953 34493 8987 34527
rect 8987 34493 8996 34527
rect 8944 34484 8996 34493
rect 9588 34484 9640 34536
rect 9772 34484 9824 34536
rect 9864 34484 9916 34536
rect 3792 34416 3844 34468
rect 6460 34416 6512 34468
rect 5632 34348 5684 34400
rect 6184 34348 6236 34400
rect 7380 34348 7432 34400
rect 8392 34348 8444 34400
rect 10692 34348 10744 34400
rect 12072 34484 12124 34536
rect 12348 34484 12400 34536
rect 13176 34484 13228 34536
rect 14280 34484 14332 34536
rect 14464 34527 14516 34536
rect 14464 34493 14473 34527
rect 14473 34493 14507 34527
rect 14507 34493 14516 34527
rect 14464 34484 14516 34493
rect 15752 34484 15804 34536
rect 16580 34484 16632 34536
rect 17132 34484 17184 34536
rect 19984 34484 20036 34536
rect 20076 34484 20128 34536
rect 19064 34348 19116 34400
rect 19156 34348 19208 34400
rect 21916 34348 21968 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 6644 34144 6696 34196
rect 8208 34144 8260 34196
rect 8300 34144 8352 34196
rect 12256 34144 12308 34196
rect 12348 34144 12400 34196
rect 3516 34008 3568 34060
rect 3884 34008 3936 34060
rect 5724 33940 5776 33992
rect 8944 34008 8996 34060
rect 11428 34076 11480 34128
rect 16212 34144 16264 34196
rect 17224 34144 17276 34196
rect 19064 34144 19116 34196
rect 21088 34144 21140 34196
rect 22928 34187 22980 34196
rect 22928 34153 22937 34187
rect 22937 34153 22971 34187
rect 22971 34153 22980 34187
rect 22928 34144 22980 34153
rect 14372 34076 14424 34128
rect 14464 34076 14516 34128
rect 19156 34076 19208 34128
rect 10692 34008 10744 34060
rect 11612 34051 11664 34060
rect 11612 34017 11621 34051
rect 11621 34017 11655 34051
rect 11655 34017 11664 34051
rect 11612 34008 11664 34017
rect 12256 34008 12308 34060
rect 12532 34008 12584 34060
rect 12624 34008 12676 34060
rect 2136 33872 2188 33924
rect 4252 33915 4304 33924
rect 1584 33804 1636 33856
rect 4252 33881 4261 33915
rect 4261 33881 4295 33915
rect 4295 33881 4304 33915
rect 4252 33872 4304 33881
rect 4988 33872 5040 33924
rect 5816 33872 5868 33924
rect 6460 33872 6512 33924
rect 10784 33940 10836 33992
rect 14556 33940 14608 33992
rect 15660 33940 15712 33992
rect 17040 34008 17092 34060
rect 18604 34008 18656 34060
rect 19892 34008 19944 34060
rect 8484 33872 8536 33924
rect 9128 33872 9180 33924
rect 8576 33804 8628 33856
rect 9036 33804 9088 33856
rect 14464 33915 14516 33924
rect 14464 33881 14473 33915
rect 14473 33881 14507 33915
rect 14507 33881 14516 33915
rect 14464 33872 14516 33881
rect 15384 33915 15436 33924
rect 15384 33881 15393 33915
rect 15393 33881 15427 33915
rect 15427 33881 15436 33915
rect 15384 33872 15436 33881
rect 15936 33872 15988 33924
rect 17316 33940 17368 33992
rect 17960 33940 18012 33992
rect 18052 33940 18104 33992
rect 20168 33940 20220 33992
rect 20628 34008 20680 34060
rect 31668 34008 31720 34060
rect 10784 33804 10836 33856
rect 12716 33804 12768 33856
rect 13268 33804 13320 33856
rect 13452 33804 13504 33856
rect 19064 33804 19116 33856
rect 19524 33804 19576 33856
rect 22008 33872 22060 33924
rect 21824 33847 21876 33856
rect 21824 33813 21833 33847
rect 21833 33813 21867 33847
rect 21867 33813 21876 33847
rect 21824 33804 21876 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 1860 33600 1912 33652
rect 11336 33600 11388 33652
rect 2688 33532 2740 33584
rect 6000 33532 6052 33584
rect 6828 33532 6880 33584
rect 8392 33532 8444 33584
rect 8576 33532 8628 33584
rect 15108 33600 15160 33652
rect 3516 33507 3568 33516
rect 3516 33473 3525 33507
rect 3525 33473 3559 33507
rect 3559 33473 3568 33507
rect 3516 33464 3568 33473
rect 1952 33396 2004 33448
rect 3240 33439 3292 33448
rect 3240 33405 3249 33439
rect 3249 33405 3283 33439
rect 3283 33405 3292 33439
rect 3240 33396 3292 33405
rect 2228 33260 2280 33312
rect 4712 33396 4764 33448
rect 5724 33396 5776 33448
rect 7840 33396 7892 33448
rect 8944 33464 8996 33516
rect 10784 33464 10836 33516
rect 11888 33532 11940 33584
rect 15568 33600 15620 33652
rect 16396 33600 16448 33652
rect 17408 33600 17460 33652
rect 20076 33600 20128 33652
rect 20720 33643 20772 33652
rect 20720 33609 20729 33643
rect 20729 33609 20763 33643
rect 20763 33609 20772 33643
rect 20720 33600 20772 33609
rect 21916 33600 21968 33652
rect 22928 33600 22980 33652
rect 24768 33643 24820 33652
rect 24768 33609 24777 33643
rect 24777 33609 24811 33643
rect 24811 33609 24820 33643
rect 24768 33600 24820 33609
rect 11612 33464 11664 33516
rect 13728 33507 13780 33516
rect 13728 33473 13737 33507
rect 13737 33473 13771 33507
rect 13771 33473 13780 33507
rect 13728 33464 13780 33473
rect 13912 33464 13964 33516
rect 14372 33464 14424 33516
rect 16948 33532 17000 33584
rect 18420 33532 18472 33584
rect 18696 33532 18748 33584
rect 19064 33532 19116 33584
rect 19984 33532 20036 33584
rect 17316 33507 17368 33516
rect 17316 33473 17325 33507
rect 17325 33473 17359 33507
rect 17359 33473 17368 33507
rect 17316 33464 17368 33473
rect 9864 33396 9916 33448
rect 11244 33396 11296 33448
rect 12716 33396 12768 33448
rect 15660 33439 15712 33448
rect 15660 33405 15669 33439
rect 15669 33405 15703 33439
rect 15703 33405 15712 33439
rect 15660 33396 15712 33405
rect 17224 33396 17276 33448
rect 18604 33439 18656 33448
rect 18604 33405 18613 33439
rect 18613 33405 18647 33439
rect 18647 33405 18656 33439
rect 18604 33396 18656 33405
rect 19800 33439 19852 33448
rect 8300 33260 8352 33312
rect 14556 33328 14608 33380
rect 19800 33405 19809 33439
rect 19809 33405 19843 33439
rect 19843 33405 19852 33439
rect 19800 33396 19852 33405
rect 11796 33260 11848 33312
rect 13452 33260 13504 33312
rect 15384 33260 15436 33312
rect 19340 33328 19392 33380
rect 19524 33260 19576 33312
rect 19616 33260 19668 33312
rect 24584 33532 24636 33584
rect 38200 33507 38252 33516
rect 38200 33473 38209 33507
rect 38209 33473 38243 33507
rect 38243 33473 38252 33507
rect 38200 33464 38252 33473
rect 23664 33371 23716 33380
rect 23664 33337 23673 33371
rect 23673 33337 23707 33371
rect 23707 33337 23716 33371
rect 23664 33328 23716 33337
rect 34520 33328 34572 33380
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 1768 33056 1820 33108
rect 7564 33056 7616 33108
rect 8668 33056 8720 33108
rect 9496 33056 9548 33108
rect 10784 32988 10836 33040
rect 12348 33056 12400 33108
rect 13268 32988 13320 33040
rect 3516 32920 3568 32972
rect 9312 32920 9364 32972
rect 11244 32920 11296 32972
rect 11520 32920 11572 32972
rect 4068 32895 4120 32904
rect 4068 32861 4077 32895
rect 4077 32861 4111 32895
rect 4111 32861 4120 32895
rect 4068 32852 4120 32861
rect 4896 32852 4948 32904
rect 5724 32852 5776 32904
rect 7196 32852 7248 32904
rect 7380 32852 7432 32904
rect 8668 32852 8720 32904
rect 9588 32895 9640 32904
rect 9588 32861 9597 32895
rect 9597 32861 9631 32895
rect 9631 32861 9640 32895
rect 9588 32852 9640 32861
rect 2596 32784 2648 32836
rect 4252 32827 4304 32836
rect 4252 32793 4261 32827
rect 4261 32793 4295 32827
rect 4295 32793 4304 32827
rect 4252 32784 4304 32793
rect 6092 32827 6144 32836
rect 6092 32793 6101 32827
rect 6101 32793 6135 32827
rect 6135 32793 6144 32827
rect 6092 32784 6144 32793
rect 8116 32784 8168 32836
rect 9496 32784 9548 32836
rect 12808 32852 12860 32904
rect 15108 33056 15160 33108
rect 18512 33056 18564 33108
rect 19524 33099 19576 33108
rect 19524 33065 19533 33099
rect 19533 33065 19567 33099
rect 19567 33065 19576 33099
rect 19524 33056 19576 33065
rect 20168 33099 20220 33108
rect 20168 33065 20177 33099
rect 20177 33065 20211 33099
rect 20211 33065 20220 33099
rect 20168 33056 20220 33065
rect 22928 33056 22980 33108
rect 13912 32988 13964 33040
rect 15936 33031 15988 33040
rect 15936 32997 15945 33031
rect 15945 32997 15979 33031
rect 15979 32997 15988 33031
rect 15936 32988 15988 32997
rect 17684 32988 17736 33040
rect 18144 32988 18196 33040
rect 19156 32988 19208 33040
rect 20904 32988 20956 33040
rect 13728 32920 13780 32972
rect 14832 32920 14884 32972
rect 16212 32920 16264 32972
rect 16488 32963 16540 32972
rect 16488 32929 16497 32963
rect 16497 32929 16531 32963
rect 16531 32929 16540 32963
rect 16488 32920 16540 32929
rect 17316 32920 17368 32972
rect 21824 32920 21876 32972
rect 15200 32852 15252 32904
rect 17040 32895 17092 32904
rect 17040 32861 17049 32895
rect 17049 32861 17083 32895
rect 17083 32861 17092 32895
rect 17040 32852 17092 32861
rect 17224 32852 17276 32904
rect 18144 32895 18196 32904
rect 18144 32861 18153 32895
rect 18153 32861 18187 32895
rect 18187 32861 18196 32895
rect 18144 32852 18196 32861
rect 18236 32852 18288 32904
rect 19248 32852 19300 32904
rect 10048 32784 10100 32836
rect 12440 32784 12492 32836
rect 13084 32784 13136 32836
rect 17132 32784 17184 32836
rect 17316 32827 17368 32836
rect 17316 32793 17325 32827
rect 17325 32793 17359 32827
rect 17359 32793 17368 32827
rect 17316 32784 17368 32793
rect 18052 32784 18104 32836
rect 19156 32784 19208 32836
rect 20720 32852 20772 32904
rect 20996 32852 21048 32904
rect 21088 32784 21140 32836
rect 4712 32716 4764 32768
rect 9956 32716 10008 32768
rect 11796 32716 11848 32768
rect 11888 32716 11940 32768
rect 13452 32716 13504 32768
rect 13636 32759 13688 32768
rect 13636 32725 13645 32759
rect 13645 32725 13679 32759
rect 13679 32725 13688 32759
rect 13636 32716 13688 32725
rect 14832 32716 14884 32768
rect 17500 32716 17552 32768
rect 19800 32716 19852 32768
rect 23296 32716 23348 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 7288 32512 7340 32564
rect 9496 32512 9548 32564
rect 9588 32512 9640 32564
rect 11152 32512 11204 32564
rect 13636 32512 13688 32564
rect 2688 32444 2740 32496
rect 5908 32444 5960 32496
rect 6000 32487 6052 32496
rect 6000 32453 6009 32487
rect 6009 32453 6043 32487
rect 6043 32453 6052 32487
rect 6000 32444 6052 32453
rect 6552 32444 6604 32496
rect 3516 32419 3568 32428
rect 3516 32385 3525 32419
rect 3525 32385 3559 32419
rect 3559 32385 3568 32419
rect 3516 32376 3568 32385
rect 3792 32376 3844 32428
rect 1768 32215 1820 32224
rect 1768 32181 1777 32215
rect 1777 32181 1811 32215
rect 1811 32181 1820 32215
rect 1768 32172 1820 32181
rect 4804 32308 4856 32360
rect 6552 32351 6604 32360
rect 6552 32317 6561 32351
rect 6561 32317 6595 32351
rect 6595 32317 6604 32351
rect 6552 32308 6604 32317
rect 7012 32444 7064 32496
rect 9680 32444 9732 32496
rect 11520 32444 11572 32496
rect 12624 32444 12676 32496
rect 13176 32487 13228 32496
rect 13176 32453 13185 32487
rect 13185 32453 13219 32487
rect 13219 32453 13228 32487
rect 13176 32444 13228 32453
rect 14096 32487 14148 32496
rect 14096 32453 14105 32487
rect 14105 32453 14139 32487
rect 14139 32453 14148 32487
rect 14096 32444 14148 32453
rect 15476 32487 15528 32496
rect 15476 32453 15485 32487
rect 15485 32453 15519 32487
rect 15519 32453 15528 32487
rect 15476 32444 15528 32453
rect 21640 32512 21692 32564
rect 22928 32512 22980 32564
rect 18420 32487 18472 32496
rect 18420 32453 18429 32487
rect 18429 32453 18463 32487
rect 18463 32453 18472 32487
rect 18420 32444 18472 32453
rect 19248 32444 19300 32496
rect 20720 32444 20772 32496
rect 9312 32419 9364 32428
rect 9312 32385 9321 32419
rect 9321 32385 9355 32419
rect 9355 32385 9364 32419
rect 9312 32376 9364 32385
rect 14648 32419 14700 32428
rect 14648 32385 14657 32419
rect 14657 32385 14691 32419
rect 14691 32385 14700 32419
rect 14648 32376 14700 32385
rect 9128 32308 9180 32360
rect 9588 32351 9640 32360
rect 9588 32317 9597 32351
rect 9597 32317 9631 32351
rect 9631 32317 9640 32351
rect 9588 32308 9640 32317
rect 11244 32308 11296 32360
rect 13728 32308 13780 32360
rect 9312 32240 9364 32292
rect 11888 32240 11940 32292
rect 13544 32240 13596 32292
rect 15476 32308 15528 32360
rect 16672 32308 16724 32360
rect 17408 32376 17460 32428
rect 19156 32376 19208 32428
rect 20904 32376 20956 32428
rect 38200 32419 38252 32428
rect 38200 32385 38209 32419
rect 38209 32385 38243 32419
rect 38243 32385 38252 32419
rect 38200 32376 38252 32385
rect 16304 32240 16356 32292
rect 20076 32308 20128 32360
rect 23572 32240 23624 32292
rect 38016 32283 38068 32292
rect 38016 32249 38025 32283
rect 38025 32249 38059 32283
rect 38059 32249 38068 32283
rect 38016 32240 38068 32249
rect 7288 32172 7340 32224
rect 8668 32172 8720 32224
rect 10968 32172 11020 32224
rect 11152 32172 11204 32224
rect 12624 32172 12676 32224
rect 12992 32172 13044 32224
rect 16948 32172 17000 32224
rect 17316 32172 17368 32224
rect 17408 32172 17460 32224
rect 20168 32172 20220 32224
rect 22468 32172 22520 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 7564 31968 7616 32020
rect 3056 31832 3108 31884
rect 3608 31832 3660 31884
rect 4896 31832 4948 31884
rect 5080 31832 5132 31884
rect 6736 31900 6788 31952
rect 9496 31943 9548 31952
rect 9496 31909 9505 31943
rect 9505 31909 9539 31943
rect 9539 31909 9548 31943
rect 9496 31900 9548 31909
rect 11428 31900 11480 31952
rect 2780 31764 2832 31816
rect 3148 31764 3200 31816
rect 3424 31807 3476 31816
rect 3424 31773 3433 31807
rect 3433 31773 3467 31807
rect 3467 31773 3476 31807
rect 3424 31764 3476 31773
rect 5724 31807 5776 31816
rect 5724 31773 5733 31807
rect 5733 31773 5767 31807
rect 5767 31773 5776 31807
rect 9680 31832 9732 31884
rect 10968 31832 11020 31884
rect 11244 31875 11296 31884
rect 11244 31841 11253 31875
rect 11253 31841 11287 31875
rect 11287 31841 11296 31875
rect 11244 31832 11296 31841
rect 11796 31832 11848 31884
rect 13360 31832 13412 31884
rect 5724 31764 5776 31773
rect 8668 31764 8720 31816
rect 4896 31696 4948 31748
rect 5448 31696 5500 31748
rect 5908 31696 5960 31748
rect 6368 31696 6420 31748
rect 6920 31696 6972 31748
rect 8116 31696 8168 31748
rect 4804 31628 4856 31680
rect 7932 31628 7984 31680
rect 9864 31764 9916 31816
rect 11336 31764 11388 31816
rect 13084 31807 13136 31816
rect 13084 31773 13093 31807
rect 13093 31773 13127 31807
rect 13127 31773 13136 31807
rect 13084 31764 13136 31773
rect 13636 31968 13688 32020
rect 16948 31968 17000 32020
rect 15292 31900 15344 31952
rect 15476 31832 15528 31884
rect 16304 31900 16356 31952
rect 16396 31900 16448 31952
rect 20720 31943 20772 31952
rect 14096 31764 14148 31816
rect 15108 31764 15160 31816
rect 12164 31696 12216 31748
rect 13176 31696 13228 31748
rect 13544 31696 13596 31748
rect 14648 31739 14700 31748
rect 14648 31705 14657 31739
rect 14657 31705 14691 31739
rect 14691 31705 14700 31739
rect 14648 31696 14700 31705
rect 15292 31739 15344 31748
rect 15292 31705 15302 31739
rect 15302 31705 15336 31739
rect 15336 31705 15344 31739
rect 15292 31696 15344 31705
rect 16120 31832 16172 31884
rect 17684 31832 17736 31884
rect 20076 31875 20128 31884
rect 20076 31841 20085 31875
rect 20085 31841 20119 31875
rect 20119 31841 20128 31875
rect 20076 31832 20128 31841
rect 20720 31909 20729 31943
rect 20729 31909 20763 31943
rect 20763 31909 20772 31943
rect 20720 31900 20772 31909
rect 22928 31968 22980 32020
rect 16672 31764 16724 31816
rect 17224 31764 17276 31816
rect 20996 31764 21048 31816
rect 21272 31807 21324 31816
rect 21272 31773 21281 31807
rect 21281 31773 21315 31807
rect 21315 31773 21324 31807
rect 21272 31764 21324 31773
rect 17592 31739 17644 31748
rect 17592 31705 17601 31739
rect 17601 31705 17635 31739
rect 17635 31705 17644 31739
rect 17592 31696 17644 31705
rect 17868 31696 17920 31748
rect 18880 31696 18932 31748
rect 19984 31739 20036 31748
rect 19984 31705 19993 31739
rect 19993 31705 20027 31739
rect 20027 31705 20036 31739
rect 19984 31696 20036 31705
rect 12256 31628 12308 31680
rect 13452 31628 13504 31680
rect 14924 31628 14976 31680
rect 15568 31628 15620 31680
rect 20996 31628 21048 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 1676 31467 1728 31476
rect 1676 31433 1685 31467
rect 1685 31433 1719 31467
rect 1719 31433 1728 31467
rect 1676 31424 1728 31433
rect 7104 31424 7156 31476
rect 9128 31424 9180 31476
rect 10140 31424 10192 31476
rect 12164 31424 12216 31476
rect 16580 31424 16632 31476
rect 16856 31424 16908 31476
rect 16948 31424 17000 31476
rect 18236 31424 18288 31476
rect 18604 31424 18656 31476
rect 4712 31356 4764 31408
rect 5816 31356 5868 31408
rect 7012 31356 7064 31408
rect 9496 31356 9548 31408
rect 10416 31356 10468 31408
rect 10600 31356 10652 31408
rect 2320 31288 2372 31340
rect 3424 31288 3476 31340
rect 3792 31288 3844 31340
rect 2780 31220 2832 31272
rect 5264 31220 5316 31272
rect 5540 31220 5592 31272
rect 5816 31220 5868 31272
rect 6736 31220 6788 31272
rect 8668 31331 8720 31340
rect 8668 31297 8677 31331
rect 8677 31297 8711 31331
rect 8711 31297 8720 31331
rect 8668 31288 8720 31297
rect 11244 31288 11296 31340
rect 13176 31356 13228 31408
rect 13544 31356 13596 31408
rect 14924 31356 14976 31408
rect 10784 31220 10836 31272
rect 11980 31220 12032 31272
rect 6092 31084 6144 31136
rect 6276 31084 6328 31136
rect 11244 31152 11296 31204
rect 13728 31331 13780 31340
rect 13728 31297 13737 31331
rect 13737 31297 13771 31331
rect 13771 31297 13780 31331
rect 13728 31288 13780 31297
rect 15568 31288 15620 31340
rect 15844 31288 15896 31340
rect 16304 31288 16356 31340
rect 17960 31288 18012 31340
rect 14280 31220 14332 31272
rect 16028 31220 16080 31272
rect 17868 31263 17920 31272
rect 17868 31229 17877 31263
rect 17877 31229 17911 31263
rect 17911 31229 17920 31263
rect 17868 31220 17920 31229
rect 19984 31424 20036 31476
rect 20996 31467 21048 31476
rect 20996 31433 21005 31467
rect 21005 31433 21039 31467
rect 21039 31433 21048 31467
rect 20996 31424 21048 31433
rect 21272 31424 21324 31476
rect 22928 31424 22980 31476
rect 20628 31356 20680 31408
rect 20536 31288 20588 31340
rect 20904 31331 20956 31340
rect 20904 31297 20913 31331
rect 20913 31297 20947 31331
rect 20947 31297 20956 31331
rect 20904 31288 20956 31297
rect 13360 31084 13412 31136
rect 15752 31084 15804 31136
rect 17776 31152 17828 31204
rect 18880 31220 18932 31272
rect 22100 31220 22152 31272
rect 22468 31220 22520 31272
rect 18420 31152 18472 31204
rect 18512 31127 18564 31136
rect 18512 31093 18521 31127
rect 18521 31093 18555 31127
rect 18555 31093 18564 31127
rect 18512 31084 18564 31093
rect 18604 31084 18656 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 6920 30880 6972 30932
rect 7932 30880 7984 30932
rect 11520 30880 11572 30932
rect 11980 30880 12032 30932
rect 6368 30812 6420 30864
rect 4252 30744 4304 30796
rect 5448 30787 5500 30796
rect 5448 30753 5457 30787
rect 5457 30753 5491 30787
rect 5491 30753 5500 30787
rect 5448 30744 5500 30753
rect 9312 30812 9364 30864
rect 10600 30812 10652 30864
rect 10876 30812 10928 30864
rect 1952 30676 2004 30728
rect 2872 30676 2924 30728
rect 4068 30676 4120 30728
rect 5724 30719 5776 30728
rect 5724 30685 5733 30719
rect 5733 30685 5767 30719
rect 5767 30685 5776 30719
rect 5724 30676 5776 30685
rect 8668 30676 8720 30728
rect 4804 30608 4856 30660
rect 5540 30608 5592 30660
rect 6920 30608 6972 30660
rect 1676 30583 1728 30592
rect 1676 30549 1685 30583
rect 1685 30549 1719 30583
rect 1719 30549 1728 30583
rect 1676 30540 1728 30549
rect 1860 30540 1912 30592
rect 2412 30583 2464 30592
rect 2412 30549 2421 30583
rect 2421 30549 2455 30583
rect 2455 30549 2464 30583
rect 2412 30540 2464 30549
rect 3240 30540 3292 30592
rect 11612 30744 11664 30796
rect 12348 30744 12400 30796
rect 12716 30880 12768 30932
rect 15660 30880 15712 30932
rect 16028 30880 16080 30932
rect 18420 30880 18472 30932
rect 23020 30923 23072 30932
rect 12808 30812 12860 30864
rect 13728 30812 13780 30864
rect 14556 30812 14608 30864
rect 15568 30812 15620 30864
rect 13452 30744 13504 30796
rect 9588 30719 9640 30728
rect 9588 30685 9597 30719
rect 9597 30685 9631 30719
rect 9631 30685 9640 30719
rect 9588 30676 9640 30685
rect 10232 30719 10284 30728
rect 10232 30685 10241 30719
rect 10241 30685 10275 30719
rect 10275 30685 10284 30719
rect 10232 30676 10284 30685
rect 10600 30676 10652 30728
rect 12808 30676 12860 30728
rect 13084 30719 13136 30728
rect 13084 30685 13093 30719
rect 13093 30685 13127 30719
rect 13127 30685 13136 30719
rect 13084 30676 13136 30685
rect 16672 30719 16724 30728
rect 10508 30608 10560 30660
rect 9680 30583 9732 30592
rect 9680 30549 9689 30583
rect 9689 30549 9723 30583
rect 9723 30549 9732 30583
rect 9680 30540 9732 30549
rect 11612 30540 11664 30592
rect 12716 30608 12768 30660
rect 16672 30685 16681 30719
rect 16681 30685 16715 30719
rect 16715 30685 16724 30719
rect 16672 30676 16724 30685
rect 18420 30676 18472 30728
rect 15476 30651 15528 30660
rect 15476 30617 15485 30651
rect 15485 30617 15519 30651
rect 15519 30617 15528 30651
rect 15476 30608 15528 30617
rect 17040 30608 17092 30660
rect 17316 30651 17368 30660
rect 17316 30617 17325 30651
rect 17325 30617 17359 30651
rect 17359 30617 17368 30651
rect 17316 30608 17368 30617
rect 18788 30608 18840 30660
rect 19984 30608 20036 30660
rect 20536 30744 20588 30796
rect 20904 30676 20956 30728
rect 23020 30889 23029 30923
rect 23029 30889 23063 30923
rect 23063 30889 23072 30923
rect 23020 30880 23072 30889
rect 25688 30744 25740 30796
rect 24124 30676 24176 30728
rect 15660 30540 15712 30592
rect 16580 30583 16632 30592
rect 16580 30549 16589 30583
rect 16589 30549 16623 30583
rect 16623 30549 16632 30583
rect 16580 30540 16632 30549
rect 18420 30583 18472 30592
rect 18420 30549 18429 30583
rect 18429 30549 18463 30583
rect 18463 30549 18472 30583
rect 18420 30540 18472 30549
rect 19340 30540 19392 30592
rect 23020 30608 23072 30660
rect 20720 30583 20772 30592
rect 20720 30549 20729 30583
rect 20729 30549 20763 30583
rect 20763 30549 20772 30583
rect 20720 30540 20772 30549
rect 22100 30540 22152 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 4252 30336 4304 30388
rect 5908 30336 5960 30388
rect 6368 30336 6420 30388
rect 9680 30336 9732 30388
rect 14004 30336 14056 30388
rect 14280 30336 14332 30388
rect 15936 30336 15988 30388
rect 16856 30336 16908 30388
rect 18788 30336 18840 30388
rect 19064 30336 19116 30388
rect 20720 30336 20772 30388
rect 3424 30268 3476 30320
rect 3608 30268 3660 30320
rect 6828 30268 6880 30320
rect 8668 30268 8720 30320
rect 2412 30200 2464 30252
rect 3792 30243 3844 30252
rect 3792 30209 3801 30243
rect 3801 30209 3835 30243
rect 3835 30209 3844 30243
rect 3792 30200 3844 30209
rect 6000 30243 6052 30252
rect 6000 30209 6009 30243
rect 6009 30209 6043 30243
rect 6043 30209 6052 30243
rect 6000 30200 6052 30209
rect 6736 30200 6788 30252
rect 3424 30132 3476 30184
rect 5264 30132 5316 30184
rect 7104 30132 7156 30184
rect 7288 30132 7340 30184
rect 7748 30132 7800 30184
rect 8300 30132 8352 30184
rect 11888 30268 11940 30320
rect 11980 30311 12032 30320
rect 11980 30277 11989 30311
rect 11989 30277 12023 30311
rect 12023 30277 12032 30311
rect 11980 30268 12032 30277
rect 10048 30200 10100 30252
rect 10324 30243 10376 30252
rect 10324 30209 10333 30243
rect 10333 30209 10367 30243
rect 10367 30209 10376 30243
rect 10324 30200 10376 30209
rect 10968 30243 11020 30252
rect 10968 30209 10977 30243
rect 10977 30209 11011 30243
rect 11011 30209 11020 30243
rect 10968 30200 11020 30209
rect 11060 30200 11112 30252
rect 11612 30200 11664 30252
rect 13084 30200 13136 30252
rect 11336 30132 11388 30184
rect 11704 30175 11756 30184
rect 11704 30141 11713 30175
rect 11713 30141 11747 30175
rect 11747 30141 11756 30175
rect 11704 30132 11756 30141
rect 12072 30132 12124 30184
rect 15844 30268 15896 30320
rect 17776 30268 17828 30320
rect 19340 30268 19392 30320
rect 19524 30311 19576 30320
rect 19524 30277 19533 30311
rect 19533 30277 19567 30311
rect 19567 30277 19576 30311
rect 19524 30268 19576 30277
rect 19800 30268 19852 30320
rect 22100 30268 22152 30320
rect 14280 30200 14332 30252
rect 14924 30200 14976 30252
rect 16672 30200 16724 30252
rect 14556 30132 14608 30184
rect 15568 30175 15620 30184
rect 9312 30064 9364 30116
rect 13452 30107 13504 30116
rect 4620 29996 4672 30048
rect 5540 29996 5592 30048
rect 6000 29996 6052 30048
rect 6276 29996 6328 30048
rect 10324 29996 10376 30048
rect 11060 30039 11112 30048
rect 11060 30005 11069 30039
rect 11069 30005 11103 30039
rect 11103 30005 11112 30039
rect 11060 29996 11112 30005
rect 13452 30073 13461 30107
rect 13461 30073 13495 30107
rect 13495 30073 13504 30107
rect 13452 30064 13504 30073
rect 14648 30064 14700 30116
rect 15568 30141 15577 30175
rect 15577 30141 15611 30175
rect 15611 30141 15620 30175
rect 15568 30132 15620 30141
rect 16764 30132 16816 30184
rect 17868 30175 17920 30184
rect 17868 30141 17877 30175
rect 17877 30141 17911 30175
rect 17911 30141 17920 30175
rect 17868 30132 17920 30141
rect 18052 30132 18104 30184
rect 19156 30132 19208 30184
rect 19800 30064 19852 30116
rect 21548 30200 21600 30252
rect 20076 30132 20128 30184
rect 20720 30064 20772 30116
rect 13176 29996 13228 30048
rect 13728 29996 13780 30048
rect 14832 29996 14884 30048
rect 17132 29996 17184 30048
rect 18328 29996 18380 30048
rect 19892 29996 19944 30048
rect 37832 30132 37884 30184
rect 38292 30175 38344 30184
rect 38292 30141 38301 30175
rect 38301 30141 38335 30175
rect 38335 30141 38344 30175
rect 38292 30132 38344 30141
rect 20904 30064 20956 30116
rect 22928 29996 22980 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 1768 29792 1820 29844
rect 6644 29792 6696 29844
rect 6828 29792 6880 29844
rect 11336 29792 11388 29844
rect 13084 29792 13136 29844
rect 18512 29792 18564 29844
rect 19524 29792 19576 29844
rect 38292 29835 38344 29844
rect 38292 29801 38301 29835
rect 38301 29801 38335 29835
rect 38335 29801 38344 29835
rect 38292 29792 38344 29801
rect 2412 29656 2464 29708
rect 3608 29656 3660 29708
rect 3792 29656 3844 29708
rect 5540 29656 5592 29708
rect 5724 29656 5776 29708
rect 6736 29656 6788 29708
rect 9864 29724 9916 29776
rect 12624 29724 12676 29776
rect 13452 29724 13504 29776
rect 8300 29656 8352 29708
rect 10416 29656 10468 29708
rect 3056 29588 3108 29640
rect 6276 29588 6328 29640
rect 9312 29631 9364 29640
rect 1676 29452 1728 29504
rect 3240 29452 3292 29504
rect 3792 29452 3844 29504
rect 6828 29520 6880 29572
rect 4620 29452 4672 29504
rect 4896 29452 4948 29504
rect 5632 29452 5684 29504
rect 5816 29452 5868 29504
rect 6000 29452 6052 29504
rect 6920 29452 6972 29504
rect 9312 29597 9321 29631
rect 9321 29597 9355 29631
rect 9355 29597 9364 29631
rect 9312 29588 9364 29597
rect 9588 29588 9640 29640
rect 11244 29656 11296 29708
rect 11704 29656 11756 29708
rect 13268 29699 13320 29708
rect 13268 29665 13277 29699
rect 13277 29665 13311 29699
rect 13311 29665 13320 29699
rect 13268 29656 13320 29665
rect 9128 29520 9180 29572
rect 9496 29520 9548 29572
rect 9680 29520 9732 29572
rect 10140 29520 10192 29572
rect 10232 29520 10284 29572
rect 11612 29520 11664 29572
rect 11796 29520 11848 29572
rect 13176 29563 13228 29572
rect 13176 29529 13185 29563
rect 13185 29529 13219 29563
rect 13219 29529 13228 29563
rect 13176 29520 13228 29529
rect 7932 29452 7984 29504
rect 8024 29452 8076 29504
rect 8484 29452 8536 29504
rect 8760 29452 8812 29504
rect 15476 29724 15528 29776
rect 16212 29724 16264 29776
rect 16672 29724 16724 29776
rect 20904 29724 20956 29776
rect 13820 29656 13872 29708
rect 14648 29699 14700 29708
rect 14648 29665 14657 29699
rect 14657 29665 14691 29699
rect 14691 29665 14700 29699
rect 14648 29656 14700 29665
rect 18052 29656 18104 29708
rect 18788 29699 18840 29708
rect 18788 29665 18797 29699
rect 18797 29665 18831 29699
rect 18831 29665 18840 29699
rect 18788 29656 18840 29665
rect 18972 29656 19024 29708
rect 20076 29656 20128 29708
rect 20444 29656 20496 29708
rect 13912 29588 13964 29640
rect 22100 29656 22152 29708
rect 21916 29588 21968 29640
rect 14924 29520 14976 29572
rect 13912 29452 13964 29504
rect 14464 29452 14516 29504
rect 15936 29520 15988 29572
rect 16396 29520 16448 29572
rect 17040 29563 17092 29572
rect 17040 29529 17049 29563
rect 17049 29529 17083 29563
rect 17083 29529 17092 29563
rect 17040 29520 17092 29529
rect 17132 29563 17184 29572
rect 17132 29529 17141 29563
rect 17141 29529 17175 29563
rect 17175 29529 17184 29563
rect 17132 29520 17184 29529
rect 17776 29520 17828 29572
rect 18696 29563 18748 29572
rect 18696 29529 18705 29563
rect 18705 29529 18739 29563
rect 18739 29529 18748 29563
rect 18696 29520 18748 29529
rect 20076 29520 20128 29572
rect 20260 29520 20312 29572
rect 16580 29452 16632 29504
rect 16672 29452 16724 29504
rect 19064 29452 19116 29504
rect 19892 29452 19944 29504
rect 20444 29563 20496 29572
rect 20444 29529 20453 29563
rect 20453 29529 20487 29563
rect 20487 29529 20496 29563
rect 20444 29520 20496 29529
rect 20996 29452 21048 29504
rect 21732 29495 21784 29504
rect 21732 29461 21741 29495
rect 21741 29461 21775 29495
rect 21775 29461 21784 29495
rect 21732 29452 21784 29461
rect 38016 29452 38068 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 1676 29291 1728 29300
rect 1676 29257 1685 29291
rect 1685 29257 1719 29291
rect 1719 29257 1728 29291
rect 1676 29248 1728 29257
rect 4804 29248 4856 29300
rect 5632 29248 5684 29300
rect 6000 29248 6052 29300
rect 5356 29180 5408 29232
rect 8760 29248 8812 29300
rect 6644 29223 6696 29232
rect 6644 29189 6653 29223
rect 6653 29189 6687 29223
rect 6687 29189 6696 29223
rect 6644 29180 6696 29189
rect 8668 29180 8720 29232
rect 9772 29180 9824 29232
rect 10416 29248 10468 29300
rect 11060 29248 11112 29300
rect 1860 29112 1912 29164
rect 2412 29112 2464 29164
rect 3240 29155 3292 29164
rect 3240 29121 3249 29155
rect 3249 29121 3283 29155
rect 3283 29121 3292 29155
rect 3240 29112 3292 29121
rect 4620 29112 4672 29164
rect 2780 29044 2832 29096
rect 4528 29044 4580 29096
rect 6736 29112 6788 29164
rect 7380 29112 7432 29164
rect 8208 29112 8260 29164
rect 6644 29044 6696 29096
rect 6276 28976 6328 29028
rect 3608 28908 3660 28960
rect 4528 28908 4580 28960
rect 4804 28908 4856 28960
rect 10508 29044 10560 29096
rect 11244 29180 11296 29232
rect 11520 29112 11572 29164
rect 13544 29180 13596 29232
rect 13728 29223 13780 29232
rect 13728 29189 13737 29223
rect 13737 29189 13771 29223
rect 13771 29189 13780 29223
rect 13728 29180 13780 29189
rect 14556 29223 14608 29232
rect 14556 29189 14565 29223
rect 14565 29189 14599 29223
rect 14599 29189 14608 29223
rect 15752 29223 15804 29232
rect 14556 29180 14608 29189
rect 15752 29189 15761 29223
rect 15761 29189 15795 29223
rect 15795 29189 15804 29223
rect 15752 29180 15804 29189
rect 15936 29180 15988 29232
rect 16304 29223 16356 29232
rect 16304 29189 16313 29223
rect 16313 29189 16347 29223
rect 16347 29189 16356 29223
rect 16304 29180 16356 29189
rect 19156 29248 19208 29300
rect 11704 29044 11756 29096
rect 11060 29019 11112 29028
rect 11060 28985 11069 29019
rect 11069 28985 11103 29019
rect 11103 28985 11112 29019
rect 11060 28976 11112 28985
rect 11336 28976 11388 29028
rect 11796 28976 11848 29028
rect 13176 29044 13228 29096
rect 14464 29044 14516 29096
rect 18420 29180 18472 29232
rect 19248 29223 19300 29232
rect 19248 29189 19257 29223
rect 19257 29189 19291 29223
rect 19291 29189 19300 29223
rect 19248 29180 19300 29189
rect 19524 29180 19576 29232
rect 20444 29223 20496 29232
rect 20444 29189 20453 29223
rect 20453 29189 20487 29223
rect 20487 29189 20496 29223
rect 20444 29180 20496 29189
rect 20996 29248 21048 29300
rect 23204 29248 23256 29300
rect 21732 29180 21784 29232
rect 16672 29112 16724 29164
rect 20812 29112 20864 29164
rect 16580 29044 16632 29096
rect 18696 29044 18748 29096
rect 16212 28976 16264 29028
rect 16948 29019 17000 29028
rect 16948 28985 16957 29019
rect 16957 28985 16991 29019
rect 16991 28985 17000 29019
rect 16948 28976 17000 28985
rect 17776 28976 17828 29028
rect 15292 28908 15344 28960
rect 15384 28908 15436 28960
rect 18328 28908 18380 28960
rect 19340 28976 19392 29028
rect 21548 28976 21600 29028
rect 24124 29112 24176 29164
rect 38016 29087 38068 29096
rect 38016 29053 38025 29087
rect 38025 29053 38059 29087
rect 38059 29053 38068 29087
rect 38016 29044 38068 29053
rect 38292 29087 38344 29096
rect 38292 29053 38301 29087
rect 38301 29053 38335 29087
rect 38335 29053 38344 29087
rect 38292 29044 38344 29053
rect 23204 28976 23256 29028
rect 23388 28976 23440 29028
rect 36636 28976 36688 29028
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 4620 28704 4672 28756
rect 11796 28704 11848 28756
rect 14372 28747 14424 28756
rect 14372 28713 14381 28747
rect 14381 28713 14415 28747
rect 14415 28713 14424 28747
rect 14372 28704 14424 28713
rect 14832 28704 14884 28756
rect 17224 28704 17276 28756
rect 17684 28704 17736 28756
rect 3976 28636 4028 28688
rect 4160 28636 4212 28688
rect 4988 28636 5040 28688
rect 5356 28679 5408 28688
rect 5356 28645 5365 28679
rect 5365 28645 5399 28679
rect 5399 28645 5408 28679
rect 5356 28636 5408 28645
rect 7012 28636 7064 28688
rect 7288 28636 7340 28688
rect 10232 28636 10284 28688
rect 16120 28636 16172 28688
rect 17776 28636 17828 28688
rect 19248 28704 19300 28756
rect 20444 28704 20496 28756
rect 22560 28704 22612 28756
rect 23296 28747 23348 28756
rect 23296 28713 23305 28747
rect 23305 28713 23339 28747
rect 23339 28713 23348 28747
rect 23296 28704 23348 28713
rect 17960 28636 18012 28688
rect 4712 28568 4764 28620
rect 6644 28568 6696 28620
rect 2412 28500 2464 28552
rect 4620 28543 4672 28552
rect 4620 28509 4629 28543
rect 4629 28509 4663 28543
rect 4663 28509 4672 28543
rect 5264 28543 5316 28552
rect 4620 28500 4672 28509
rect 5264 28509 5273 28543
rect 5273 28509 5307 28543
rect 5307 28509 5316 28543
rect 5264 28500 5316 28509
rect 8668 28568 8720 28620
rect 11428 28568 11480 28620
rect 11704 28568 11756 28620
rect 15108 28568 15160 28620
rect 15752 28568 15804 28620
rect 16580 28568 16632 28620
rect 16856 28568 16908 28620
rect 7288 28500 7340 28552
rect 7932 28500 7984 28552
rect 8024 28500 8076 28552
rect 9036 28500 9088 28552
rect 6736 28432 6788 28484
rect 1676 28407 1728 28416
rect 1676 28373 1685 28407
rect 1685 28373 1719 28407
rect 1719 28373 1728 28407
rect 1676 28364 1728 28373
rect 2596 28364 2648 28416
rect 2780 28364 2832 28416
rect 4252 28364 4304 28416
rect 6828 28364 6880 28416
rect 9220 28432 9272 28484
rect 9312 28432 9364 28484
rect 12256 28500 12308 28552
rect 12992 28500 13044 28552
rect 13268 28500 13320 28552
rect 11152 28432 11204 28484
rect 9772 28364 9824 28416
rect 9956 28364 10008 28416
rect 10968 28364 11020 28416
rect 11704 28364 11756 28416
rect 13176 28432 13228 28484
rect 15200 28432 15252 28484
rect 16396 28432 16448 28484
rect 12808 28364 12860 28416
rect 13360 28364 13412 28416
rect 13728 28364 13780 28416
rect 15568 28364 15620 28416
rect 17684 28432 17736 28484
rect 19892 28568 19944 28620
rect 19984 28568 20036 28620
rect 19524 28500 19576 28552
rect 19616 28500 19668 28552
rect 20168 28500 20220 28552
rect 20812 28500 20864 28552
rect 23756 28636 23808 28688
rect 38292 28679 38344 28688
rect 38292 28645 38301 28679
rect 38301 28645 38335 28679
rect 38335 28645 38344 28679
rect 38292 28636 38344 28645
rect 21732 28611 21784 28620
rect 21732 28577 21741 28611
rect 21741 28577 21775 28611
rect 21775 28577 21784 28611
rect 21732 28568 21784 28577
rect 19524 28364 19576 28416
rect 20536 28364 20588 28416
rect 38016 28432 38068 28484
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 2780 28160 2832 28212
rect 5264 28160 5316 28212
rect 4068 28092 4120 28144
rect 1768 28024 1820 28076
rect 3240 28024 3292 28076
rect 2412 27956 2464 28008
rect 2596 27956 2648 28008
rect 2872 27956 2924 28008
rect 3792 28024 3844 28076
rect 4620 28024 4672 28076
rect 5264 28024 5316 28076
rect 7472 28160 7524 28212
rect 7656 28160 7708 28212
rect 9772 28160 9824 28212
rect 8300 28092 8352 28144
rect 10048 28092 10100 28144
rect 10232 28092 10284 28144
rect 12532 28160 12584 28212
rect 16120 28160 16172 28212
rect 14924 28092 14976 28144
rect 6828 28067 6880 28076
rect 6828 28033 6837 28067
rect 6837 28033 6871 28067
rect 6871 28033 6880 28067
rect 6828 28024 6880 28033
rect 7288 28024 7340 28076
rect 7472 28067 7524 28076
rect 7472 28033 7481 28067
rect 7481 28033 7515 28067
rect 7515 28033 7524 28067
rect 7472 28024 7524 28033
rect 11612 28024 11664 28076
rect 7196 27956 7248 28008
rect 10416 27956 10468 28008
rect 11244 27956 11296 28008
rect 11336 27956 11388 28008
rect 5080 27888 5132 27940
rect 4252 27820 4304 27872
rect 6276 27888 6328 27940
rect 8668 27888 8720 27940
rect 11152 27888 11204 27940
rect 13636 27888 13688 27940
rect 14832 27888 14884 27940
rect 15384 27956 15436 28008
rect 15660 27888 15712 27940
rect 9036 27863 9088 27872
rect 9036 27829 9045 27863
rect 9045 27829 9079 27863
rect 9079 27829 9088 27863
rect 9036 27820 9088 27829
rect 9956 27820 10008 27872
rect 11520 27820 11572 27872
rect 12348 27820 12400 27872
rect 13084 27820 13136 27872
rect 15200 27820 15252 27872
rect 17408 28135 17460 28144
rect 17408 28101 17417 28135
rect 17417 28101 17451 28135
rect 17451 28101 17460 28135
rect 17408 28092 17460 28101
rect 23756 28203 23808 28212
rect 23756 28169 23765 28203
rect 23765 28169 23799 28203
rect 23799 28169 23808 28203
rect 23756 28160 23808 28169
rect 19432 28092 19484 28144
rect 23388 28092 23440 28144
rect 20444 28024 20496 28076
rect 20720 28024 20772 28076
rect 21732 28024 21784 28076
rect 18328 27999 18380 28008
rect 18328 27965 18337 27999
rect 18337 27965 18371 27999
rect 18371 27965 18380 27999
rect 18328 27956 18380 27965
rect 18512 27956 18564 28008
rect 18604 27956 18656 28008
rect 21364 27999 21416 28008
rect 21364 27965 21373 27999
rect 21373 27965 21407 27999
rect 21407 27965 21416 27999
rect 21364 27956 21416 27965
rect 16488 27888 16540 27940
rect 18880 27888 18932 27940
rect 17592 27820 17644 27872
rect 20444 27888 20496 27940
rect 24676 28024 24728 28076
rect 23388 27888 23440 27940
rect 37740 27888 37792 27940
rect 19524 27863 19576 27872
rect 19524 27829 19533 27863
rect 19533 27829 19567 27863
rect 19567 27829 19576 27863
rect 19524 27820 19576 27829
rect 19984 27820 20036 27872
rect 22560 27820 22612 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 3424 27616 3476 27668
rect 10140 27616 10192 27668
rect 10416 27616 10468 27668
rect 12992 27616 13044 27668
rect 3056 27548 3108 27600
rect 4068 27591 4120 27600
rect 4068 27557 4077 27591
rect 4077 27557 4111 27591
rect 4111 27557 4120 27591
rect 4068 27548 4120 27557
rect 5724 27548 5776 27600
rect 6092 27548 6144 27600
rect 2688 27480 2740 27532
rect 3792 27480 3844 27532
rect 1676 27412 1728 27464
rect 2688 27344 2740 27396
rect 4344 27412 4396 27464
rect 5264 27480 5316 27532
rect 10048 27548 10100 27600
rect 9864 27480 9916 27532
rect 12164 27548 12216 27600
rect 8116 27412 8168 27464
rect 3240 27344 3292 27396
rect 3792 27344 3844 27396
rect 6828 27344 6880 27396
rect 8760 27344 8812 27396
rect 11428 27523 11480 27532
rect 11428 27489 11437 27523
rect 11437 27489 11471 27523
rect 11471 27489 11480 27523
rect 11428 27480 11480 27489
rect 12440 27480 12492 27532
rect 12808 27480 12860 27532
rect 12900 27455 12952 27464
rect 12900 27421 12909 27455
rect 12909 27421 12943 27455
rect 12943 27421 12952 27455
rect 12900 27412 12952 27421
rect 14556 27548 14608 27600
rect 16856 27616 16908 27668
rect 20352 27616 20404 27668
rect 15384 27548 15436 27600
rect 16396 27591 16448 27600
rect 16396 27557 16405 27591
rect 16405 27557 16439 27591
rect 16439 27557 16448 27591
rect 16396 27548 16448 27557
rect 18788 27548 18840 27600
rect 14372 27523 14424 27532
rect 14372 27489 14381 27523
rect 14381 27489 14415 27523
rect 14415 27489 14424 27523
rect 17592 27523 17644 27532
rect 14372 27480 14424 27489
rect 14188 27412 14240 27464
rect 16120 27412 16172 27464
rect 17592 27489 17601 27523
rect 17601 27489 17635 27523
rect 17635 27489 17644 27523
rect 17592 27480 17644 27489
rect 19524 27480 19576 27532
rect 20628 27480 20680 27532
rect 19984 27412 20036 27464
rect 10508 27387 10560 27396
rect 10508 27353 10517 27387
rect 10517 27353 10551 27387
rect 10551 27353 10560 27387
rect 10508 27344 10560 27353
rect 11520 27344 11572 27396
rect 5540 27276 5592 27328
rect 6644 27276 6696 27328
rect 6920 27276 6972 27328
rect 7380 27276 7432 27328
rect 9128 27276 9180 27328
rect 9772 27276 9824 27328
rect 13084 27344 13136 27396
rect 13268 27344 13320 27396
rect 13360 27344 13412 27396
rect 12532 27276 12584 27328
rect 12716 27276 12768 27328
rect 13452 27276 13504 27328
rect 15568 27344 15620 27396
rect 16396 27344 16448 27396
rect 17500 27387 17552 27396
rect 17500 27353 17509 27387
rect 17509 27353 17543 27387
rect 17543 27353 17552 27387
rect 17500 27344 17552 27353
rect 18696 27387 18748 27396
rect 15292 27276 15344 27328
rect 18696 27353 18705 27387
rect 18705 27353 18739 27387
rect 18739 27353 18748 27387
rect 18696 27344 18748 27353
rect 20536 27344 20588 27396
rect 20996 27344 21048 27396
rect 21272 27548 21324 27600
rect 22008 27548 22060 27600
rect 21640 27412 21692 27464
rect 34520 27344 34572 27396
rect 19340 27276 19392 27328
rect 19984 27276 20036 27328
rect 21272 27276 21324 27328
rect 21824 27319 21876 27328
rect 21824 27285 21833 27319
rect 21833 27285 21867 27319
rect 21867 27285 21876 27319
rect 21824 27276 21876 27285
rect 23388 27319 23440 27328
rect 23388 27285 23397 27319
rect 23397 27285 23431 27319
rect 23431 27285 23440 27319
rect 23388 27276 23440 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 2228 27072 2280 27124
rect 3700 27115 3752 27124
rect 3700 27081 3709 27115
rect 3709 27081 3743 27115
rect 3743 27081 3752 27115
rect 3700 27072 3752 27081
rect 7104 27072 7156 27124
rect 7564 27072 7616 27124
rect 10508 27072 10560 27124
rect 12072 27072 12124 27124
rect 8484 27004 8536 27056
rect 8576 27004 8628 27056
rect 9496 27047 9548 27056
rect 9496 27013 9505 27047
rect 9505 27013 9539 27047
rect 9539 27013 9548 27047
rect 9496 27004 9548 27013
rect 11152 27004 11204 27056
rect 12440 27047 12492 27056
rect 12440 27013 12449 27047
rect 12449 27013 12483 27047
rect 12483 27013 12492 27047
rect 13728 27047 13780 27056
rect 12440 27004 12492 27013
rect 13728 27013 13737 27047
rect 13737 27013 13771 27047
rect 13771 27013 13780 27047
rect 13728 27004 13780 27013
rect 15108 27072 15160 27124
rect 14556 27047 14608 27056
rect 14556 27013 14565 27047
rect 14565 27013 14599 27047
rect 14599 27013 14608 27047
rect 14556 27004 14608 27013
rect 16948 27004 17000 27056
rect 17868 27004 17920 27056
rect 20720 27072 20772 27124
rect 19340 27004 19392 27056
rect 19800 27004 19852 27056
rect 22652 27004 22704 27056
rect 23296 27004 23348 27056
rect 2872 26936 2924 26988
rect 3792 26979 3844 26988
rect 3792 26945 3801 26979
rect 3801 26945 3835 26979
rect 3835 26945 3844 26979
rect 3792 26936 3844 26945
rect 10232 26936 10284 26988
rect 10968 26979 11020 26988
rect 10968 26945 10977 26979
rect 10977 26945 11011 26979
rect 11011 26945 11020 26979
rect 10968 26936 11020 26945
rect 16396 26936 16448 26988
rect 21364 26979 21416 26988
rect 21364 26945 21373 26979
rect 21373 26945 21407 26979
rect 21407 26945 21416 26979
rect 21364 26936 21416 26945
rect 5080 26868 5132 26920
rect 8024 26868 8076 26920
rect 9864 26868 9916 26920
rect 11152 26868 11204 26920
rect 14280 26868 14332 26920
rect 6828 26800 6880 26852
rect 7472 26843 7524 26852
rect 7472 26809 7481 26843
rect 7481 26809 7515 26843
rect 7515 26809 7524 26843
rect 7472 26800 7524 26809
rect 1676 26775 1728 26784
rect 1676 26741 1685 26775
rect 1685 26741 1719 26775
rect 1719 26741 1728 26775
rect 1676 26732 1728 26741
rect 4344 26775 4396 26784
rect 4344 26741 4353 26775
rect 4353 26741 4387 26775
rect 4387 26741 4396 26775
rect 4344 26732 4396 26741
rect 4620 26732 4672 26784
rect 5080 26732 5132 26784
rect 5356 26775 5408 26784
rect 5356 26741 5365 26775
rect 5365 26741 5399 26775
rect 5399 26741 5408 26775
rect 5356 26732 5408 26741
rect 5540 26732 5592 26784
rect 6000 26732 6052 26784
rect 9128 26732 9180 26784
rect 9956 26732 10008 26784
rect 10692 26732 10744 26784
rect 12072 26800 12124 26852
rect 12532 26732 12584 26784
rect 13084 26732 13136 26784
rect 16120 26868 16172 26920
rect 14740 26732 14792 26784
rect 15292 26732 15344 26784
rect 15844 26800 15896 26852
rect 17592 26868 17644 26920
rect 18420 26911 18472 26920
rect 18420 26877 18429 26911
rect 18429 26877 18463 26911
rect 18463 26877 18472 26911
rect 18420 26868 18472 26877
rect 18972 26868 19024 26920
rect 19432 26868 19484 26920
rect 20260 26911 20312 26920
rect 20260 26877 20269 26911
rect 20269 26877 20303 26911
rect 20303 26877 20312 26911
rect 20260 26868 20312 26877
rect 20628 26868 20680 26920
rect 36636 26936 36688 26988
rect 19524 26732 19576 26784
rect 21640 26800 21692 26852
rect 21824 26800 21876 26852
rect 23572 26911 23624 26920
rect 22468 26800 22520 26852
rect 23572 26877 23581 26911
rect 23581 26877 23615 26911
rect 23615 26877 23624 26911
rect 23572 26868 23624 26877
rect 20260 26732 20312 26784
rect 29828 26732 29880 26784
rect 38200 26775 38252 26784
rect 38200 26741 38209 26775
rect 38209 26741 38243 26775
rect 38243 26741 38252 26775
rect 38200 26732 38252 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 2044 26528 2096 26580
rect 2136 26528 2188 26580
rect 3332 26528 3384 26580
rect 4804 26528 4856 26580
rect 12440 26528 12492 26580
rect 12532 26571 12584 26580
rect 12532 26537 12541 26571
rect 12541 26537 12575 26571
rect 12575 26537 12584 26571
rect 12532 26528 12584 26537
rect 12716 26528 12768 26580
rect 13084 26460 13136 26512
rect 17408 26528 17460 26580
rect 18236 26528 18288 26580
rect 18420 26528 18472 26580
rect 22468 26528 22520 26580
rect 22652 26571 22704 26580
rect 22652 26537 22661 26571
rect 22661 26537 22695 26571
rect 22695 26537 22704 26571
rect 22652 26528 22704 26537
rect 23296 26571 23348 26580
rect 23296 26537 23305 26571
rect 23305 26537 23339 26571
rect 23339 26537 23348 26571
rect 23296 26528 23348 26537
rect 29828 26571 29880 26580
rect 29828 26537 29837 26571
rect 29837 26537 29871 26571
rect 29871 26537 29880 26571
rect 29828 26528 29880 26537
rect 6552 26392 6604 26444
rect 2228 26324 2280 26376
rect 2688 26367 2740 26376
rect 2688 26333 2697 26367
rect 2697 26333 2731 26367
rect 2731 26333 2740 26367
rect 2688 26324 2740 26333
rect 2872 26324 2924 26376
rect 7288 26367 7340 26376
rect 7288 26333 7297 26367
rect 7297 26333 7331 26367
rect 7331 26333 7340 26367
rect 7288 26324 7340 26333
rect 8392 26367 8444 26376
rect 2596 26256 2648 26308
rect 5540 26299 5592 26308
rect 5540 26265 5549 26299
rect 5549 26265 5583 26299
rect 5583 26265 5592 26299
rect 5540 26256 5592 26265
rect 8392 26333 8401 26367
rect 8401 26333 8435 26367
rect 8435 26333 8444 26367
rect 8392 26324 8444 26333
rect 9036 26324 9088 26376
rect 8944 26256 8996 26308
rect 9220 26299 9272 26308
rect 9220 26265 9229 26299
rect 9229 26265 9263 26299
rect 9263 26265 9272 26299
rect 9220 26256 9272 26265
rect 9312 26299 9364 26308
rect 9312 26265 9321 26299
rect 9321 26265 9355 26299
rect 9355 26265 9364 26299
rect 9312 26256 9364 26265
rect 9864 26256 9916 26308
rect 10232 26299 10284 26308
rect 10232 26265 10241 26299
rect 10241 26265 10275 26299
rect 10275 26265 10284 26299
rect 10232 26256 10284 26265
rect 10508 26392 10560 26444
rect 10784 26392 10836 26444
rect 11336 26435 11388 26444
rect 11336 26401 11345 26435
rect 11345 26401 11379 26435
rect 11379 26401 11388 26435
rect 11336 26392 11388 26401
rect 11796 26392 11848 26444
rect 12716 26324 12768 26376
rect 13084 26299 13136 26308
rect 13084 26265 13093 26299
rect 13093 26265 13127 26299
rect 13127 26265 13136 26299
rect 13084 26256 13136 26265
rect 13360 26256 13412 26308
rect 13728 26299 13780 26308
rect 13728 26265 13737 26299
rect 13737 26265 13771 26299
rect 13771 26265 13780 26299
rect 13728 26256 13780 26265
rect 14004 26460 14056 26512
rect 15384 26460 15436 26512
rect 15752 26460 15804 26512
rect 16488 26392 16540 26444
rect 14740 26324 14792 26376
rect 4988 26188 5040 26240
rect 5356 26188 5408 26240
rect 8392 26188 8444 26240
rect 9128 26188 9180 26240
rect 11336 26188 11388 26240
rect 14832 26256 14884 26308
rect 15384 26256 15436 26308
rect 16304 26324 16356 26376
rect 17592 26392 17644 26444
rect 20628 26460 20680 26512
rect 20536 26392 20588 26444
rect 26240 26392 26292 26444
rect 18788 26367 18840 26376
rect 18788 26333 18797 26367
rect 18797 26333 18831 26367
rect 18831 26333 18840 26367
rect 18788 26324 18840 26333
rect 19340 26324 19392 26376
rect 20904 26367 20956 26376
rect 20904 26333 20913 26367
rect 20913 26333 20947 26367
rect 20947 26333 20956 26367
rect 20904 26324 20956 26333
rect 22744 26367 22796 26376
rect 22744 26333 22753 26367
rect 22753 26333 22787 26367
rect 22787 26333 22796 26367
rect 22744 26324 22796 26333
rect 23204 26367 23256 26376
rect 23204 26333 23213 26367
rect 23213 26333 23247 26367
rect 23247 26333 23256 26367
rect 23204 26324 23256 26333
rect 37924 26324 37976 26376
rect 17316 26299 17368 26308
rect 17316 26265 17325 26299
rect 17325 26265 17359 26299
rect 17359 26265 17368 26299
rect 17316 26256 17368 26265
rect 18236 26188 18288 26240
rect 19156 26188 19208 26240
rect 19524 26188 19576 26240
rect 21364 26256 21416 26308
rect 19800 26188 19852 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 1308 25984 1360 26036
rect 2504 25984 2556 26036
rect 7748 25984 7800 26036
rect 11796 26027 11848 26036
rect 3884 25916 3936 25968
rect 2872 25848 2924 25900
rect 5816 25891 5868 25900
rect 5816 25857 5825 25891
rect 5825 25857 5859 25891
rect 5859 25857 5868 25891
rect 5816 25848 5868 25857
rect 7104 25891 7156 25900
rect 7104 25857 7113 25891
rect 7113 25857 7147 25891
rect 7147 25857 7156 25891
rect 7104 25848 7156 25857
rect 7656 25848 7708 25900
rect 7932 25916 7984 25968
rect 9404 25916 9456 25968
rect 10508 25916 10560 25968
rect 11796 25993 11805 26027
rect 11805 25993 11839 26027
rect 11839 25993 11848 26027
rect 11796 25984 11848 25993
rect 11888 25984 11940 26036
rect 11152 25959 11204 25968
rect 11152 25925 11161 25959
rect 11161 25925 11195 25959
rect 11195 25925 11204 25959
rect 11152 25916 11204 25925
rect 12532 25959 12584 25968
rect 6184 25780 6236 25832
rect 8576 25780 8628 25832
rect 9128 25823 9180 25832
rect 9128 25789 9137 25823
rect 9137 25789 9171 25823
rect 9171 25789 9180 25823
rect 9128 25780 9180 25789
rect 9864 25780 9916 25832
rect 5816 25712 5868 25764
rect 8208 25712 8260 25764
rect 9220 25712 9272 25764
rect 11152 25712 11204 25764
rect 12532 25925 12541 25959
rect 12541 25925 12575 25959
rect 12575 25925 12584 25959
rect 12532 25916 12584 25925
rect 13452 25916 13504 25968
rect 14372 25916 14424 25968
rect 14464 25916 14516 25968
rect 15292 25959 15344 25968
rect 15292 25925 15301 25959
rect 15301 25925 15335 25959
rect 15335 25925 15344 25959
rect 15292 25916 15344 25925
rect 15752 25916 15804 25968
rect 17316 25984 17368 26036
rect 17500 25984 17552 26036
rect 18696 25984 18748 26036
rect 20720 26027 20772 26036
rect 20720 25993 20729 26027
rect 20729 25993 20763 26027
rect 20763 25993 20772 26027
rect 20720 25984 20772 25993
rect 20996 25984 21048 26036
rect 19340 25916 19392 25968
rect 20076 25916 20128 25968
rect 22744 25984 22796 26036
rect 23204 25984 23256 26036
rect 14648 25848 14700 25900
rect 16212 25848 16264 25900
rect 16856 25848 16908 25900
rect 17132 25891 17184 25900
rect 17132 25857 17141 25891
rect 17141 25857 17175 25891
rect 17175 25857 17184 25891
rect 17132 25848 17184 25857
rect 17960 25891 18012 25900
rect 17960 25857 17969 25891
rect 17969 25857 18003 25891
rect 18003 25857 18012 25891
rect 17960 25848 18012 25857
rect 18144 25848 18196 25900
rect 20628 25891 20680 25900
rect 20628 25857 20637 25891
rect 20637 25857 20671 25891
rect 20671 25857 20680 25891
rect 20628 25848 20680 25857
rect 22836 25848 22888 25900
rect 4620 25644 4672 25696
rect 5540 25644 5592 25696
rect 7196 25687 7248 25696
rect 7196 25653 7205 25687
rect 7205 25653 7239 25687
rect 7239 25653 7248 25687
rect 7196 25644 7248 25653
rect 9772 25644 9824 25696
rect 12164 25712 12216 25764
rect 12716 25644 12768 25696
rect 13452 25712 13504 25764
rect 14464 25712 14516 25764
rect 14740 25712 14792 25764
rect 14648 25644 14700 25696
rect 16028 25712 16080 25764
rect 20076 25780 20128 25832
rect 20168 25823 20220 25832
rect 20168 25789 20177 25823
rect 20177 25789 20211 25823
rect 20211 25789 20220 25823
rect 22652 25823 22704 25832
rect 20168 25780 20220 25789
rect 22652 25789 22661 25823
rect 22661 25789 22695 25823
rect 22695 25789 22704 25823
rect 22652 25780 22704 25789
rect 19340 25712 19392 25764
rect 23572 25712 23624 25764
rect 15384 25644 15436 25696
rect 17408 25644 17460 25696
rect 23112 25644 23164 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 2228 25483 2280 25492
rect 2228 25449 2237 25483
rect 2237 25449 2271 25483
rect 2271 25449 2280 25483
rect 2228 25440 2280 25449
rect 4988 25483 5040 25492
rect 4988 25449 4997 25483
rect 4997 25449 5031 25483
rect 5031 25449 5040 25483
rect 4988 25440 5040 25449
rect 5080 25440 5132 25492
rect 9128 25440 9180 25492
rect 12532 25440 12584 25492
rect 12624 25440 12676 25492
rect 14740 25440 14792 25492
rect 15016 25440 15068 25492
rect 7196 25372 7248 25424
rect 5632 25236 5684 25288
rect 8392 25304 8444 25356
rect 9404 25304 9456 25356
rect 10140 25304 10192 25356
rect 10416 25304 10468 25356
rect 12164 25372 12216 25424
rect 18880 25440 18932 25492
rect 22652 25440 22704 25492
rect 20628 25372 20680 25424
rect 11612 25304 11664 25356
rect 16304 25304 16356 25356
rect 16488 25347 16540 25356
rect 16488 25313 16497 25347
rect 16497 25313 16531 25347
rect 16531 25313 16540 25347
rect 16488 25304 16540 25313
rect 16764 25347 16816 25356
rect 16764 25313 16773 25347
rect 16773 25313 16807 25347
rect 16807 25313 16816 25347
rect 16764 25304 16816 25313
rect 18420 25304 18472 25356
rect 19524 25304 19576 25356
rect 14280 25236 14332 25288
rect 19156 25236 19208 25288
rect 19340 25236 19392 25288
rect 22100 25279 22152 25288
rect 22100 25245 22109 25279
rect 22109 25245 22143 25279
rect 22143 25245 22152 25279
rect 22100 25236 22152 25245
rect 37832 25236 37884 25288
rect 2872 25168 2924 25220
rect 8484 25168 8536 25220
rect 3424 25143 3476 25152
rect 3424 25109 3433 25143
rect 3433 25109 3467 25143
rect 3467 25109 3476 25143
rect 3424 25100 3476 25109
rect 4620 25100 4672 25152
rect 6184 25143 6236 25152
rect 6184 25109 6193 25143
rect 6193 25109 6227 25143
rect 6227 25109 6236 25143
rect 6184 25100 6236 25109
rect 6736 25100 6788 25152
rect 10600 25100 10652 25152
rect 11796 25168 11848 25220
rect 12072 25100 12124 25152
rect 12440 25168 12492 25220
rect 13728 25211 13780 25220
rect 13728 25177 13737 25211
rect 13737 25177 13771 25211
rect 13771 25177 13780 25211
rect 13728 25168 13780 25177
rect 12256 25100 12308 25152
rect 12624 25100 12676 25152
rect 12716 25100 12768 25152
rect 15016 25168 15068 25220
rect 15384 25211 15436 25220
rect 15384 25177 15393 25211
rect 15393 25177 15427 25211
rect 15427 25177 15436 25211
rect 15384 25168 15436 25177
rect 14464 25143 14516 25152
rect 14464 25109 14473 25143
rect 14473 25109 14507 25143
rect 14507 25109 14516 25143
rect 14464 25100 14516 25109
rect 16672 25168 16724 25220
rect 18512 25211 18564 25220
rect 18512 25177 18521 25211
rect 18521 25177 18555 25211
rect 18555 25177 18564 25211
rect 18512 25168 18564 25177
rect 20260 25211 20312 25220
rect 20260 25177 20269 25211
rect 20269 25177 20303 25211
rect 20303 25177 20312 25211
rect 20260 25168 20312 25177
rect 19248 25100 19300 25152
rect 22192 25168 22244 25220
rect 23112 25211 23164 25220
rect 23112 25177 23121 25211
rect 23121 25177 23155 25211
rect 23155 25177 23164 25211
rect 24032 25211 24084 25220
rect 23112 25168 23164 25177
rect 24032 25177 24041 25211
rect 24041 25177 24075 25211
rect 24075 25177 24084 25211
rect 24032 25168 24084 25177
rect 32956 25168 33008 25220
rect 38292 25143 38344 25152
rect 38292 25109 38301 25143
rect 38301 25109 38335 25143
rect 38335 25109 38344 25143
rect 38292 25100 38344 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 4988 24896 5040 24948
rect 9864 24939 9916 24948
rect 9864 24905 9873 24939
rect 9873 24905 9907 24939
rect 9907 24905 9916 24939
rect 9864 24896 9916 24905
rect 11612 24896 11664 24948
rect 1584 24803 1636 24812
rect 1584 24769 1593 24803
rect 1593 24769 1627 24803
rect 1627 24769 1636 24803
rect 1584 24760 1636 24769
rect 2872 24803 2924 24812
rect 2872 24769 2881 24803
rect 2881 24769 2915 24803
rect 2915 24769 2924 24803
rect 2872 24760 2924 24769
rect 3332 24760 3384 24812
rect 4896 24760 4948 24812
rect 6460 24760 6512 24812
rect 6736 24760 6788 24812
rect 7840 24803 7892 24812
rect 7840 24769 7849 24803
rect 7849 24769 7883 24803
rect 7883 24769 7892 24803
rect 7840 24760 7892 24769
rect 7932 24803 7984 24812
rect 7932 24769 7941 24803
rect 7941 24769 7975 24803
rect 7975 24769 7984 24803
rect 7932 24760 7984 24769
rect 8668 24760 8720 24812
rect 8852 24760 8904 24812
rect 10508 24828 10560 24880
rect 11888 24871 11940 24880
rect 11888 24837 11897 24871
rect 11897 24837 11931 24871
rect 11931 24837 11940 24871
rect 12164 24896 12216 24948
rect 13912 24896 13964 24948
rect 11888 24828 11940 24837
rect 12624 24828 12676 24880
rect 10324 24760 10376 24812
rect 12532 24760 12584 24812
rect 13820 24760 13872 24812
rect 9312 24692 9364 24744
rect 10048 24692 10100 24744
rect 12164 24692 12216 24744
rect 1952 24624 2004 24676
rect 5632 24624 5684 24676
rect 3424 24556 3476 24608
rect 4620 24556 4672 24608
rect 7932 24556 7984 24608
rect 9496 24556 9548 24608
rect 10600 24624 10652 24676
rect 15936 24896 15988 24948
rect 16488 24896 16540 24948
rect 18512 24896 18564 24948
rect 14372 24828 14424 24880
rect 20168 24896 20220 24948
rect 22744 24939 22796 24948
rect 22744 24905 22753 24939
rect 22753 24905 22787 24939
rect 22787 24905 22796 24939
rect 22744 24896 22796 24905
rect 23112 24896 23164 24948
rect 15660 24760 15712 24812
rect 16396 24760 16448 24812
rect 14372 24735 14424 24744
rect 14372 24701 14381 24735
rect 14381 24701 14415 24735
rect 14415 24701 14424 24735
rect 14372 24692 14424 24701
rect 15568 24692 15620 24744
rect 17592 24803 17644 24812
rect 17592 24769 17601 24803
rect 17601 24769 17635 24803
rect 17635 24769 17644 24803
rect 17592 24760 17644 24769
rect 18144 24760 18196 24812
rect 17316 24692 17368 24744
rect 19892 24760 19944 24812
rect 21272 24803 21324 24812
rect 21272 24769 21281 24803
rect 21281 24769 21315 24803
rect 21315 24769 21324 24803
rect 21272 24760 21324 24769
rect 21364 24803 21416 24812
rect 21364 24769 21373 24803
rect 21373 24769 21407 24803
rect 21407 24769 21416 24803
rect 21364 24760 21416 24769
rect 21548 24760 21600 24812
rect 19432 24692 19484 24744
rect 20260 24692 20312 24744
rect 13912 24624 13964 24676
rect 16304 24624 16356 24676
rect 17224 24624 17276 24676
rect 20076 24624 20128 24676
rect 20720 24667 20772 24676
rect 20720 24633 20729 24667
rect 20729 24633 20763 24667
rect 20763 24633 20772 24667
rect 20720 24624 20772 24633
rect 21916 24692 21968 24744
rect 30012 24692 30064 24744
rect 37924 24692 37976 24744
rect 38292 24735 38344 24744
rect 38292 24701 38301 24735
rect 38301 24701 38335 24735
rect 38335 24701 38344 24735
rect 38292 24692 38344 24701
rect 11796 24556 11848 24608
rect 14188 24556 14240 24608
rect 15568 24556 15620 24608
rect 15752 24556 15804 24608
rect 16212 24599 16264 24608
rect 16212 24565 16221 24599
rect 16221 24565 16255 24599
rect 16255 24565 16264 24599
rect 16212 24556 16264 24565
rect 17592 24556 17644 24608
rect 36544 24556 36596 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 1676 24395 1728 24404
rect 1676 24361 1685 24395
rect 1685 24361 1719 24395
rect 1719 24361 1728 24395
rect 1676 24352 1728 24361
rect 2596 24352 2648 24404
rect 3332 24395 3384 24404
rect 3332 24361 3341 24395
rect 3341 24361 3375 24395
rect 3375 24361 3384 24395
rect 3332 24352 3384 24361
rect 3884 24352 3936 24404
rect 6828 24352 6880 24404
rect 10508 24352 10560 24404
rect 13728 24352 13780 24404
rect 15844 24352 15896 24404
rect 16396 24352 16448 24404
rect 33600 24395 33652 24404
rect 33600 24361 33609 24395
rect 33609 24361 33643 24395
rect 33643 24361 33652 24395
rect 33600 24352 33652 24361
rect 2228 24327 2280 24336
rect 2228 24293 2237 24327
rect 2237 24293 2271 24327
rect 2271 24293 2280 24327
rect 2228 24284 2280 24293
rect 5908 24284 5960 24336
rect 11888 24284 11940 24336
rect 12624 24284 12676 24336
rect 14924 24284 14976 24336
rect 5724 24216 5776 24268
rect 7932 24216 7984 24268
rect 9680 24216 9732 24268
rect 10416 24216 10468 24268
rect 12164 24216 12216 24268
rect 13820 24216 13872 24268
rect 14280 24216 14332 24268
rect 16764 24284 16816 24336
rect 16396 24216 16448 24268
rect 24032 24284 24084 24336
rect 19248 24216 19300 24268
rect 21272 24259 21324 24268
rect 21272 24225 21281 24259
rect 21281 24225 21315 24259
rect 21315 24225 21324 24259
rect 21272 24216 21324 24225
rect 21916 24259 21968 24268
rect 21916 24225 21925 24259
rect 21925 24225 21959 24259
rect 21959 24225 21968 24259
rect 21916 24216 21968 24225
rect 22192 24259 22244 24268
rect 22192 24225 22201 24259
rect 22201 24225 22235 24259
rect 22235 24225 22244 24259
rect 22192 24216 22244 24225
rect 8392 24191 8444 24200
rect 8392 24157 8401 24191
rect 8401 24157 8435 24191
rect 8435 24157 8444 24191
rect 8392 24148 8444 24157
rect 8944 24148 8996 24200
rect 10968 24148 11020 24200
rect 19064 24148 19116 24200
rect 20352 24148 20404 24200
rect 27252 24148 27304 24200
rect 37832 24191 37884 24200
rect 2872 24012 2924 24064
rect 4620 24012 4672 24064
rect 6644 24055 6696 24064
rect 6644 24021 6653 24055
rect 6653 24021 6687 24055
rect 6687 24021 6696 24055
rect 6644 24012 6696 24021
rect 9956 24012 10008 24064
rect 10140 24080 10192 24132
rect 11336 24080 11388 24132
rect 11428 24080 11480 24132
rect 12256 24123 12308 24132
rect 12256 24089 12265 24123
rect 12265 24089 12299 24123
rect 12299 24089 12308 24123
rect 12256 24080 12308 24089
rect 13084 24123 13136 24132
rect 13084 24089 13093 24123
rect 13093 24089 13127 24123
rect 13127 24089 13136 24123
rect 13084 24080 13136 24089
rect 13268 24080 13320 24132
rect 14740 24123 14792 24132
rect 14740 24089 14749 24123
rect 14749 24089 14783 24123
rect 14783 24089 14792 24123
rect 14740 24080 14792 24089
rect 14832 24123 14884 24132
rect 14832 24089 14841 24123
rect 14841 24089 14875 24123
rect 14875 24089 14884 24123
rect 14832 24080 14884 24089
rect 15844 24080 15896 24132
rect 18604 24123 18656 24132
rect 13544 24012 13596 24064
rect 18604 24089 18613 24123
rect 18613 24089 18647 24123
rect 18647 24089 18656 24123
rect 18604 24080 18656 24089
rect 19892 24080 19944 24132
rect 21180 24080 21232 24132
rect 16580 24012 16632 24064
rect 18512 24055 18564 24064
rect 18512 24021 18521 24055
rect 18521 24021 18555 24055
rect 18555 24021 18564 24055
rect 18512 24012 18564 24021
rect 37832 24157 37841 24191
rect 37841 24157 37875 24191
rect 37875 24157 37884 24191
rect 37832 24148 37884 24157
rect 37556 24012 37608 24064
rect 38016 24055 38068 24064
rect 38016 24021 38025 24055
rect 38025 24021 38059 24055
rect 38059 24021 38068 24055
rect 38016 24012 38068 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 2228 23808 2280 23860
rect 3240 23808 3292 23860
rect 3884 23851 3936 23860
rect 3884 23817 3893 23851
rect 3893 23817 3927 23851
rect 3927 23817 3936 23851
rect 3884 23808 3936 23817
rect 5908 23851 5960 23860
rect 5908 23817 5917 23851
rect 5917 23817 5951 23851
rect 5951 23817 5960 23851
rect 5908 23808 5960 23817
rect 10140 23808 10192 23860
rect 6644 23740 6696 23792
rect 1952 23715 2004 23724
rect 1952 23681 1961 23715
rect 1961 23681 1995 23715
rect 1995 23681 2004 23715
rect 1952 23672 2004 23681
rect 3608 23672 3660 23724
rect 8300 23740 8352 23792
rect 10968 23808 11020 23860
rect 12440 23808 12492 23860
rect 9680 23715 9732 23724
rect 9680 23681 9689 23715
rect 9689 23681 9723 23715
rect 9723 23681 9732 23715
rect 9680 23672 9732 23681
rect 14832 23808 14884 23860
rect 18604 23808 18656 23860
rect 21732 23808 21784 23860
rect 26240 23851 26292 23860
rect 26240 23817 26249 23851
rect 26249 23817 26283 23851
rect 26283 23817 26292 23851
rect 26240 23808 26292 23817
rect 27252 23851 27304 23860
rect 27252 23817 27261 23851
rect 27261 23817 27295 23851
rect 27295 23817 27304 23851
rect 27252 23808 27304 23817
rect 30012 23851 30064 23860
rect 30012 23817 30021 23851
rect 30021 23817 30055 23851
rect 30055 23817 30064 23851
rect 30012 23808 30064 23817
rect 12716 23783 12768 23792
rect 12716 23749 12725 23783
rect 12725 23749 12759 23783
rect 12759 23749 12768 23783
rect 12716 23740 12768 23749
rect 13452 23740 13504 23792
rect 13544 23740 13596 23792
rect 15476 23740 15528 23792
rect 16396 23740 16448 23792
rect 17316 23783 17368 23792
rect 17316 23749 17325 23783
rect 17325 23749 17359 23783
rect 17359 23749 17368 23783
rect 17316 23740 17368 23749
rect 18052 23740 18104 23792
rect 20352 23740 20404 23792
rect 10876 23672 10928 23724
rect 11060 23672 11112 23724
rect 11980 23672 12032 23724
rect 20628 23672 20680 23724
rect 37832 23672 37884 23724
rect 38016 23715 38068 23724
rect 38016 23681 38025 23715
rect 38025 23681 38059 23715
rect 38059 23681 38068 23715
rect 38016 23672 38068 23681
rect 5080 23604 5132 23656
rect 8392 23604 8444 23656
rect 9404 23604 9456 23656
rect 12256 23604 12308 23656
rect 12440 23604 12492 23656
rect 13820 23647 13872 23656
rect 13820 23613 13829 23647
rect 13829 23613 13863 23647
rect 13863 23613 13872 23647
rect 13820 23604 13872 23613
rect 15016 23604 15068 23656
rect 16488 23604 16540 23656
rect 5816 23536 5868 23588
rect 10876 23536 10928 23588
rect 11888 23536 11940 23588
rect 14372 23579 14424 23588
rect 14372 23545 14381 23579
rect 14381 23545 14415 23579
rect 14415 23545 14424 23579
rect 14372 23536 14424 23545
rect 17040 23536 17092 23588
rect 17500 23536 17552 23588
rect 1860 23468 1912 23520
rect 4620 23511 4672 23520
rect 4620 23477 4629 23511
rect 4629 23477 4663 23511
rect 4663 23477 4672 23511
rect 4620 23468 4672 23477
rect 11612 23468 11664 23520
rect 11980 23511 12032 23520
rect 11980 23477 11989 23511
rect 11989 23477 12023 23511
rect 12023 23477 12032 23511
rect 11980 23468 12032 23477
rect 12624 23468 12676 23520
rect 15752 23468 15804 23520
rect 17132 23468 17184 23520
rect 21272 23536 21324 23588
rect 20720 23511 20772 23520
rect 20720 23477 20729 23511
rect 20729 23477 20763 23511
rect 20763 23477 20772 23511
rect 20720 23468 20772 23477
rect 38200 23511 38252 23520
rect 38200 23477 38209 23511
rect 38209 23477 38243 23511
rect 38243 23477 38252 23511
rect 38200 23468 38252 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 1676 23307 1728 23316
rect 1676 23273 1685 23307
rect 1685 23273 1719 23307
rect 1719 23273 1728 23307
rect 1676 23264 1728 23273
rect 2412 23264 2464 23316
rect 3240 23307 3292 23316
rect 3240 23273 3249 23307
rect 3249 23273 3283 23307
rect 3283 23273 3292 23307
rect 3240 23264 3292 23273
rect 8300 23264 8352 23316
rect 8484 23307 8536 23316
rect 8484 23273 8493 23307
rect 8493 23273 8527 23307
rect 8527 23273 8536 23307
rect 8484 23264 8536 23273
rect 11244 23264 11296 23316
rect 14740 23264 14792 23316
rect 15292 23264 15344 23316
rect 16856 23264 16908 23316
rect 17776 23264 17828 23316
rect 18052 23307 18104 23316
rect 18052 23273 18061 23307
rect 18061 23273 18095 23307
rect 18095 23273 18104 23307
rect 18052 23264 18104 23273
rect 19156 23264 19208 23316
rect 19984 23264 20036 23316
rect 3792 22992 3844 23044
rect 10876 23196 10928 23248
rect 12808 23196 12860 23248
rect 8852 23128 8904 23180
rect 9404 23171 9456 23180
rect 9404 23137 9413 23171
rect 9413 23137 9447 23171
rect 9447 23137 9456 23171
rect 9404 23128 9456 23137
rect 10048 23128 10100 23180
rect 11520 23128 11572 23180
rect 11888 23128 11940 23180
rect 13820 23128 13872 23180
rect 14556 23196 14608 23248
rect 17868 23196 17920 23248
rect 16028 23128 16080 23180
rect 13452 23103 13504 23112
rect 6368 22992 6420 23044
rect 13452 23069 13461 23103
rect 13461 23069 13495 23103
rect 13495 23069 13504 23103
rect 13452 23060 13504 23069
rect 15568 23060 15620 23112
rect 17224 23128 17276 23180
rect 8668 22992 8720 23044
rect 11796 23035 11848 23044
rect 3424 22924 3476 22976
rect 4620 22924 4672 22976
rect 5540 22967 5592 22976
rect 5540 22933 5549 22967
rect 5549 22933 5583 22967
rect 5583 22933 5592 22967
rect 5540 22924 5592 22933
rect 7564 22967 7616 22976
rect 7564 22933 7573 22967
rect 7573 22933 7607 22967
rect 7607 22933 7616 22967
rect 7564 22924 7616 22933
rect 9864 22924 9916 22976
rect 11796 23001 11805 23035
rect 11805 23001 11839 23035
rect 11839 23001 11848 23035
rect 11796 22992 11848 23001
rect 10784 22924 10836 22976
rect 13912 22992 13964 23044
rect 15016 23035 15068 23044
rect 12624 22924 12676 22976
rect 15016 23001 15025 23035
rect 15025 23001 15059 23035
rect 15059 23001 15068 23035
rect 15016 22992 15068 23001
rect 14556 22924 14608 22976
rect 16764 23060 16816 23112
rect 17776 23060 17828 23112
rect 18236 23060 18288 23112
rect 18972 23060 19024 23112
rect 19340 23060 19392 23112
rect 20720 23060 20772 23112
rect 20904 23103 20956 23112
rect 20904 23069 20913 23103
rect 20913 23069 20947 23103
rect 20947 23069 20956 23103
rect 20904 23060 20956 23069
rect 16120 22992 16172 23044
rect 17684 22992 17736 23044
rect 31760 23128 31812 23180
rect 22928 23060 22980 23112
rect 18420 22924 18472 22976
rect 18604 22924 18656 22976
rect 20076 22967 20128 22976
rect 20076 22933 20085 22967
rect 20085 22933 20119 22967
rect 20119 22933 20128 22967
rect 20076 22924 20128 22933
rect 38016 22924 38068 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 3792 22763 3844 22772
rect 3792 22729 3801 22763
rect 3801 22729 3835 22763
rect 3835 22729 3844 22763
rect 3792 22720 3844 22729
rect 4068 22720 4120 22772
rect 5448 22763 5500 22772
rect 5448 22729 5457 22763
rect 5457 22729 5491 22763
rect 5491 22729 5500 22763
rect 5448 22720 5500 22729
rect 8668 22763 8720 22772
rect 8668 22729 8677 22763
rect 8677 22729 8711 22763
rect 8711 22729 8720 22763
rect 8668 22720 8720 22729
rect 12532 22720 12584 22772
rect 12716 22720 12768 22772
rect 13268 22720 13320 22772
rect 13452 22720 13504 22772
rect 6000 22652 6052 22704
rect 11612 22652 11664 22704
rect 12164 22652 12216 22704
rect 15200 22720 15252 22772
rect 18052 22763 18104 22772
rect 18052 22729 18061 22763
rect 18061 22729 18095 22763
rect 18095 22729 18104 22763
rect 18052 22720 18104 22729
rect 8576 22627 8628 22636
rect 1952 22516 2004 22568
rect 8576 22593 8585 22627
rect 8585 22593 8619 22627
rect 8619 22593 8628 22627
rect 8576 22584 8628 22593
rect 9404 22627 9456 22636
rect 9404 22593 9413 22627
rect 9413 22593 9447 22627
rect 9447 22593 9456 22627
rect 9404 22584 9456 22593
rect 10876 22584 10928 22636
rect 9680 22516 9732 22568
rect 10692 22559 10744 22568
rect 1676 22491 1728 22500
rect 1676 22457 1685 22491
rect 1685 22457 1719 22491
rect 1719 22457 1728 22491
rect 1676 22448 1728 22457
rect 2044 22448 2096 22500
rect 10692 22525 10701 22559
rect 10701 22525 10735 22559
rect 10735 22525 10744 22559
rect 10692 22516 10744 22525
rect 11888 22516 11940 22568
rect 5540 22380 5592 22432
rect 6460 22380 6512 22432
rect 11060 22423 11112 22432
rect 11060 22389 11069 22423
rect 11069 22389 11103 22423
rect 11103 22389 11112 22423
rect 11060 22380 11112 22389
rect 12256 22448 12308 22500
rect 14924 22695 14976 22704
rect 14924 22661 14933 22695
rect 14933 22661 14967 22695
rect 14967 22661 14976 22695
rect 14924 22652 14976 22661
rect 16304 22652 16356 22704
rect 22192 22720 22244 22772
rect 20168 22695 20220 22704
rect 20168 22661 20177 22695
rect 20177 22661 20211 22695
rect 20211 22661 20220 22695
rect 20168 22652 20220 22661
rect 16028 22584 16080 22636
rect 17592 22627 17644 22636
rect 17592 22593 17601 22627
rect 17601 22593 17635 22627
rect 17635 22593 17644 22627
rect 17592 22584 17644 22593
rect 15384 22516 15436 22568
rect 16856 22516 16908 22568
rect 18328 22516 18380 22568
rect 20076 22559 20128 22568
rect 20076 22525 20085 22559
rect 20085 22525 20119 22559
rect 20119 22525 20128 22559
rect 20076 22516 20128 22525
rect 20352 22516 20404 22568
rect 20812 22652 20864 22704
rect 14556 22448 14608 22500
rect 12900 22380 12952 22432
rect 15292 22380 15344 22432
rect 23572 22380 23624 22432
rect 37832 22380 37884 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 2412 22219 2464 22228
rect 2412 22185 2421 22219
rect 2421 22185 2455 22219
rect 2455 22185 2464 22219
rect 2412 22176 2464 22185
rect 12440 22176 12492 22228
rect 15568 22176 15620 22228
rect 20444 22176 20496 22228
rect 6460 22151 6512 22160
rect 6460 22117 6469 22151
rect 6469 22117 6503 22151
rect 6503 22117 6512 22151
rect 6460 22108 6512 22117
rect 11244 22108 11296 22160
rect 12624 22108 12676 22160
rect 1768 22040 1820 22092
rect 2964 21972 3016 22024
rect 13636 22083 13688 22092
rect 9772 22015 9824 22024
rect 9772 21981 9781 22015
rect 9781 21981 9815 22015
rect 9815 21981 9824 22015
rect 9772 21972 9824 21981
rect 10140 21972 10192 22024
rect 10324 22015 10376 22024
rect 4804 21904 4856 21956
rect 10324 21981 10333 22015
rect 10333 21981 10367 22015
rect 10367 21981 10376 22015
rect 10324 21972 10376 21981
rect 13636 22049 13645 22083
rect 13645 22049 13679 22083
rect 13679 22049 13688 22083
rect 13636 22040 13688 22049
rect 14556 22015 14608 22024
rect 14556 21981 14565 22015
rect 14565 21981 14599 22015
rect 14599 21981 14608 22015
rect 14556 21972 14608 21981
rect 15384 21972 15436 22024
rect 16212 21972 16264 22024
rect 4068 21879 4120 21888
rect 4068 21845 4077 21879
rect 4077 21845 4111 21879
rect 4111 21845 4120 21879
rect 4068 21836 4120 21845
rect 5264 21879 5316 21888
rect 5264 21845 5273 21879
rect 5273 21845 5307 21879
rect 5307 21845 5316 21879
rect 5264 21836 5316 21845
rect 8208 21836 8260 21888
rect 10968 21836 11020 21888
rect 11152 21947 11204 21956
rect 11152 21913 11161 21947
rect 11161 21913 11195 21947
rect 11195 21913 11204 21947
rect 12992 21947 13044 21956
rect 11152 21904 11204 21913
rect 12992 21913 13001 21947
rect 13001 21913 13035 21947
rect 13035 21913 13044 21947
rect 12992 21904 13044 21913
rect 15936 21947 15988 21956
rect 11796 21836 11848 21888
rect 11980 21836 12032 21888
rect 15936 21913 15945 21947
rect 15945 21913 15979 21947
rect 15979 21913 15988 21947
rect 15936 21904 15988 21913
rect 18328 22040 18380 22092
rect 20352 22040 20404 22092
rect 21180 22083 21232 22092
rect 21180 22049 21189 22083
rect 21189 22049 21223 22083
rect 21223 22049 21232 22083
rect 21180 22040 21232 22049
rect 17132 22015 17184 22024
rect 17132 21981 17141 22015
rect 17141 21981 17175 22015
rect 17175 21981 17184 22015
rect 17132 21972 17184 21981
rect 18972 21972 19024 22024
rect 37832 21972 37884 22024
rect 15384 21836 15436 21888
rect 16028 21879 16080 21888
rect 16028 21845 16037 21879
rect 16037 21845 16071 21879
rect 16071 21845 16080 21879
rect 16028 21836 16080 21845
rect 17040 21879 17092 21888
rect 17040 21845 17049 21879
rect 17049 21845 17083 21879
rect 17083 21845 17092 21879
rect 17040 21836 17092 21845
rect 17224 21904 17276 21956
rect 19432 21879 19484 21888
rect 19432 21845 19441 21879
rect 19441 21845 19475 21879
rect 19475 21845 19484 21879
rect 19432 21836 19484 21845
rect 19984 21879 20036 21888
rect 19984 21845 19993 21879
rect 19993 21845 20027 21879
rect 20027 21845 20036 21879
rect 19984 21836 20036 21845
rect 37372 21836 37424 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 2504 21675 2556 21684
rect 2504 21641 2513 21675
rect 2513 21641 2547 21675
rect 2547 21641 2556 21675
rect 2504 21632 2556 21641
rect 3424 21632 3476 21684
rect 3608 21675 3660 21684
rect 3608 21641 3617 21675
rect 3617 21641 3651 21675
rect 3651 21641 3660 21675
rect 3608 21632 3660 21641
rect 4068 21632 4120 21684
rect 6460 21632 6512 21684
rect 9680 21632 9732 21684
rect 9772 21632 9824 21684
rect 5172 21607 5224 21616
rect 5172 21573 5181 21607
rect 5181 21573 5215 21607
rect 5215 21573 5224 21607
rect 5172 21564 5224 21573
rect 10692 21564 10744 21616
rect 10968 21607 11020 21616
rect 10968 21573 10977 21607
rect 10977 21573 11011 21607
rect 11011 21573 11020 21607
rect 10968 21564 11020 21573
rect 17040 21632 17092 21684
rect 18328 21675 18380 21684
rect 18328 21641 18337 21675
rect 18337 21641 18371 21675
rect 18371 21641 18380 21675
rect 18328 21632 18380 21641
rect 20168 21632 20220 21684
rect 15476 21564 15528 21616
rect 1860 21539 1912 21548
rect 1860 21505 1869 21539
rect 1869 21505 1903 21539
rect 1903 21505 1912 21539
rect 1860 21496 1912 21505
rect 1952 21428 2004 21480
rect 8576 21496 8628 21548
rect 9404 21539 9456 21548
rect 9404 21505 9413 21539
rect 9413 21505 9447 21539
rect 9447 21505 9456 21539
rect 9404 21496 9456 21505
rect 17960 21564 18012 21616
rect 9680 21428 9732 21480
rect 10232 21428 10284 21480
rect 11060 21471 11112 21480
rect 11060 21437 11069 21471
rect 11069 21437 11103 21471
rect 11103 21437 11112 21471
rect 11060 21428 11112 21437
rect 11980 21428 12032 21480
rect 11244 21360 11296 21412
rect 12440 21428 12492 21480
rect 12808 21403 12860 21412
rect 12808 21369 12817 21403
rect 12817 21369 12851 21403
rect 12851 21369 12860 21403
rect 12808 21360 12860 21369
rect 14280 21428 14332 21480
rect 15016 21471 15068 21480
rect 15016 21437 15025 21471
rect 15025 21437 15059 21471
rect 15059 21437 15068 21471
rect 15016 21428 15068 21437
rect 15660 21471 15712 21480
rect 15660 21437 15669 21471
rect 15669 21437 15703 21471
rect 15703 21437 15712 21471
rect 15660 21428 15712 21437
rect 17684 21496 17736 21548
rect 21456 21564 21508 21616
rect 19064 21496 19116 21548
rect 38016 21539 38068 21548
rect 38016 21505 38025 21539
rect 38025 21505 38059 21539
rect 38059 21505 38068 21539
rect 38016 21496 38068 21505
rect 16028 21428 16080 21480
rect 26516 21428 26568 21480
rect 17592 21360 17644 21412
rect 17960 21360 18012 21412
rect 18972 21360 19024 21412
rect 1676 21335 1728 21344
rect 1676 21301 1685 21335
rect 1685 21301 1719 21335
rect 1719 21301 1728 21335
rect 1676 21292 1728 21301
rect 10324 21292 10376 21344
rect 15936 21292 15988 21344
rect 17684 21335 17736 21344
rect 17684 21301 17693 21335
rect 17693 21301 17727 21335
rect 17727 21301 17736 21335
rect 17684 21292 17736 21301
rect 38200 21335 38252 21344
rect 38200 21301 38209 21335
rect 38209 21301 38243 21335
rect 38243 21301 38252 21335
rect 38200 21292 38252 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 2228 21131 2280 21140
rect 2228 21097 2237 21131
rect 2237 21097 2271 21131
rect 2271 21097 2280 21131
rect 2228 21088 2280 21097
rect 3056 21088 3108 21140
rect 4068 21131 4120 21140
rect 4068 21097 4077 21131
rect 4077 21097 4111 21131
rect 4111 21097 4120 21131
rect 4068 21088 4120 21097
rect 8116 21088 8168 21140
rect 9496 21088 9548 21140
rect 10784 21088 10836 21140
rect 13268 21088 13320 21140
rect 15568 21088 15620 21140
rect 15936 21088 15988 21140
rect 19984 21088 20036 21140
rect 10232 21063 10284 21072
rect 10232 21029 10241 21063
rect 10241 21029 10275 21063
rect 10275 21029 10284 21063
rect 10232 21020 10284 21029
rect 12808 21020 12860 21072
rect 17500 21020 17552 21072
rect 18236 21020 18288 21072
rect 6920 20952 6972 21004
rect 12440 20952 12492 21004
rect 13084 20952 13136 21004
rect 13728 20995 13780 21004
rect 13728 20961 13737 20995
rect 13737 20961 13771 20995
rect 13771 20961 13780 20995
rect 13728 20952 13780 20961
rect 14372 20952 14424 21004
rect 15660 20952 15712 21004
rect 9496 20927 9548 20936
rect 9496 20893 9505 20927
rect 9505 20893 9539 20927
rect 9539 20893 9548 20927
rect 9496 20884 9548 20893
rect 12900 20884 12952 20936
rect 16856 20927 16908 20936
rect 9956 20748 10008 20800
rect 10784 20859 10836 20868
rect 10784 20825 10793 20859
rect 10793 20825 10827 20859
rect 10827 20825 10836 20859
rect 10784 20816 10836 20825
rect 12624 20816 12676 20868
rect 13176 20859 13228 20868
rect 13176 20825 13185 20859
rect 13185 20825 13219 20859
rect 13219 20825 13228 20859
rect 13176 20816 13228 20825
rect 16856 20893 16865 20927
rect 16865 20893 16899 20927
rect 16899 20893 16908 20927
rect 16856 20884 16908 20893
rect 17500 20927 17552 20936
rect 17500 20893 17509 20927
rect 17509 20893 17543 20927
rect 17543 20893 17552 20927
rect 17500 20884 17552 20893
rect 18880 20884 18932 20936
rect 11980 20748 12032 20800
rect 16212 20748 16264 20800
rect 16948 20816 17000 20868
rect 19064 20816 19116 20868
rect 17316 20791 17368 20800
rect 17316 20757 17325 20791
rect 17325 20757 17359 20791
rect 17359 20757 17368 20791
rect 17316 20748 17368 20757
rect 18696 20791 18748 20800
rect 18696 20757 18705 20791
rect 18705 20757 18739 20791
rect 18739 20757 18748 20791
rect 18696 20748 18748 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 5080 20544 5132 20596
rect 9864 20587 9916 20596
rect 9864 20553 9873 20587
rect 9873 20553 9907 20587
rect 9907 20553 9916 20587
rect 9864 20544 9916 20553
rect 12348 20544 12400 20596
rect 13544 20587 13596 20596
rect 10876 20476 10928 20528
rect 11060 20476 11112 20528
rect 12072 20476 12124 20528
rect 12808 20519 12860 20528
rect 12808 20485 12817 20519
rect 12817 20485 12851 20519
rect 12851 20485 12860 20519
rect 12808 20476 12860 20485
rect 9772 20451 9824 20460
rect 9772 20417 9781 20451
rect 9781 20417 9815 20451
rect 9815 20417 9824 20451
rect 9772 20408 9824 20417
rect 13544 20553 13553 20587
rect 13553 20553 13587 20587
rect 13587 20553 13596 20587
rect 13544 20544 13596 20553
rect 15384 20587 15436 20596
rect 13268 20476 13320 20528
rect 13728 20476 13780 20528
rect 14280 20519 14332 20528
rect 14280 20485 14289 20519
rect 14289 20485 14323 20519
rect 14323 20485 14332 20519
rect 14280 20476 14332 20485
rect 15384 20553 15393 20587
rect 15393 20553 15427 20587
rect 15427 20553 15436 20587
rect 15384 20544 15436 20553
rect 15476 20544 15528 20596
rect 17132 20544 17184 20596
rect 15844 20408 15896 20460
rect 16120 20476 16172 20528
rect 17500 20408 17552 20460
rect 17868 20408 17920 20460
rect 10784 20383 10836 20392
rect 10784 20349 10793 20383
rect 10793 20349 10827 20383
rect 10827 20349 10836 20383
rect 10784 20340 10836 20349
rect 11244 20340 11296 20392
rect 14188 20383 14240 20392
rect 14188 20349 14197 20383
rect 14197 20349 14231 20383
rect 14231 20349 14240 20383
rect 14188 20340 14240 20349
rect 14372 20340 14424 20392
rect 19156 20544 19208 20596
rect 37924 20408 37976 20460
rect 9404 20204 9456 20256
rect 13268 20272 13320 20324
rect 14924 20272 14976 20324
rect 14832 20204 14884 20256
rect 17868 20204 17920 20256
rect 38108 20204 38160 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 9772 20000 9824 20052
rect 11152 20000 11204 20052
rect 9404 19932 9456 19984
rect 13360 19932 13412 19984
rect 13728 20000 13780 20052
rect 16304 20000 16356 20052
rect 17960 20000 18012 20052
rect 21456 20043 21508 20052
rect 21456 20009 21465 20043
rect 21465 20009 21499 20043
rect 21499 20009 21508 20043
rect 21456 20000 21508 20009
rect 23296 19932 23348 19984
rect 11428 19864 11480 19916
rect 12624 19864 12676 19916
rect 14556 19864 14608 19916
rect 16488 19864 16540 19916
rect 16856 19864 16908 19916
rect 7840 19796 7892 19848
rect 10140 19796 10192 19848
rect 10876 19796 10928 19848
rect 15752 19796 15804 19848
rect 21456 19796 21508 19848
rect 11428 19728 11480 19780
rect 13084 19771 13136 19780
rect 1860 19660 1912 19712
rect 13084 19737 13093 19771
rect 13093 19737 13127 19771
rect 13127 19737 13136 19771
rect 13084 19728 13136 19737
rect 13544 19728 13596 19780
rect 14832 19771 14884 19780
rect 13636 19660 13688 19712
rect 14832 19737 14841 19771
rect 14841 19737 14875 19771
rect 14875 19737 14884 19771
rect 14832 19728 14884 19737
rect 15292 19728 15344 19780
rect 17868 19728 17920 19780
rect 37464 19864 37516 19916
rect 36544 19796 36596 19848
rect 16304 19660 16356 19712
rect 33692 19728 33744 19780
rect 36728 19660 36780 19712
rect 38200 19703 38252 19712
rect 38200 19669 38209 19703
rect 38209 19669 38243 19703
rect 38243 19669 38252 19703
rect 38200 19660 38252 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 10876 19456 10928 19508
rect 11060 19499 11112 19508
rect 11060 19465 11069 19499
rect 11069 19465 11103 19499
rect 11103 19465 11112 19499
rect 11060 19456 11112 19465
rect 11980 19499 12032 19508
rect 11980 19465 11989 19499
rect 11989 19465 12023 19499
rect 12023 19465 12032 19499
rect 11980 19456 12032 19465
rect 13544 19499 13596 19508
rect 13544 19465 13553 19499
rect 13553 19465 13587 19499
rect 13587 19465 13596 19499
rect 13544 19456 13596 19465
rect 1860 19363 1912 19372
rect 1860 19329 1869 19363
rect 1869 19329 1903 19363
rect 1903 19329 1912 19363
rect 1860 19320 1912 19329
rect 13728 19388 13780 19440
rect 14188 19431 14240 19440
rect 14188 19397 14197 19431
rect 14197 19397 14231 19431
rect 14231 19397 14240 19431
rect 14188 19388 14240 19397
rect 16304 19456 16356 19508
rect 22744 19456 22796 19508
rect 12624 19363 12676 19372
rect 12624 19329 12633 19363
rect 12633 19329 12667 19363
rect 12667 19329 12676 19363
rect 12624 19320 12676 19329
rect 13636 19363 13688 19372
rect 13636 19329 13645 19363
rect 13645 19329 13679 19363
rect 13679 19329 13688 19363
rect 13636 19320 13688 19329
rect 11428 19252 11480 19304
rect 15016 19252 15068 19304
rect 12992 19184 13044 19236
rect 15752 19320 15804 19372
rect 15292 19184 15344 19236
rect 17224 19320 17276 19372
rect 1676 19159 1728 19168
rect 1676 19125 1685 19159
rect 1685 19125 1719 19159
rect 1719 19125 1728 19159
rect 1676 19116 1728 19125
rect 11336 19116 11388 19168
rect 14648 19116 14700 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 7104 18912 7156 18964
rect 10140 18955 10192 18964
rect 10140 18921 10149 18955
rect 10149 18921 10183 18955
rect 10183 18921 10192 18955
rect 10140 18912 10192 18921
rect 12624 18912 12676 18964
rect 12900 18912 12952 18964
rect 14188 18912 14240 18964
rect 15200 18955 15252 18964
rect 15200 18921 15209 18955
rect 15209 18921 15243 18955
rect 15243 18921 15252 18955
rect 15200 18912 15252 18921
rect 16212 18912 16264 18964
rect 16488 18955 16540 18964
rect 16488 18921 16497 18955
rect 16497 18921 16531 18955
rect 16531 18921 16540 18955
rect 16488 18912 16540 18921
rect 13636 18844 13688 18896
rect 9496 18776 9548 18828
rect 11612 18776 11664 18828
rect 11520 18708 11572 18760
rect 13912 18776 13964 18828
rect 15108 18776 15160 18828
rect 13544 18751 13596 18760
rect 13544 18717 13553 18751
rect 13553 18717 13587 18751
rect 13587 18717 13596 18751
rect 13544 18708 13596 18717
rect 14648 18751 14700 18760
rect 14648 18717 14657 18751
rect 14657 18717 14691 18751
rect 14691 18717 14700 18751
rect 14648 18708 14700 18717
rect 15200 18708 15252 18760
rect 20904 18776 20956 18828
rect 7472 18640 7524 18692
rect 17316 18640 17368 18692
rect 3976 18615 4028 18624
rect 3976 18581 3985 18615
rect 3985 18581 4019 18615
rect 4019 18581 4028 18615
rect 3976 18572 4028 18581
rect 11520 18615 11572 18624
rect 11520 18581 11529 18615
rect 11529 18581 11563 18615
rect 11563 18581 11572 18615
rect 11520 18572 11572 18581
rect 11612 18572 11664 18624
rect 12992 18572 13044 18624
rect 13728 18572 13780 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 7472 18368 7524 18420
rect 12808 18368 12860 18420
rect 13176 18368 13228 18420
rect 14280 18368 14332 18420
rect 15108 18368 15160 18420
rect 9220 18300 9272 18352
rect 13544 18300 13596 18352
rect 15292 18343 15344 18352
rect 15292 18309 15301 18343
rect 15301 18309 15335 18343
rect 15335 18309 15344 18343
rect 15292 18300 15344 18309
rect 10232 18232 10284 18284
rect 5448 18164 5500 18216
rect 13728 18275 13780 18284
rect 13728 18241 13737 18275
rect 13737 18241 13771 18275
rect 13771 18241 13780 18275
rect 13728 18232 13780 18241
rect 13912 18164 13964 18216
rect 1676 18071 1728 18080
rect 1676 18037 1685 18071
rect 1685 18037 1719 18071
rect 1719 18037 1728 18071
rect 1676 18028 1728 18037
rect 3332 18028 3384 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 12992 17867 13044 17876
rect 12992 17833 13001 17867
rect 13001 17833 13035 17867
rect 13035 17833 13044 17867
rect 12992 17824 13044 17833
rect 15200 17824 15252 17876
rect 14832 17731 14884 17740
rect 14832 17697 14841 17731
rect 14841 17697 14875 17731
rect 14875 17697 14884 17731
rect 14832 17688 14884 17697
rect 38016 17620 38068 17672
rect 14556 17552 14608 17604
rect 16488 17484 16540 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 13912 17323 13964 17332
rect 13912 17289 13921 17323
rect 13921 17289 13955 17323
rect 13955 17289 13964 17323
rect 13912 17280 13964 17289
rect 14556 17323 14608 17332
rect 14556 17289 14565 17323
rect 14565 17289 14599 17323
rect 14599 17289 14608 17323
rect 14556 17280 14608 17289
rect 15292 17280 15344 17332
rect 15016 17144 15068 17196
rect 34796 16940 34848 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 18604 16532 18656 16584
rect 24584 16600 24636 16652
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 3976 16056 4028 16108
rect 38108 16056 38160 16108
rect 1676 15895 1728 15904
rect 1676 15861 1685 15895
rect 1685 15861 1719 15895
rect 1719 15861 1728 15895
rect 1676 15852 1728 15861
rect 38200 15895 38252 15904
rect 38200 15861 38209 15895
rect 38209 15861 38243 15895
rect 38243 15861 38252 15895
rect 38200 15852 38252 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 38016 14467 38068 14476
rect 38016 14433 38025 14467
rect 38025 14433 38059 14467
rect 38059 14433 38068 14467
rect 38016 14424 38068 14433
rect 38292 14399 38344 14408
rect 38292 14365 38301 14399
rect 38301 14365 38335 14399
rect 38335 14365 38344 14399
rect 38292 14356 38344 14365
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 38292 14059 38344 14068
rect 38292 14025 38301 14059
rect 38301 14025 38335 14059
rect 38335 14025 38344 14059
rect 38292 14016 38344 14025
rect 5264 13880 5316 13932
rect 1676 13719 1728 13728
rect 1676 13685 1685 13719
rect 1685 13685 1719 13719
rect 1719 13685 1728 13719
rect 1676 13676 1728 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 13268 13515 13320 13524
rect 13268 13481 13277 13515
rect 13277 13481 13311 13515
rect 13311 13481 13320 13515
rect 13268 13472 13320 13481
rect 20444 13515 20496 13524
rect 20444 13481 20453 13515
rect 20453 13481 20487 13515
rect 20487 13481 20496 13515
rect 20444 13472 20496 13481
rect 13452 13268 13504 13320
rect 20444 13268 20496 13320
rect 20076 13132 20128 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 3332 12792 3384 12844
rect 21824 12928 21876 12980
rect 37464 12767 37516 12776
rect 37464 12733 37473 12767
rect 37473 12733 37507 12767
rect 37507 12733 37516 12767
rect 37464 12724 37516 12733
rect 1676 12631 1728 12640
rect 1676 12597 1685 12631
rect 1685 12597 1719 12631
rect 1719 12597 1728 12631
rect 1676 12588 1728 12597
rect 16120 12631 16172 12640
rect 16120 12597 16129 12631
rect 16129 12597 16163 12631
rect 16163 12597 16172 12631
rect 16120 12588 16172 12597
rect 38200 12631 38252 12640
rect 38200 12597 38209 12631
rect 38209 12597 38243 12631
rect 38243 12597 38252 12631
rect 38200 12588 38252 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 16856 12316 16908 12368
rect 15568 12180 15620 12232
rect 38016 12180 38068 12232
rect 38016 12087 38068 12096
rect 38016 12053 38025 12087
rect 38025 12053 38059 12087
rect 38059 12053 38068 12087
rect 38016 12044 38068 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 18788 11840 18840 11892
rect 24952 11704 25004 11756
rect 24952 11543 25004 11552
rect 24952 11509 24961 11543
rect 24961 11509 24995 11543
rect 24995 11509 25004 11543
rect 24952 11500 25004 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 38108 11024 38160 11076
rect 38200 11067 38252 11076
rect 38200 11033 38209 11067
rect 38209 11033 38243 11067
rect 38243 11033 38252 11067
rect 38200 11024 38252 11033
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 13084 10752 13136 10804
rect 18512 10684 18564 10736
rect 1676 10455 1728 10464
rect 1676 10421 1685 10455
rect 1685 10421 1719 10455
rect 1719 10421 1728 10455
rect 1676 10412 1728 10421
rect 13820 10455 13872 10464
rect 13820 10421 13829 10455
rect 13829 10421 13863 10455
rect 13863 10421 13872 10455
rect 13820 10412 13872 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 10048 10208 10100 10260
rect 12716 10251 12768 10260
rect 12716 10217 12725 10251
rect 12725 10217 12759 10251
rect 12759 10217 12768 10251
rect 12716 10208 12768 10217
rect 8576 10004 8628 10056
rect 12716 10004 12768 10056
rect 13268 9911 13320 9920
rect 13268 9877 13277 9911
rect 13277 9877 13311 9911
rect 13311 9877 13320 9911
rect 13268 9868 13320 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 13820 9664 13872 9716
rect 19984 9664 20036 9716
rect 20260 9596 20312 9648
rect 24768 9324 24820 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 38016 8959 38068 8968
rect 38016 8925 38025 8959
rect 38025 8925 38059 8959
rect 38059 8925 38068 8959
rect 38016 8916 38068 8925
rect 1676 8891 1728 8900
rect 1676 8857 1685 8891
rect 1685 8857 1719 8891
rect 1719 8857 1728 8891
rect 1676 8848 1728 8857
rect 17684 8780 17736 8832
rect 38200 8823 38252 8832
rect 38200 8789 38209 8823
rect 38209 8789 38243 8823
rect 38243 8789 38252 8823
rect 38200 8780 38252 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 1676 8619 1728 8628
rect 1676 8585 1685 8619
rect 1685 8585 1719 8619
rect 1719 8585 1728 8619
rect 1676 8576 1728 8585
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 4804 7420 4856 7472
rect 37740 7420 37792 7472
rect 1584 7352 1636 7404
rect 38200 7395 38252 7404
rect 38200 7361 38209 7395
rect 38209 7361 38243 7395
rect 38243 7361 38252 7395
rect 38200 7352 38252 7361
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 1584 6987 1636 6996
rect 1584 6953 1593 6987
rect 1593 6953 1627 6987
rect 1627 6953 1636 6987
rect 1584 6944 1636 6953
rect 9680 6808 9732 6860
rect 24676 6740 24728 6792
rect 2780 6604 2832 6656
rect 25228 6672 25280 6724
rect 24676 6647 24728 6656
rect 24676 6613 24685 6647
rect 24685 6613 24719 6647
rect 24719 6613 24728 6647
rect 24676 6604 24728 6613
rect 38108 6604 38160 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 32956 6443 33008 6452
rect 32956 6409 32965 6443
rect 32965 6409 32999 6443
rect 32999 6409 33008 6443
rect 32956 6400 33008 6409
rect 34520 6128 34572 6180
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 37924 5788 37976 5840
rect 38200 5627 38252 5636
rect 38200 5593 38209 5627
rect 38209 5593 38243 5627
rect 38243 5593 38252 5627
rect 38200 5584 38252 5593
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 1768 5355 1820 5364
rect 1768 5321 1777 5355
rect 1777 5321 1811 5355
rect 1811 5321 1820 5355
rect 1768 5312 1820 5321
rect 1584 5176 1636 5228
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 1584 4811 1636 4820
rect 1584 4777 1593 4811
rect 1593 4777 1627 4811
rect 1627 4777 1636 4811
rect 1584 4768 1636 4777
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 2780 3476 2832 3528
rect 1952 3408 2004 3460
rect 18696 3408 18748 3460
rect 1676 3383 1728 3392
rect 1676 3349 1685 3383
rect 1685 3349 1719 3383
rect 1719 3349 1728 3383
rect 1676 3340 1728 3349
rect 37464 3383 37516 3392
rect 37464 3349 37473 3383
rect 37473 3349 37507 3383
rect 37507 3349 37516 3383
rect 37464 3340 37516 3349
rect 38200 3383 38252 3392
rect 38200 3349 38209 3383
rect 38209 3349 38243 3383
rect 38243 3349 38252 3383
rect 38200 3340 38252 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 5540 3136 5592 3188
rect 7564 3136 7616 3188
rect 34796 3136 34848 3188
rect 1676 3043 1728 3052
rect 1676 3009 1685 3043
rect 1685 3009 1719 3043
rect 1719 3009 1728 3043
rect 1676 3000 1728 3009
rect 8576 3043 8628 3052
rect 8576 3009 8585 3043
rect 8585 3009 8619 3043
rect 8619 3009 8628 3043
rect 8576 3000 8628 3009
rect 12716 3000 12768 3052
rect 13452 3043 13504 3052
rect 13452 3009 13461 3043
rect 13461 3009 13495 3043
rect 13495 3009 13504 3043
rect 13452 3000 13504 3009
rect 19984 3043 20036 3052
rect 19984 3009 19993 3043
rect 19993 3009 20027 3043
rect 20027 3009 20036 3043
rect 19984 3000 20036 3009
rect 33876 3043 33928 3052
rect 33876 3009 33885 3043
rect 33885 3009 33919 3043
rect 33919 3009 33928 3043
rect 33876 3000 33928 3009
rect 34520 3000 34572 3052
rect 37464 2932 37516 2984
rect 11520 2864 11572 2916
rect 27344 2864 27396 2916
rect 35900 2864 35952 2916
rect 2412 2839 2464 2848
rect 2412 2805 2421 2839
rect 2421 2805 2455 2839
rect 2455 2805 2464 2839
rect 2412 2796 2464 2805
rect 8300 2796 8352 2848
rect 29644 2839 29696 2848
rect 29644 2805 29653 2839
rect 29653 2805 29687 2839
rect 29687 2805 29696 2839
rect 29644 2796 29696 2805
rect 36820 2796 36872 2848
rect 37648 2796 37700 2848
rect 38016 2796 38068 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 11888 2635 11940 2644
rect 11888 2601 11897 2635
rect 11897 2601 11931 2635
rect 11931 2601 11940 2635
rect 11888 2592 11940 2601
rect 14464 2592 14516 2644
rect 15200 2567 15252 2576
rect 8576 2456 8628 2508
rect 15200 2533 15209 2567
rect 15209 2533 15243 2567
rect 15243 2533 15252 2567
rect 15200 2524 15252 2533
rect 16488 2592 16540 2644
rect 32404 2635 32456 2644
rect 32404 2601 32413 2635
rect 32413 2601 32447 2635
rect 32447 2601 32456 2635
rect 32404 2592 32456 2601
rect 33692 2635 33744 2644
rect 33692 2601 33701 2635
rect 33701 2601 33735 2635
rect 33735 2601 33744 2635
rect 33692 2592 33744 2601
rect 36728 2635 36780 2644
rect 36728 2601 36737 2635
rect 36737 2601 36771 2635
rect 36771 2601 36780 2635
rect 36728 2592 36780 2601
rect 37556 2635 37608 2644
rect 37556 2601 37565 2635
rect 37565 2601 37599 2635
rect 37599 2601 37608 2635
rect 37556 2592 37608 2601
rect 23296 2567 23348 2576
rect 19984 2456 20036 2508
rect 1952 2388 2004 2440
rect 2412 2363 2464 2372
rect 2412 2329 2421 2363
rect 2421 2329 2455 2363
rect 2455 2329 2464 2363
rect 2412 2320 2464 2329
rect 1308 2252 1360 2304
rect 3240 2252 3292 2304
rect 5540 2431 5592 2440
rect 5540 2397 5549 2431
rect 5549 2397 5583 2431
rect 5583 2397 5592 2431
rect 5540 2388 5592 2397
rect 8300 2431 8352 2440
rect 8300 2397 8309 2431
rect 8309 2397 8343 2431
rect 8343 2397 8352 2431
rect 8300 2388 8352 2397
rect 9680 2388 9732 2440
rect 12716 2388 12768 2440
rect 13268 2431 13320 2440
rect 13268 2397 13277 2431
rect 13277 2397 13311 2431
rect 13311 2397 13320 2431
rect 13268 2388 13320 2397
rect 4528 2252 4580 2304
rect 6460 2252 6512 2304
rect 8392 2252 8444 2304
rect 11612 2320 11664 2372
rect 16120 2388 16172 2440
rect 16856 2431 16908 2440
rect 16856 2397 16865 2431
rect 16865 2397 16899 2431
rect 16899 2397 16908 2431
rect 16856 2388 16908 2397
rect 20076 2431 20128 2440
rect 20076 2397 20085 2431
rect 20085 2397 20119 2431
rect 20119 2397 20128 2431
rect 20076 2388 20128 2397
rect 23296 2533 23305 2567
rect 23305 2533 23339 2567
rect 23339 2533 23348 2567
rect 23296 2524 23348 2533
rect 24952 2456 25004 2508
rect 33876 2456 33928 2508
rect 25228 2431 25280 2440
rect 25228 2397 25237 2431
rect 25237 2397 25271 2431
rect 25271 2397 25280 2431
rect 25228 2388 25280 2397
rect 14832 2320 14884 2372
rect 18052 2320 18104 2372
rect 23204 2320 23256 2372
rect 24768 2320 24820 2372
rect 27344 2388 27396 2440
rect 29644 2388 29696 2440
rect 34796 2388 34848 2440
rect 35900 2431 35952 2440
rect 35900 2397 35909 2431
rect 35909 2397 35943 2431
rect 35943 2397 35952 2431
rect 35900 2388 35952 2397
rect 37280 2388 37332 2440
rect 33508 2320 33560 2372
rect 36820 2363 36872 2372
rect 36820 2329 36829 2363
rect 36829 2329 36863 2363
rect 36863 2329 36872 2363
rect 36820 2320 36872 2329
rect 12900 2252 12952 2304
rect 16764 2252 16816 2304
rect 19984 2252 20036 2304
rect 21640 2252 21692 2304
rect 25136 2252 25188 2304
rect 26424 2252 26476 2304
rect 28356 2252 28408 2304
rect 31760 2295 31812 2304
rect 31760 2261 31769 2295
rect 31769 2261 31803 2295
rect 31803 2261 31812 2295
rect 31760 2252 31812 2261
rect 34796 2252 34848 2304
rect 35808 2252 35860 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 20 1300 72 1352
rect 2412 1300 2464 1352
<< metal2 >>
rect 18 39200 74 39800
rect 1950 39200 2006 39800
rect 3882 39200 3938 39800
rect 5170 39200 5226 39800
rect 7102 39200 7158 39800
rect 8390 39200 8446 39800
rect 10322 39200 10378 39800
rect 12254 39200 12310 39800
rect 13542 39200 13598 39800
rect 13648 39222 13860 39250
rect 32 37670 60 39200
rect 20 37664 72 37670
rect 20 37606 72 37612
rect 1584 36848 1636 36854
rect 1584 36790 1636 36796
rect 1308 36712 1360 36718
rect 1308 36654 1360 36660
rect 1320 26042 1348 36654
rect 1596 33862 1624 36790
rect 1676 36780 1728 36786
rect 1676 36722 1728 36728
rect 1688 36242 1716 36722
rect 1676 36236 1728 36242
rect 1676 36178 1728 36184
rect 1688 35154 1716 36178
rect 1768 36032 1820 36038
rect 1768 35974 1820 35980
rect 1676 35148 1728 35154
rect 1676 35090 1728 35096
rect 1688 34610 1716 35090
rect 1676 34604 1728 34610
rect 1676 34546 1728 34552
rect 1584 33856 1636 33862
rect 1584 33798 1636 33804
rect 1596 30841 1624 33798
rect 1780 33114 1808 35974
rect 1964 35698 1992 39200
rect 2410 38856 2466 38865
rect 2410 38791 2466 38800
rect 2044 37256 2096 37262
rect 2044 37198 2096 37204
rect 1952 35692 2004 35698
rect 1952 35634 2004 35640
rect 1860 35556 1912 35562
rect 1860 35498 1912 35504
rect 1952 35556 2004 35562
rect 1952 35498 2004 35504
rect 1872 33658 1900 35498
rect 1964 35018 1992 35498
rect 1952 35012 2004 35018
rect 1952 34954 2004 34960
rect 1860 33652 1912 33658
rect 1860 33594 1912 33600
rect 1964 33454 1992 34954
rect 1952 33448 2004 33454
rect 1952 33390 2004 33396
rect 1768 33108 1820 33114
rect 1768 33050 1820 33056
rect 1768 32224 1820 32230
rect 1768 32166 1820 32172
rect 1676 31476 1728 31482
rect 1676 31418 1728 31424
rect 1688 31385 1716 31418
rect 1674 31376 1730 31385
rect 1674 31311 1730 31320
rect 1582 30832 1638 30841
rect 1582 30767 1638 30776
rect 1676 30592 1728 30598
rect 1676 30534 1728 30540
rect 1688 30025 1716 30534
rect 1674 30016 1730 30025
rect 1674 29951 1730 29960
rect 1780 29850 1808 32166
rect 1952 30728 2004 30734
rect 1952 30670 2004 30676
rect 1860 30592 1912 30598
rect 1860 30534 1912 30540
rect 1768 29844 1820 29850
rect 1768 29786 1820 29792
rect 1676 29504 1728 29510
rect 1676 29446 1728 29452
rect 1688 29306 1716 29446
rect 1676 29300 1728 29306
rect 1676 29242 1728 29248
rect 1872 29170 1900 30534
rect 1860 29164 1912 29170
rect 1860 29106 1912 29112
rect 1676 28416 1728 28422
rect 1676 28358 1728 28364
rect 1688 27470 1716 28358
rect 1768 28076 1820 28082
rect 1768 28018 1820 28024
rect 1780 27985 1808 28018
rect 1766 27976 1822 27985
rect 1766 27911 1822 27920
rect 1676 27464 1728 27470
rect 1676 27406 1728 27412
rect 1676 26784 1728 26790
rect 1676 26726 1728 26732
rect 1688 26625 1716 26726
rect 1674 26616 1730 26625
rect 1674 26551 1730 26560
rect 1308 26036 1360 26042
rect 1308 25978 1360 25984
rect 1584 24812 1636 24818
rect 1584 24754 1636 24760
rect 1596 24585 1624 24754
rect 1582 24576 1638 24585
rect 1582 24511 1638 24520
rect 1676 24404 1728 24410
rect 1676 24346 1728 24352
rect 1688 23322 1716 24346
rect 1676 23316 1728 23322
rect 1676 23258 1728 23264
rect 1674 22536 1730 22545
rect 1674 22471 1676 22480
rect 1728 22471 1730 22480
rect 1676 22442 1728 22448
rect 1780 22098 1808 27911
rect 1964 24834 1992 30670
rect 2056 26586 2084 37198
rect 2136 33924 2188 33930
rect 2136 33866 2188 33872
rect 2148 26586 2176 33866
rect 2228 33312 2280 33318
rect 2228 33254 2280 33260
rect 2240 27130 2268 33254
rect 2424 31754 2452 38791
rect 3896 37330 3924 39200
rect 4804 37800 4856 37806
rect 4804 37742 4856 37748
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4816 37330 4844 37742
rect 4896 37664 4948 37670
rect 4896 37606 4948 37612
rect 3148 37324 3200 37330
rect 3148 37266 3200 37272
rect 3884 37324 3936 37330
rect 3884 37266 3936 37272
rect 4804 37324 4856 37330
rect 4804 37266 4856 37272
rect 3160 37210 3188 37266
rect 3160 37182 3372 37210
rect 2870 36816 2926 36825
rect 2870 36751 2926 36760
rect 2504 36100 2556 36106
rect 2504 36042 2556 36048
rect 2332 31726 2452 31754
rect 2332 31346 2360 31726
rect 2320 31340 2372 31346
rect 2320 31282 2372 31288
rect 2228 27124 2280 27130
rect 2228 27066 2280 27072
rect 2044 26580 2096 26586
rect 2044 26522 2096 26528
rect 2136 26580 2188 26586
rect 2136 26522 2188 26528
rect 2228 26376 2280 26382
rect 2228 26318 2280 26324
rect 2240 25498 2268 26318
rect 2228 25492 2280 25498
rect 2228 25434 2280 25440
rect 1964 24806 2084 24834
rect 1952 24676 2004 24682
rect 1952 24618 2004 24624
rect 1964 23730 1992 24618
rect 1952 23724 2004 23730
rect 1952 23666 2004 23672
rect 1860 23520 1912 23526
rect 1860 23462 1912 23468
rect 1768 22092 1820 22098
rect 1768 22034 1820 22040
rect 1872 21554 1900 23462
rect 1952 22568 2004 22574
rect 1952 22510 2004 22516
rect 1860 21548 1912 21554
rect 1860 21490 1912 21496
rect 1964 21486 1992 22510
rect 2056 22506 2084 24806
rect 2240 24342 2268 25434
rect 2228 24336 2280 24342
rect 2228 24278 2280 24284
rect 2240 23866 2268 24278
rect 2228 23860 2280 23866
rect 2228 23802 2280 23808
rect 2044 22500 2096 22506
rect 2044 22442 2096 22448
rect 2332 22094 2360 31282
rect 2412 30592 2464 30598
rect 2412 30534 2464 30540
rect 2424 30258 2452 30534
rect 2412 30252 2464 30258
rect 2412 30194 2464 30200
rect 2412 29708 2464 29714
rect 2412 29650 2464 29656
rect 2424 29617 2452 29650
rect 2410 29608 2466 29617
rect 2410 29543 2466 29552
rect 2412 29164 2464 29170
rect 2412 29106 2464 29112
rect 2424 28558 2452 29106
rect 2412 28552 2464 28558
rect 2412 28494 2464 28500
rect 2424 28014 2452 28494
rect 2412 28008 2464 28014
rect 2412 27950 2464 27956
rect 2516 26042 2544 36042
rect 2884 35766 2912 36751
rect 3344 36582 3372 37182
rect 3700 36848 3752 36854
rect 3700 36790 3752 36796
rect 3332 36576 3384 36582
rect 3332 36518 3384 36524
rect 2872 35760 2924 35766
rect 2872 35702 2924 35708
rect 2780 35692 2832 35698
rect 2780 35634 2832 35640
rect 2688 33584 2740 33590
rect 2686 33552 2688 33561
rect 2740 33552 2742 33561
rect 2686 33487 2742 33496
rect 2596 32836 2648 32842
rect 2596 32778 2648 32784
rect 2608 28422 2636 32778
rect 2688 32496 2740 32502
rect 2688 32438 2740 32444
rect 2596 28416 2648 28422
rect 2596 28358 2648 28364
rect 2596 28008 2648 28014
rect 2596 27950 2648 27956
rect 2608 26314 2636 27950
rect 2700 27538 2728 32438
rect 2792 31822 2820 35634
rect 2872 35624 2924 35630
rect 2872 35566 2924 35572
rect 2780 31816 2832 31822
rect 2780 31758 2832 31764
rect 2884 31754 2912 35566
rect 3240 33448 3292 33454
rect 3240 33390 3292 33396
rect 3252 33289 3280 33390
rect 3238 33280 3294 33289
rect 3238 33215 3294 33224
rect 3344 33130 3372 36518
rect 3516 36100 3568 36106
rect 3252 33102 3372 33130
rect 3436 36060 3516 36088
rect 3054 32464 3110 32473
rect 3054 32399 3110 32408
rect 3068 31890 3096 32399
rect 3056 31884 3108 31890
rect 3056 31826 3108 31832
rect 3148 31816 3200 31822
rect 3148 31758 3200 31764
rect 2884 31726 3004 31754
rect 2780 31272 2832 31278
rect 2780 31214 2832 31220
rect 2792 29102 2820 31214
rect 2872 30728 2924 30734
rect 2872 30670 2924 30676
rect 2780 29096 2832 29102
rect 2780 29038 2832 29044
rect 2780 28416 2832 28422
rect 2780 28358 2832 28364
rect 2792 28218 2820 28358
rect 2780 28212 2832 28218
rect 2780 28154 2832 28160
rect 2884 28014 2912 30670
rect 2872 28008 2924 28014
rect 2872 27950 2924 27956
rect 2688 27532 2740 27538
rect 2688 27474 2740 27480
rect 2688 27396 2740 27402
rect 2688 27338 2740 27344
rect 2700 26382 2728 27338
rect 2884 26994 2912 27950
rect 2872 26988 2924 26994
rect 2872 26930 2924 26936
rect 2884 26382 2912 26930
rect 2688 26376 2740 26382
rect 2688 26318 2740 26324
rect 2872 26376 2924 26382
rect 2872 26318 2924 26324
rect 2596 26308 2648 26314
rect 2596 26250 2648 26256
rect 2504 26036 2556 26042
rect 2504 25978 2556 25984
rect 2608 24410 2636 26250
rect 2884 25906 2912 26318
rect 2872 25900 2924 25906
rect 2872 25842 2924 25848
rect 2884 25226 2912 25842
rect 2872 25220 2924 25226
rect 2872 25162 2924 25168
rect 2884 24818 2912 25162
rect 2872 24812 2924 24818
rect 2872 24754 2924 24760
rect 2596 24404 2648 24410
rect 2596 24346 2648 24352
rect 2884 24070 2912 24754
rect 2872 24064 2924 24070
rect 2872 24006 2924 24012
rect 2412 23316 2464 23322
rect 2412 23258 2464 23264
rect 2424 22234 2452 23258
rect 2412 22228 2464 22234
rect 2412 22170 2464 22176
rect 2240 22066 2360 22094
rect 2424 22094 2452 22170
rect 2424 22066 2544 22094
rect 1952 21480 2004 21486
rect 1952 21422 2004 21428
rect 1676 21344 1728 21350
rect 1676 21286 1728 21292
rect 1688 21185 1716 21286
rect 1674 21176 1730 21185
rect 1674 21111 1730 21120
rect 1860 19712 1912 19718
rect 1860 19654 1912 19660
rect 1872 19378 1900 19654
rect 1860 19372 1912 19378
rect 1860 19314 1912 19320
rect 1676 19168 1728 19174
rect 1674 19136 1676 19145
rect 1728 19136 1730 19145
rect 1674 19071 1730 19080
rect 1676 18080 1728 18086
rect 1676 18022 1728 18028
rect 1688 17785 1716 18022
rect 1674 17776 1730 17785
rect 1674 17711 1730 17720
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 1688 15745 1716 15846
rect 1674 15736 1730 15745
rect 1674 15671 1730 15680
rect 1676 13728 1728 13734
rect 1674 13696 1676 13705
rect 1728 13696 1730 13705
rect 1674 13631 1730 13640
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 1688 12345 1716 12582
rect 1674 12336 1730 12345
rect 1674 12271 1730 12280
rect 1676 10464 1728 10470
rect 1676 10406 1728 10412
rect 1688 10305 1716 10406
rect 1674 10296 1730 10305
rect 1674 10231 1730 10240
rect 1674 8936 1730 8945
rect 1674 8871 1676 8880
rect 1728 8871 1730 8880
rect 1676 8842 1728 8848
rect 1688 8634 1716 8842
rect 1676 8628 1728 8634
rect 1676 8570 1728 8576
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 1596 7002 1624 7346
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1596 6905 1624 6938
rect 1964 6914 1992 21422
rect 2240 21146 2268 22066
rect 2516 21690 2544 22066
rect 2976 22030 3004 31726
rect 3056 29640 3108 29646
rect 3056 29582 3108 29588
rect 3068 27606 3096 29582
rect 3056 27600 3108 27606
rect 3056 27542 3108 27548
rect 3160 22094 3188 31758
rect 3252 30598 3280 33102
rect 3436 33028 3464 36060
rect 3516 36042 3568 36048
rect 3516 35828 3568 35834
rect 3516 35770 3568 35776
rect 3528 35290 3556 35770
rect 3608 35488 3660 35494
rect 3608 35430 3660 35436
rect 3516 35284 3568 35290
rect 3516 35226 3568 35232
rect 3516 34060 3568 34066
rect 3516 34002 3568 34008
rect 3528 33522 3556 34002
rect 3516 33516 3568 33522
rect 3516 33458 3568 33464
rect 3344 33000 3464 33028
rect 3240 30592 3292 30598
rect 3240 30534 3292 30540
rect 3240 29504 3292 29510
rect 3240 29446 3292 29452
rect 3252 29170 3280 29446
rect 3240 29164 3292 29170
rect 3240 29106 3292 29112
rect 3240 28076 3292 28082
rect 3240 28018 3292 28024
rect 3252 27402 3280 28018
rect 3240 27396 3292 27402
rect 3240 27338 3292 27344
rect 3344 26586 3372 33000
rect 3528 32978 3556 33458
rect 3516 32972 3568 32978
rect 3516 32914 3568 32920
rect 3528 32434 3556 32914
rect 3516 32428 3568 32434
rect 3516 32370 3568 32376
rect 3620 32314 3648 35430
rect 3528 32286 3648 32314
rect 3424 31816 3476 31822
rect 3422 31784 3424 31793
rect 3476 31784 3478 31793
rect 3422 31719 3478 31728
rect 3424 31340 3476 31346
rect 3424 31282 3476 31288
rect 3436 30433 3464 31282
rect 3422 30424 3478 30433
rect 3422 30359 3478 30368
rect 3424 30320 3476 30326
rect 3424 30262 3476 30268
rect 3436 30190 3464 30262
rect 3424 30184 3476 30190
rect 3424 30126 3476 30132
rect 3436 27674 3464 30126
rect 3528 29050 3556 32286
rect 3608 31884 3660 31890
rect 3608 31826 3660 31832
rect 3620 30326 3648 31826
rect 3608 30320 3660 30326
rect 3608 30262 3660 30268
rect 3606 29744 3662 29753
rect 3606 29679 3608 29688
rect 3660 29679 3662 29688
rect 3608 29650 3660 29656
rect 3528 29022 3648 29050
rect 3620 28966 3648 29022
rect 3608 28960 3660 28966
rect 3608 28902 3660 28908
rect 3424 27668 3476 27674
rect 3424 27610 3476 27616
rect 3332 26580 3384 26586
rect 3332 26522 3384 26528
rect 3424 25152 3476 25158
rect 3424 25094 3476 25100
rect 3332 24812 3384 24818
rect 3332 24754 3384 24760
rect 3344 24410 3372 24754
rect 3436 24614 3464 25094
rect 3424 24608 3476 24614
rect 3424 24550 3476 24556
rect 3332 24404 3384 24410
rect 3332 24346 3384 24352
rect 3240 23860 3292 23866
rect 3240 23802 3292 23808
rect 3252 23322 3280 23802
rect 3620 23730 3648 28902
rect 3712 27130 3740 36790
rect 3896 36242 3924 37266
rect 4620 36576 4672 36582
rect 4620 36518 4672 36524
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4632 36378 4660 36518
rect 4816 36394 4844 37266
rect 4620 36372 4672 36378
rect 4620 36314 4672 36320
rect 4724 36366 4844 36394
rect 3884 36236 3936 36242
rect 3884 36178 3936 36184
rect 3792 35760 3844 35766
rect 3896 35737 3924 36178
rect 4724 36038 4752 36366
rect 4804 36236 4856 36242
rect 4804 36178 4856 36184
rect 4712 36032 4764 36038
rect 4712 35974 4764 35980
rect 3792 35702 3844 35708
rect 3882 35728 3938 35737
rect 3804 35601 3832 35702
rect 3882 35663 3938 35672
rect 3976 35692 4028 35698
rect 3790 35592 3846 35601
rect 3790 35527 3846 35536
rect 3792 34944 3844 34950
rect 3792 34886 3844 34892
rect 3804 34474 3832 34886
rect 3896 34610 3924 35663
rect 3976 35634 4028 35640
rect 3884 34604 3936 34610
rect 3884 34546 3936 34552
rect 3792 34468 3844 34474
rect 3792 34410 3844 34416
rect 3804 33946 3832 34410
rect 3896 34066 3924 34546
rect 3884 34060 3936 34066
rect 3884 34002 3936 34008
rect 3804 33918 3924 33946
rect 3792 32428 3844 32434
rect 3792 32370 3844 32376
rect 3804 31346 3832 32370
rect 3792 31340 3844 31346
rect 3792 31282 3844 31288
rect 3804 30258 3832 31282
rect 3792 30252 3844 30258
rect 3792 30194 3844 30200
rect 3804 29714 3832 30194
rect 3792 29708 3844 29714
rect 3792 29650 3844 29656
rect 3804 29510 3832 29650
rect 3792 29504 3844 29510
rect 3792 29446 3844 29452
rect 3792 28076 3844 28082
rect 3792 28018 3844 28024
rect 3804 27538 3832 28018
rect 3792 27532 3844 27538
rect 3792 27474 3844 27480
rect 3792 27396 3844 27402
rect 3792 27338 3844 27344
rect 3700 27124 3752 27130
rect 3700 27066 3752 27072
rect 3804 26994 3832 27338
rect 3792 26988 3844 26994
rect 3792 26930 3844 26936
rect 3896 25974 3924 33918
rect 3988 28694 4016 35634
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4066 35048 4122 35057
rect 4066 34983 4068 34992
rect 4120 34983 4122 34992
rect 4068 34954 4120 34960
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4252 33924 4304 33930
rect 4252 33866 4304 33872
rect 4264 33833 4292 33866
rect 4250 33824 4306 33833
rect 4250 33759 4306 33768
rect 4712 33448 4764 33454
rect 4712 33390 4764 33396
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4066 33144 4122 33153
rect 4214 33147 4522 33156
rect 4066 33079 4122 33088
rect 4080 32910 4108 33079
rect 4068 32904 4120 32910
rect 4068 32846 4120 32852
rect 4252 32836 4304 32842
rect 4252 32778 4304 32784
rect 4264 32337 4292 32778
rect 4724 32774 4752 33390
rect 4712 32768 4764 32774
rect 4712 32710 4764 32716
rect 4250 32328 4306 32337
rect 4250 32263 4306 32272
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4724 31754 4752 32710
rect 4816 32366 4844 36178
rect 4908 32910 4936 37606
rect 5080 35624 5132 35630
rect 5184 35612 5212 39200
rect 5540 37256 5592 37262
rect 5540 37198 5592 37204
rect 5356 36712 5408 36718
rect 5356 36654 5408 36660
rect 5368 35737 5396 36654
rect 5448 35760 5500 35766
rect 5354 35728 5410 35737
rect 5448 35702 5500 35708
rect 5354 35663 5356 35672
rect 5408 35663 5410 35672
rect 5356 35634 5408 35640
rect 5132 35584 5212 35612
rect 5080 35566 5132 35572
rect 5368 35018 5396 35634
rect 5356 35012 5408 35018
rect 5356 34954 5408 34960
rect 5356 34604 5408 34610
rect 5356 34546 5408 34552
rect 4988 33924 5040 33930
rect 4988 33866 5040 33872
rect 4896 32904 4948 32910
rect 4896 32846 4948 32852
rect 4804 32360 4856 32366
rect 4804 32302 4856 32308
rect 4632 31726 4752 31754
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4252 30796 4304 30802
rect 4252 30738 4304 30744
rect 4068 30728 4120 30734
rect 4066 30696 4068 30705
rect 4120 30696 4122 30705
rect 4066 30631 4122 30640
rect 4264 30394 4292 30738
rect 4252 30388 4304 30394
rect 4252 30330 4304 30336
rect 4632 30161 4660 31726
rect 4816 31686 4844 32302
rect 4908 31890 4936 32846
rect 4896 31884 4948 31890
rect 4896 31826 4948 31832
rect 4896 31748 4948 31754
rect 4896 31690 4948 31696
rect 4804 31680 4856 31686
rect 4804 31622 4856 31628
rect 4712 31408 4764 31414
rect 4712 31350 4764 31356
rect 4618 30152 4674 30161
rect 4618 30087 4674 30096
rect 4620 30048 4672 30054
rect 4620 29990 4672 29996
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4632 29510 4660 29990
rect 4620 29504 4672 29510
rect 4620 29446 4672 29452
rect 4620 29164 4672 29170
rect 4620 29106 4672 29112
rect 4528 29096 4580 29102
rect 4528 29038 4580 29044
rect 4540 28966 4568 29038
rect 4528 28960 4580 28966
rect 4528 28902 4580 28908
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4632 28762 4660 29106
rect 4620 28756 4672 28762
rect 4620 28698 4672 28704
rect 3976 28688 4028 28694
rect 3976 28630 4028 28636
rect 4160 28688 4212 28694
rect 4160 28630 4212 28636
rect 4068 28144 4120 28150
rect 4172 28098 4200 28630
rect 4724 28626 4752 31350
rect 4804 30660 4856 30666
rect 4804 30602 4856 30608
rect 4816 29306 4844 30602
rect 4908 29594 4936 31690
rect 5000 29730 5028 33866
rect 5080 31884 5132 31890
rect 5080 31826 5132 31832
rect 5092 31754 5120 31826
rect 5092 31726 5212 31754
rect 5000 29702 5120 29730
rect 4908 29566 5028 29594
rect 4896 29504 4948 29510
rect 4896 29446 4948 29452
rect 4804 29300 4856 29306
rect 4804 29242 4856 29248
rect 4804 28960 4856 28966
rect 4804 28902 4856 28908
rect 4712 28620 4764 28626
rect 4712 28562 4764 28568
rect 4620 28552 4672 28558
rect 4620 28494 4672 28500
rect 4710 28520 4766 28529
rect 4252 28416 4304 28422
rect 4252 28358 4304 28364
rect 4120 28092 4200 28098
rect 4068 28086 4200 28092
rect 4080 28070 4200 28086
rect 4264 27878 4292 28358
rect 4632 28082 4660 28494
rect 4710 28455 4766 28464
rect 4620 28076 4672 28082
rect 4620 28018 4672 28024
rect 4252 27872 4304 27878
rect 4252 27814 4304 27820
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4068 27600 4120 27606
rect 4066 27568 4068 27577
rect 4120 27568 4122 27577
rect 4066 27503 4122 27512
rect 4344 27464 4396 27470
rect 4344 27406 4396 27412
rect 4356 26790 4384 27406
rect 4632 26790 4660 28018
rect 4344 26784 4396 26790
rect 4344 26726 4396 26732
rect 4620 26784 4672 26790
rect 4620 26726 4672 26732
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 3884 25968 3936 25974
rect 3884 25910 3936 25916
rect 4632 25702 4660 26726
rect 4724 26330 4752 28455
rect 4816 26586 4844 28902
rect 4804 26580 4856 26586
rect 4804 26522 4856 26528
rect 4724 26302 4844 26330
rect 4620 25696 4672 25702
rect 4620 25638 4672 25644
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4632 25158 4660 25638
rect 4620 25152 4672 25158
rect 4620 25094 4672 25100
rect 4632 24614 4660 25094
rect 4816 24698 4844 26302
rect 4908 24818 4936 29446
rect 5000 28694 5028 29566
rect 4988 28688 5040 28694
rect 4988 28630 5040 28636
rect 5092 27946 5120 29702
rect 5080 27940 5132 27946
rect 5080 27882 5132 27888
rect 5080 26920 5132 26926
rect 5080 26862 5132 26868
rect 5092 26790 5120 26862
rect 5080 26784 5132 26790
rect 5080 26726 5132 26732
rect 4988 26240 5040 26246
rect 4988 26182 5040 26188
rect 5000 25498 5028 26182
rect 5092 25498 5120 26726
rect 4988 25492 5040 25498
rect 4988 25434 5040 25440
rect 5080 25492 5132 25498
rect 5080 25434 5132 25440
rect 5000 24954 5028 25434
rect 4988 24948 5040 24954
rect 4988 24890 5040 24896
rect 4896 24812 4948 24818
rect 4896 24754 4948 24760
rect 4816 24670 5120 24698
rect 4620 24608 4672 24614
rect 4620 24550 4672 24556
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 3884 24404 3936 24410
rect 3884 24346 3936 24352
rect 3896 23866 3924 24346
rect 4632 24070 4660 24550
rect 4620 24064 4672 24070
rect 4620 24006 4672 24012
rect 3884 23860 3936 23866
rect 3884 23802 3936 23808
rect 3608 23724 3660 23730
rect 3608 23666 3660 23672
rect 3240 23316 3292 23322
rect 3240 23258 3292 23264
rect 3792 23044 3844 23050
rect 3792 22986 3844 22992
rect 3424 22976 3476 22982
rect 3424 22918 3476 22924
rect 3068 22066 3188 22094
rect 2964 22024 3016 22030
rect 2964 21966 3016 21972
rect 2504 21684 2556 21690
rect 2504 21626 2556 21632
rect 3068 21146 3096 22066
rect 3436 21690 3464 22918
rect 3804 22778 3832 22986
rect 3792 22772 3844 22778
rect 3792 22714 3844 22720
rect 3896 22094 3924 23802
rect 4632 23526 4660 24006
rect 5092 23662 5120 24670
rect 5080 23656 5132 23662
rect 5080 23598 5132 23604
rect 4620 23520 4672 23526
rect 4620 23462 4672 23468
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4632 22982 4660 23462
rect 4620 22976 4672 22982
rect 4620 22918 4672 22924
rect 4068 22772 4120 22778
rect 4068 22714 4120 22720
rect 3620 22066 3924 22094
rect 3620 21690 3648 22066
rect 4080 21894 4108 22714
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4804 21956 4856 21962
rect 4804 21898 4856 21904
rect 4068 21888 4120 21894
rect 4068 21830 4120 21836
rect 4080 21690 4108 21830
rect 3424 21684 3476 21690
rect 3424 21626 3476 21632
rect 3608 21684 3660 21690
rect 3608 21626 3660 21632
rect 4068 21684 4120 21690
rect 4068 21626 4120 21632
rect 4080 21146 4108 21626
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 2228 21140 2280 21146
rect 2228 21082 2280 21088
rect 3056 21140 3108 21146
rect 3056 21082 3108 21088
rect 4068 21140 4120 21146
rect 4068 21082 4120 21088
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 3976 18624 4028 18630
rect 3976 18566 4028 18572
rect 3332 18080 3384 18086
rect 3332 18022 3384 18028
rect 3344 12850 3372 18022
rect 3988 16114 4016 18566
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 3976 16108 4028 16114
rect 3976 16050 4028 16056
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 3332 12844 3384 12850
rect 3332 12786 3384 12792
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4816 7478 4844 21898
rect 5092 20602 5120 23598
rect 5184 21622 5212 31726
rect 5264 31272 5316 31278
rect 5264 31214 5316 31220
rect 5276 30190 5304 31214
rect 5264 30184 5316 30190
rect 5264 30126 5316 30132
rect 5276 29073 5304 30126
rect 5368 29238 5396 34546
rect 5460 31754 5488 35702
rect 5448 31748 5500 31754
rect 5448 31690 5500 31696
rect 5552 31278 5580 37198
rect 5724 37188 5776 37194
rect 5724 37130 5776 37136
rect 5736 36854 5764 37130
rect 5816 37120 5868 37126
rect 5816 37062 5868 37068
rect 6736 37120 6788 37126
rect 6736 37062 6788 37068
rect 6828 37120 6880 37126
rect 6828 37062 6880 37068
rect 5724 36848 5776 36854
rect 5724 36790 5776 36796
rect 5632 35488 5684 35494
rect 5632 35430 5684 35436
rect 5644 34950 5672 35430
rect 5828 35018 5856 37062
rect 6748 36961 6776 37062
rect 6734 36952 6790 36961
rect 6734 36887 6790 36896
rect 6840 36718 6868 37062
rect 6828 36712 6880 36718
rect 6828 36654 6880 36660
rect 6644 35692 6696 35698
rect 6644 35634 6696 35640
rect 5908 35488 5960 35494
rect 5908 35430 5960 35436
rect 5816 35012 5868 35018
rect 5816 34954 5868 34960
rect 5632 34944 5684 34950
rect 5632 34886 5684 34892
rect 5632 34400 5684 34406
rect 5632 34342 5684 34348
rect 5540 31272 5592 31278
rect 5540 31214 5592 31220
rect 5448 30796 5500 30802
rect 5448 30738 5500 30744
rect 5356 29232 5408 29238
rect 5356 29174 5408 29180
rect 5262 29064 5318 29073
rect 5262 28999 5318 29008
rect 5354 28792 5410 28801
rect 5354 28727 5410 28736
rect 5368 28694 5396 28727
rect 5356 28688 5408 28694
rect 5356 28630 5408 28636
rect 5264 28552 5316 28558
rect 5264 28494 5316 28500
rect 5276 28218 5304 28494
rect 5264 28212 5316 28218
rect 5264 28154 5316 28160
rect 5264 28076 5316 28082
rect 5264 28018 5316 28024
rect 5276 27538 5304 28018
rect 5264 27532 5316 27538
rect 5264 27474 5316 27480
rect 5356 26784 5408 26790
rect 5356 26726 5408 26732
rect 5368 26246 5396 26726
rect 5356 26240 5408 26246
rect 5356 26182 5408 26188
rect 5460 22778 5488 30738
rect 5540 30660 5592 30666
rect 5540 30602 5592 30608
rect 5552 30054 5580 30602
rect 5540 30048 5592 30054
rect 5540 29990 5592 29996
rect 5552 29714 5580 29990
rect 5540 29708 5592 29714
rect 5540 29650 5592 29656
rect 5552 27334 5580 29650
rect 5644 29510 5672 34342
rect 5724 33992 5776 33998
rect 5724 33934 5776 33940
rect 5736 33454 5764 33934
rect 5816 33924 5868 33930
rect 5816 33866 5868 33872
rect 5724 33448 5776 33454
rect 5724 33390 5776 33396
rect 5736 32910 5764 33390
rect 5724 32904 5776 32910
rect 5724 32846 5776 32852
rect 5736 31822 5764 32846
rect 5724 31816 5776 31822
rect 5724 31758 5776 31764
rect 5736 30734 5764 31758
rect 5828 31414 5856 33866
rect 5920 32502 5948 35430
rect 6276 35080 6328 35086
rect 6276 35022 6328 35028
rect 6288 34610 6316 35022
rect 6552 35012 6604 35018
rect 6552 34954 6604 34960
rect 6276 34604 6328 34610
rect 6276 34546 6328 34552
rect 6460 34468 6512 34474
rect 6460 34410 6512 34416
rect 6184 34400 6236 34406
rect 6184 34342 6236 34348
rect 6000 33584 6052 33590
rect 6000 33526 6052 33532
rect 6012 32502 6040 33526
rect 6092 32836 6144 32842
rect 6092 32778 6144 32784
rect 5908 32496 5960 32502
rect 5908 32438 5960 32444
rect 6000 32496 6052 32502
rect 6000 32438 6052 32444
rect 5908 31748 5960 31754
rect 5908 31690 5960 31696
rect 5816 31408 5868 31414
rect 5816 31350 5868 31356
rect 5816 31272 5868 31278
rect 5816 31214 5868 31220
rect 5724 30728 5776 30734
rect 5724 30670 5776 30676
rect 5722 30424 5778 30433
rect 5722 30359 5778 30368
rect 5736 29714 5764 30359
rect 5724 29708 5776 29714
rect 5724 29650 5776 29656
rect 5828 29594 5856 31214
rect 5920 30394 5948 31690
rect 6012 30410 6040 32438
rect 6104 31142 6132 32778
rect 6092 31136 6144 31142
rect 6092 31078 6144 31084
rect 5908 30388 5960 30394
rect 6012 30382 6132 30410
rect 5908 30330 5960 30336
rect 6000 30252 6052 30258
rect 6000 30194 6052 30200
rect 5906 30152 5962 30161
rect 5906 30087 5962 30096
rect 5736 29566 5856 29594
rect 5632 29504 5684 29510
rect 5632 29446 5684 29452
rect 5630 29336 5686 29345
rect 5630 29271 5632 29280
rect 5684 29271 5686 29280
rect 5632 29242 5684 29248
rect 5644 27418 5672 29242
rect 5736 27606 5764 29566
rect 5816 29504 5868 29510
rect 5816 29446 5868 29452
rect 5724 27600 5776 27606
rect 5724 27542 5776 27548
rect 5644 27390 5764 27418
rect 5540 27328 5592 27334
rect 5540 27270 5592 27276
rect 5552 26790 5580 27270
rect 5540 26784 5592 26790
rect 5540 26726 5592 26732
rect 5552 26314 5580 26726
rect 5540 26308 5592 26314
rect 5540 26250 5592 26256
rect 5552 25702 5580 26250
rect 5540 25696 5592 25702
rect 5540 25638 5592 25644
rect 5552 22982 5580 25638
rect 5632 25288 5684 25294
rect 5632 25230 5684 25236
rect 5644 24682 5672 25230
rect 5632 24676 5684 24682
rect 5632 24618 5684 24624
rect 5736 24274 5764 27390
rect 5828 25906 5856 29446
rect 5920 28914 5948 30087
rect 6012 30054 6040 30194
rect 6000 30048 6052 30054
rect 6000 29990 6052 29996
rect 6000 29504 6052 29510
rect 6000 29446 6052 29452
rect 6012 29306 6040 29446
rect 6000 29300 6052 29306
rect 6000 29242 6052 29248
rect 5920 28886 6040 28914
rect 6012 26790 6040 28886
rect 6104 27606 6132 30382
rect 6196 29345 6224 34342
rect 6472 33930 6500 34410
rect 6460 33924 6512 33930
rect 6460 33866 6512 33872
rect 6368 31748 6420 31754
rect 6368 31690 6420 31696
rect 6380 31657 6408 31690
rect 6366 31648 6422 31657
rect 6366 31583 6422 31592
rect 6276 31136 6328 31142
rect 6276 31078 6328 31084
rect 6288 30054 6316 31078
rect 6380 30870 6408 31583
rect 6368 30864 6420 30870
rect 6368 30806 6420 30812
rect 6368 30388 6420 30394
rect 6368 30330 6420 30336
rect 6276 30048 6328 30054
rect 6276 29990 6328 29996
rect 6276 29640 6328 29646
rect 6276 29582 6328 29588
rect 6288 29481 6316 29582
rect 6274 29472 6330 29481
rect 6274 29407 6330 29416
rect 6182 29336 6238 29345
rect 6182 29271 6238 29280
rect 6182 29200 6238 29209
rect 6182 29135 6238 29144
rect 6092 27600 6144 27606
rect 6092 27542 6144 27548
rect 6000 26784 6052 26790
rect 6000 26726 6052 26732
rect 5816 25900 5868 25906
rect 5816 25842 5868 25848
rect 5816 25764 5868 25770
rect 5816 25706 5868 25712
rect 5724 24268 5776 24274
rect 5724 24210 5776 24216
rect 5828 23594 5856 25706
rect 5908 24336 5960 24342
rect 5908 24278 5960 24284
rect 5920 23866 5948 24278
rect 5908 23860 5960 23866
rect 5908 23802 5960 23808
rect 5816 23588 5868 23594
rect 5816 23530 5868 23536
rect 5540 22976 5592 22982
rect 5540 22918 5592 22924
rect 5448 22772 5500 22778
rect 5448 22714 5500 22720
rect 5264 21888 5316 21894
rect 5264 21830 5316 21836
rect 5172 21616 5224 21622
rect 5172 21558 5224 21564
rect 5080 20596 5132 20602
rect 5080 20538 5132 20544
rect 5276 13938 5304 21830
rect 5460 18222 5488 22714
rect 5552 22438 5580 22918
rect 6012 22710 6040 26726
rect 6196 25838 6224 29135
rect 6274 29064 6330 29073
rect 6274 28999 6276 29008
rect 6328 28999 6330 29008
rect 6276 28970 6328 28976
rect 6274 28928 6330 28937
rect 6274 28863 6330 28872
rect 6288 27946 6316 28863
rect 6276 27940 6328 27946
rect 6276 27882 6328 27888
rect 6184 25832 6236 25838
rect 6184 25774 6236 25780
rect 6196 25158 6224 25774
rect 6184 25152 6236 25158
rect 6184 25094 6236 25100
rect 6380 23050 6408 30330
rect 6472 24818 6500 33866
rect 6564 32502 6592 34954
rect 6656 34202 6684 35634
rect 7116 34542 7144 39200
rect 8404 37346 8432 39200
rect 10232 37460 10284 37466
rect 10232 37402 10284 37408
rect 8404 37318 8524 37346
rect 7840 37188 7892 37194
rect 7840 37130 7892 37136
rect 7852 36922 7880 37130
rect 7840 36916 7892 36922
rect 7840 36858 7892 36864
rect 8392 36576 8444 36582
rect 8392 36518 8444 36524
rect 8116 36236 8168 36242
rect 8116 36178 8168 36184
rect 8128 35850 8156 36178
rect 8404 36174 8432 36518
rect 8392 36168 8444 36174
rect 8392 36110 8444 36116
rect 8036 35834 8156 35850
rect 8496 35834 8524 37318
rect 9864 37324 9916 37330
rect 9864 37266 9916 37272
rect 8944 37256 8996 37262
rect 8944 37198 8996 37204
rect 8668 36848 8720 36854
rect 8668 36790 8720 36796
rect 8576 36780 8628 36786
rect 8576 36722 8628 36728
rect 8588 36242 8616 36722
rect 8576 36236 8628 36242
rect 8576 36178 8628 36184
rect 8024 35828 8156 35834
rect 8076 35822 8156 35828
rect 8024 35770 8076 35776
rect 7472 35556 7524 35562
rect 7472 35498 7524 35504
rect 7196 35488 7248 35494
rect 7484 35465 7512 35498
rect 7196 35430 7248 35436
rect 7470 35456 7526 35465
rect 7104 34536 7156 34542
rect 7104 34478 7156 34484
rect 6826 34368 6882 34377
rect 6826 34303 6882 34312
rect 6644 34196 6696 34202
rect 6644 34138 6696 34144
rect 6552 32496 6604 32502
rect 6552 32438 6604 32444
rect 6552 32360 6604 32366
rect 6552 32302 6604 32308
rect 6564 29209 6592 32302
rect 6656 30705 6684 34138
rect 6840 33590 6868 34303
rect 7208 33674 7236 35430
rect 7470 35391 7526 35400
rect 7656 35216 7708 35222
rect 7656 35158 7708 35164
rect 7288 34672 7340 34678
rect 7340 34632 7420 34660
rect 7288 34614 7340 34620
rect 7392 34406 7420 34632
rect 7380 34400 7432 34406
rect 7380 34342 7432 34348
rect 7208 33646 7328 33674
rect 6828 33584 6880 33590
rect 6828 33526 6880 33532
rect 7196 32904 7248 32910
rect 7196 32846 7248 32852
rect 7012 32496 7064 32502
rect 7012 32438 7064 32444
rect 6736 31952 6788 31958
rect 6736 31894 6788 31900
rect 6748 31278 6776 31894
rect 7024 31754 7052 32438
rect 6920 31748 6972 31754
rect 7024 31726 7144 31754
rect 6920 31690 6972 31696
rect 6736 31272 6788 31278
rect 6736 31214 6788 31220
rect 6642 30696 6698 30705
rect 6642 30631 6698 30640
rect 6748 30580 6776 31214
rect 6932 30938 6960 31690
rect 7116 31482 7144 31726
rect 7104 31476 7156 31482
rect 7104 31418 7156 31424
rect 7012 31408 7064 31414
rect 7012 31350 7064 31356
rect 6920 30932 6972 30938
rect 6920 30874 6972 30880
rect 6920 30660 6972 30666
rect 6920 30602 6972 30608
rect 6656 30552 6776 30580
rect 6656 30161 6684 30552
rect 6828 30320 6880 30326
rect 6828 30262 6880 30268
rect 6736 30252 6788 30258
rect 6736 30194 6788 30200
rect 6642 30152 6698 30161
rect 6642 30087 6698 30096
rect 6642 29880 6698 29889
rect 6642 29815 6644 29824
rect 6696 29815 6698 29824
rect 6644 29786 6696 29792
rect 6748 29714 6776 30194
rect 6840 29850 6868 30262
rect 6828 29844 6880 29850
rect 6828 29786 6880 29792
rect 6736 29708 6788 29714
rect 6736 29650 6788 29656
rect 6828 29572 6880 29578
rect 6828 29514 6880 29520
rect 6642 29472 6698 29481
rect 6642 29407 6698 29416
rect 6656 29238 6684 29407
rect 6644 29232 6696 29238
rect 6550 29200 6606 29209
rect 6644 29174 6696 29180
rect 6550 29135 6606 29144
rect 6736 29164 6788 29170
rect 6564 26450 6592 29135
rect 6736 29106 6788 29112
rect 6644 29096 6696 29102
rect 6748 29073 6776 29106
rect 6644 29038 6696 29044
rect 6734 29064 6790 29073
rect 6656 28626 6684 29038
rect 6734 28999 6790 29008
rect 6644 28620 6696 28626
rect 6644 28562 6696 28568
rect 6642 28520 6698 28529
rect 6840 28506 6868 29514
rect 6932 29510 6960 30602
rect 6920 29504 6972 29510
rect 6920 29446 6972 29452
rect 7024 28694 7052 31350
rect 7104 30184 7156 30190
rect 7104 30126 7156 30132
rect 7012 28688 7064 28694
rect 7012 28630 7064 28636
rect 7116 28506 7144 30126
rect 6748 28490 6868 28506
rect 6642 28455 6698 28464
rect 6736 28484 6868 28490
rect 6656 27334 6684 28455
rect 6788 28478 6868 28484
rect 7024 28478 7144 28506
rect 6736 28426 6788 28432
rect 6828 28416 6880 28422
rect 6880 28376 6960 28404
rect 6828 28358 6880 28364
rect 6828 28076 6880 28082
rect 6828 28018 6880 28024
rect 6840 27402 6868 28018
rect 6828 27396 6880 27402
rect 6828 27338 6880 27344
rect 6932 27334 6960 28376
rect 6644 27328 6696 27334
rect 6644 27270 6696 27276
rect 6920 27328 6972 27334
rect 6920 27270 6972 27276
rect 6552 26444 6604 26450
rect 6552 26386 6604 26392
rect 6460 24812 6512 24818
rect 6460 24754 6512 24760
rect 6656 24070 6684 27270
rect 6828 26852 6880 26858
rect 6828 26794 6880 26800
rect 6736 25152 6788 25158
rect 6736 25094 6788 25100
rect 6748 24818 6776 25094
rect 6736 24812 6788 24818
rect 6736 24754 6788 24760
rect 6840 24410 6868 26794
rect 6828 24404 6880 24410
rect 6828 24346 6880 24352
rect 6644 24064 6696 24070
rect 6644 24006 6696 24012
rect 6656 23798 6684 24006
rect 6644 23792 6696 23798
rect 6644 23734 6696 23740
rect 6368 23044 6420 23050
rect 6368 22986 6420 22992
rect 6000 22704 6052 22710
rect 6000 22646 6052 22652
rect 5540 22432 5592 22438
rect 5540 22374 5592 22380
rect 6460 22432 6512 22438
rect 6460 22374 6512 22380
rect 6472 22166 6500 22374
rect 6460 22160 6512 22166
rect 6460 22102 6512 22108
rect 6472 21690 6500 22102
rect 7024 22094 7052 28478
rect 7208 28014 7236 32846
rect 7300 32570 7328 33646
rect 7564 33108 7616 33114
rect 7564 33050 7616 33056
rect 7380 32904 7432 32910
rect 7380 32846 7432 32852
rect 7288 32564 7340 32570
rect 7288 32506 7340 32512
rect 7288 32224 7340 32230
rect 7288 32166 7340 32172
rect 7300 30190 7328 32166
rect 7288 30184 7340 30190
rect 7288 30126 7340 30132
rect 7392 29458 7420 32846
rect 7576 32026 7604 33050
rect 7564 32020 7616 32026
rect 7564 31962 7616 31968
rect 7668 30920 7696 35158
rect 8128 35086 8156 35822
rect 8484 35828 8536 35834
rect 8484 35770 8536 35776
rect 8680 35766 8708 36790
rect 8956 36582 8984 37198
rect 9128 37120 9180 37126
rect 9128 37062 9180 37068
rect 9140 36854 9168 37062
rect 9128 36848 9180 36854
rect 9128 36790 9180 36796
rect 9588 36848 9640 36854
rect 9588 36790 9640 36796
rect 9034 36680 9090 36689
rect 9034 36615 9036 36624
rect 9088 36615 9090 36624
rect 9036 36586 9088 36592
rect 8944 36576 8996 36582
rect 8944 36518 8996 36524
rect 8852 36168 8904 36174
rect 8852 36110 8904 36116
rect 8760 36100 8812 36106
rect 8760 36042 8812 36048
rect 8208 35760 8260 35766
rect 8208 35702 8260 35708
rect 8668 35760 8720 35766
rect 8668 35702 8720 35708
rect 8220 35494 8248 35702
rect 8208 35488 8260 35494
rect 8208 35430 8260 35436
rect 8116 35080 8168 35086
rect 8116 35022 8168 35028
rect 8024 35012 8076 35018
rect 8024 34954 8076 34960
rect 8300 35012 8352 35018
rect 8300 34954 8352 34960
rect 7746 34912 7802 34921
rect 7746 34847 7802 34856
rect 7300 29430 7420 29458
rect 7576 30892 7696 30920
rect 7300 28694 7328 29430
rect 7378 29336 7434 29345
rect 7378 29271 7434 29280
rect 7392 29170 7420 29271
rect 7380 29164 7432 29170
rect 7432 29124 7512 29152
rect 7380 29106 7432 29112
rect 7288 28688 7340 28694
rect 7288 28630 7340 28636
rect 7288 28552 7340 28558
rect 7288 28494 7340 28500
rect 7300 28082 7328 28494
rect 7484 28218 7512 29124
rect 7472 28212 7524 28218
rect 7472 28154 7524 28160
rect 7484 28082 7512 28154
rect 7288 28076 7340 28082
rect 7288 28018 7340 28024
rect 7472 28076 7524 28082
rect 7472 28018 7524 28024
rect 7196 28008 7248 28014
rect 7196 27950 7248 27956
rect 7380 27328 7432 27334
rect 7432 27288 7512 27316
rect 7380 27270 7432 27276
rect 7104 27124 7156 27130
rect 7104 27066 7156 27072
rect 7116 25906 7144 27066
rect 7484 26858 7512 27288
rect 7576 27130 7604 30892
rect 7760 30784 7788 34847
rect 7838 33688 7894 33697
rect 7838 33623 7894 33632
rect 7852 33454 7880 33623
rect 7840 33448 7892 33454
rect 7840 33390 7892 33396
rect 7668 30756 7788 30784
rect 7668 28218 7696 30756
rect 7748 30184 7800 30190
rect 7748 30126 7800 30132
rect 7656 28212 7708 28218
rect 7656 28154 7708 28160
rect 7564 27124 7616 27130
rect 7564 27066 7616 27072
rect 7472 26852 7524 26858
rect 7472 26794 7524 26800
rect 7484 26761 7512 26794
rect 7470 26752 7526 26761
rect 7470 26687 7526 26696
rect 7288 26376 7340 26382
rect 7288 26318 7340 26324
rect 7104 25900 7156 25906
rect 7104 25842 7156 25848
rect 6932 22066 7052 22094
rect 6460 21684 6512 21690
rect 6460 21626 6512 21632
rect 6932 21010 6960 22066
rect 6920 21004 6972 21010
rect 6920 20946 6972 20952
rect 7116 18970 7144 25842
rect 7196 25696 7248 25702
rect 7196 25638 7248 25644
rect 7208 25430 7236 25638
rect 7196 25424 7248 25430
rect 7196 25366 7248 25372
rect 7300 24857 7328 26318
rect 7760 26194 7788 30126
rect 7668 26166 7788 26194
rect 7668 25906 7696 26166
rect 7748 26036 7800 26042
rect 7852 26024 7880 33390
rect 8036 32881 8064 34954
rect 8116 34604 8168 34610
rect 8116 34546 8168 34552
rect 8128 33153 8156 34546
rect 8206 34232 8262 34241
rect 8312 34202 8340 34954
rect 8576 34536 8628 34542
rect 8576 34478 8628 34484
rect 8392 34400 8444 34406
rect 8392 34342 8444 34348
rect 8206 34167 8208 34176
rect 8260 34167 8262 34176
rect 8300 34196 8352 34202
rect 8208 34138 8260 34144
rect 8300 34138 8352 34144
rect 8404 33590 8432 34342
rect 8484 33924 8536 33930
rect 8484 33866 8536 33872
rect 8392 33584 8444 33590
rect 8206 33552 8262 33561
rect 8392 33526 8444 33532
rect 8206 33487 8262 33496
rect 8114 33144 8170 33153
rect 8114 33079 8170 33088
rect 8022 32872 8078 32881
rect 8022 32807 8078 32816
rect 8116 32836 8168 32842
rect 8116 32778 8168 32784
rect 8128 31754 8156 32778
rect 8116 31748 8168 31754
rect 8116 31690 8168 31696
rect 7932 31680 7984 31686
rect 7932 31622 7984 31628
rect 7944 30938 7972 31622
rect 7932 30932 7984 30938
rect 7932 30874 7984 30880
rect 8220 30376 8248 33487
rect 8300 33312 8352 33318
rect 8300 33254 8352 33260
rect 7944 30348 8248 30376
rect 7944 29510 7972 30348
rect 8312 30190 8340 33254
rect 8496 31754 8524 33866
rect 8588 33862 8616 34478
rect 8576 33856 8628 33862
rect 8576 33798 8628 33804
rect 8576 33584 8628 33590
rect 8576 33526 8628 33532
rect 8404 31726 8524 31754
rect 8300 30184 8352 30190
rect 8300 30126 8352 30132
rect 8300 29708 8352 29714
rect 8300 29650 8352 29656
rect 8312 29617 8340 29650
rect 8298 29608 8354 29617
rect 8298 29543 8354 29552
rect 7932 29504 7984 29510
rect 7932 29446 7984 29452
rect 8024 29504 8076 29510
rect 8024 29446 8076 29452
rect 7944 29073 7972 29446
rect 8036 29345 8064 29446
rect 8022 29336 8078 29345
rect 8022 29271 8078 29280
rect 8298 29336 8354 29345
rect 8298 29271 8354 29280
rect 8208 29164 8260 29170
rect 8208 29106 8260 29112
rect 7930 29064 7986 29073
rect 7930 28999 7986 29008
rect 7944 28558 7972 28999
rect 8220 28994 8248 29106
rect 8036 28966 8248 28994
rect 8036 28558 8064 28966
rect 7932 28552 7984 28558
rect 7932 28494 7984 28500
rect 8024 28552 8076 28558
rect 8024 28494 8076 28500
rect 8036 26926 8064 28494
rect 8312 28150 8340 29271
rect 8404 28529 8432 31726
rect 8484 29504 8536 29510
rect 8484 29446 8536 29452
rect 8390 28520 8446 28529
rect 8390 28455 8446 28464
rect 8300 28144 8352 28150
rect 8300 28086 8352 28092
rect 8116 27464 8168 27470
rect 8116 27406 8168 27412
rect 8024 26920 8076 26926
rect 8024 26862 8076 26868
rect 7800 25996 7880 26024
rect 7748 25978 7800 25984
rect 7656 25900 7708 25906
rect 7656 25842 7708 25848
rect 7286 24848 7342 24857
rect 7852 24818 7880 25996
rect 7932 25968 7984 25974
rect 7932 25910 7984 25916
rect 7944 24818 7972 25910
rect 7286 24783 7342 24792
rect 7840 24812 7892 24818
rect 7840 24754 7892 24760
rect 7932 24812 7984 24818
rect 7932 24754 7984 24760
rect 7564 22976 7616 22982
rect 7564 22918 7616 22924
rect 7104 18964 7156 18970
rect 7104 18906 7156 18912
rect 7472 18692 7524 18698
rect 7472 18634 7524 18640
rect 7484 18426 7512 18634
rect 7472 18420 7524 18426
rect 7472 18362 7524 18368
rect 5448 18216 5500 18222
rect 5448 18158 5500 18164
rect 5264 13932 5316 13938
rect 5264 13874 5316 13880
rect 4804 7472 4856 7478
rect 4804 7414 4856 7420
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 1582 6896 1638 6905
rect 1582 6831 1638 6840
rect 1780 6886 1992 6914
rect 1780 5370 1808 6886
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 1768 5364 1820 5370
rect 1768 5306 1820 5312
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1596 4865 1624 5170
rect 1582 4856 1638 4865
rect 1582 4791 1584 4800
rect 1636 4791 1638 4800
rect 1584 4762 1636 4768
rect 2792 3534 2820 6598
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 2780 3528 2832 3534
rect 1674 3496 1730 3505
rect 2780 3470 2832 3476
rect 1674 3431 1730 3440
rect 1952 3460 2004 3466
rect 1688 3398 1716 3431
rect 1952 3402 2004 3408
rect 1676 3392 1728 3398
rect 1676 3334 1728 3340
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1308 2304 1360 2310
rect 1308 2246 1360 2252
rect 20 1352 72 1358
rect 20 1294 72 1300
rect 32 800 60 1294
rect 1320 800 1348 2246
rect 1688 1465 1716 2994
rect 1964 2446 1992 3402
rect 7576 3194 7604 22918
rect 7852 19854 7880 24754
rect 7932 24608 7984 24614
rect 7932 24550 7984 24556
rect 7944 24274 7972 24550
rect 7932 24268 7984 24274
rect 7932 24210 7984 24216
rect 8128 21146 8156 27406
rect 8496 27062 8524 29446
rect 8588 27062 8616 33526
rect 8680 33114 8708 35702
rect 8668 33108 8720 33114
rect 8668 33050 8720 33056
rect 8668 32904 8720 32910
rect 8668 32846 8720 32852
rect 8680 32230 8708 32846
rect 8668 32224 8720 32230
rect 8668 32166 8720 32172
rect 8668 31816 8720 31822
rect 8668 31758 8720 31764
rect 8680 31346 8708 31758
rect 8668 31340 8720 31346
rect 8668 31282 8720 31288
rect 8680 30734 8708 31282
rect 8668 30728 8720 30734
rect 8668 30670 8720 30676
rect 8680 30326 8708 30670
rect 8668 30320 8720 30326
rect 8668 30262 8720 30268
rect 8666 29880 8722 29889
rect 8666 29815 8722 29824
rect 8680 29238 8708 29815
rect 8772 29510 8800 36042
rect 8760 29504 8812 29510
rect 8760 29446 8812 29452
rect 8760 29300 8812 29306
rect 8760 29242 8812 29248
rect 8668 29232 8720 29238
rect 8668 29174 8720 29180
rect 8668 28620 8720 28626
rect 8668 28562 8720 28568
rect 8680 27946 8708 28562
rect 8668 27940 8720 27946
rect 8668 27882 8720 27888
rect 8772 27402 8800 29242
rect 8760 27396 8812 27402
rect 8760 27338 8812 27344
rect 8484 27056 8536 27062
rect 8484 26998 8536 27004
rect 8576 27056 8628 27062
rect 8576 26998 8628 27004
rect 8392 26376 8444 26382
rect 8392 26318 8444 26324
rect 8404 26246 8432 26318
rect 8392 26240 8444 26246
rect 8392 26182 8444 26188
rect 8576 25832 8628 25838
rect 8576 25774 8628 25780
rect 8208 25764 8260 25770
rect 8208 25706 8260 25712
rect 8220 21894 8248 25706
rect 8392 25356 8444 25362
rect 8392 25298 8444 25304
rect 8404 24206 8432 25298
rect 8484 25220 8536 25226
rect 8484 25162 8536 25168
rect 8392 24200 8444 24206
rect 8392 24142 8444 24148
rect 8300 23792 8352 23798
rect 8300 23734 8352 23740
rect 8312 23322 8340 23734
rect 8392 23656 8444 23662
rect 8390 23624 8392 23633
rect 8444 23624 8446 23633
rect 8390 23559 8446 23568
rect 8496 23322 8524 25162
rect 8300 23316 8352 23322
rect 8300 23258 8352 23264
rect 8484 23316 8536 23322
rect 8484 23258 8536 23264
rect 8588 22642 8616 25774
rect 8864 24818 8892 36110
rect 8956 35698 8984 36518
rect 8944 35692 8996 35698
rect 8944 35634 8996 35640
rect 8956 34542 8984 35634
rect 9312 35624 9364 35630
rect 9312 35566 9364 35572
rect 9404 35624 9456 35630
rect 9404 35566 9456 35572
rect 9128 35080 9180 35086
rect 9128 35022 9180 35028
rect 9140 34678 9168 35022
rect 9128 34672 9180 34678
rect 9128 34614 9180 34620
rect 8944 34536 8996 34542
rect 8944 34478 8996 34484
rect 8956 34066 8984 34478
rect 9324 34105 9352 35566
rect 9310 34096 9366 34105
rect 8944 34060 8996 34066
rect 8944 34002 8996 34008
rect 9232 34054 9310 34082
rect 8956 33522 8984 34002
rect 9128 33924 9180 33930
rect 9128 33866 9180 33872
rect 9036 33856 9088 33862
rect 9036 33798 9088 33804
rect 8944 33516 8996 33522
rect 8944 33458 8996 33464
rect 9048 31754 9076 33798
rect 9140 32366 9168 33866
rect 9128 32360 9180 32366
rect 9128 32302 9180 32308
rect 8956 31726 9076 31754
rect 8956 26314 8984 31726
rect 9128 31476 9180 31482
rect 9128 31418 9180 31424
rect 9140 29578 9168 31418
rect 9128 29572 9180 29578
rect 9128 29514 9180 29520
rect 9034 29064 9090 29073
rect 9034 28999 9090 29008
rect 9048 28558 9076 28999
rect 9232 28608 9260 34054
rect 9310 34031 9366 34040
rect 9312 32972 9364 32978
rect 9312 32914 9364 32920
rect 9324 32434 9352 32914
rect 9312 32428 9364 32434
rect 9312 32370 9364 32376
rect 9310 32328 9366 32337
rect 9310 32263 9312 32272
rect 9364 32263 9366 32272
rect 9312 32234 9364 32240
rect 9312 30864 9364 30870
rect 9312 30806 9364 30812
rect 9324 30122 9352 30806
rect 9312 30116 9364 30122
rect 9312 30058 9364 30064
rect 9310 29744 9366 29753
rect 9310 29679 9366 29688
rect 9324 29646 9352 29679
rect 9312 29640 9364 29646
rect 9312 29582 9364 29588
rect 9416 28937 9444 35566
rect 9600 34542 9628 36790
rect 9876 36718 9904 37266
rect 9864 36712 9916 36718
rect 9864 36654 9916 36660
rect 9680 36100 9732 36106
rect 9680 36042 9732 36048
rect 9588 34536 9640 34542
rect 9588 34478 9640 34484
rect 9496 33108 9548 33114
rect 9496 33050 9548 33056
rect 9508 32842 9536 33050
rect 9588 32904 9640 32910
rect 9588 32846 9640 32852
rect 9496 32836 9548 32842
rect 9496 32778 9548 32784
rect 9600 32570 9628 32846
rect 9496 32564 9548 32570
rect 9496 32506 9548 32512
rect 9588 32564 9640 32570
rect 9588 32506 9640 32512
rect 9508 31958 9536 32506
rect 9600 32473 9628 32506
rect 9692 32502 9720 36042
rect 9772 35692 9824 35698
rect 9772 35634 9824 35640
rect 9784 34649 9812 35634
rect 9864 35556 9916 35562
rect 9864 35498 9916 35504
rect 9770 34640 9826 34649
rect 9770 34575 9826 34584
rect 9876 34542 9904 35498
rect 10244 34728 10272 37402
rect 10336 36310 10364 39200
rect 10600 37732 10652 37738
rect 10600 37674 10652 37680
rect 10612 37466 10640 37674
rect 10600 37460 10652 37466
rect 10600 37402 10652 37408
rect 10968 37324 11020 37330
rect 10968 37266 11020 37272
rect 10692 37188 10744 37194
rect 10692 37130 10744 37136
rect 10600 36848 10652 36854
rect 10600 36790 10652 36796
rect 10324 36304 10376 36310
rect 10324 36246 10376 36252
rect 10336 36174 10364 36246
rect 10324 36168 10376 36174
rect 10324 36110 10376 36116
rect 10612 35834 10640 36790
rect 10704 36145 10732 37130
rect 10980 37097 11008 37266
rect 11520 37256 11572 37262
rect 11520 37198 11572 37204
rect 10966 37088 11022 37097
rect 10966 37023 11022 37032
rect 11072 37046 11376 37074
rect 10876 36712 10928 36718
rect 10876 36654 10928 36660
rect 10690 36136 10746 36145
rect 10690 36071 10746 36080
rect 10600 35828 10652 35834
rect 10600 35770 10652 35776
rect 10692 35828 10744 35834
rect 10692 35770 10744 35776
rect 10704 35714 10732 35770
rect 10520 35686 10732 35714
rect 10784 35760 10836 35766
rect 10784 35702 10836 35708
rect 10520 35630 10548 35686
rect 10508 35624 10560 35630
rect 10508 35566 10560 35572
rect 10796 35442 10824 35702
rect 10888 35494 10916 36654
rect 10704 35414 10824 35442
rect 10876 35488 10928 35494
rect 10876 35430 10928 35436
rect 10704 35290 10732 35414
rect 10692 35284 10744 35290
rect 10692 35226 10744 35232
rect 10782 35184 10838 35193
rect 10782 35119 10838 35128
rect 10796 35086 10824 35119
rect 10784 35080 10836 35086
rect 10784 35022 10836 35028
rect 10876 35012 10928 35018
rect 10876 34954 10928 34960
rect 10244 34700 10548 34728
rect 10520 34610 10548 34700
rect 10888 34649 10916 34954
rect 10874 34640 10930 34649
rect 10508 34604 10560 34610
rect 10874 34575 10930 34584
rect 10508 34546 10560 34552
rect 9772 34536 9824 34542
rect 9772 34478 9824 34484
rect 9864 34536 9916 34542
rect 9864 34478 9916 34484
rect 9680 32496 9732 32502
rect 9586 32464 9642 32473
rect 9680 32438 9732 32444
rect 9586 32399 9642 32408
rect 9588 32360 9640 32366
rect 9588 32302 9640 32308
rect 9496 31952 9548 31958
rect 9494 31920 9496 31929
rect 9548 31920 9550 31929
rect 9494 31855 9550 31864
rect 9496 31408 9548 31414
rect 9496 31350 9548 31356
rect 9508 29578 9536 31350
rect 9600 30734 9628 32302
rect 9692 31890 9720 32438
rect 9680 31884 9732 31890
rect 9680 31826 9732 31832
rect 9588 30728 9640 30734
rect 9588 30670 9640 30676
rect 9680 30592 9732 30598
rect 9680 30534 9732 30540
rect 9692 30394 9720 30534
rect 9680 30388 9732 30394
rect 9680 30330 9732 30336
rect 9588 29640 9640 29646
rect 9588 29582 9640 29588
rect 9496 29572 9548 29578
rect 9496 29514 9548 29520
rect 9600 29481 9628 29582
rect 9680 29572 9732 29578
rect 9680 29514 9732 29520
rect 9586 29472 9642 29481
rect 9586 29407 9642 29416
rect 9692 29322 9720 29514
rect 9784 29481 9812 34478
rect 10692 34400 10744 34406
rect 10692 34342 10744 34348
rect 10704 34066 10732 34342
rect 10692 34060 10744 34066
rect 10692 34002 10744 34008
rect 9864 33448 9916 33454
rect 9864 33390 9916 33396
rect 9876 33289 9904 33390
rect 9862 33280 9918 33289
rect 9862 33215 9918 33224
rect 10048 32836 10100 32842
rect 10048 32778 10100 32784
rect 9956 32768 10008 32774
rect 9954 32736 9956 32745
rect 10008 32736 10010 32745
rect 9954 32671 10010 32680
rect 9864 31816 9916 31822
rect 9864 31758 9916 31764
rect 9876 29782 9904 31758
rect 10060 30258 10088 32778
rect 10230 31512 10286 31521
rect 10140 31476 10192 31482
rect 10230 31447 10286 31456
rect 10140 31418 10192 31424
rect 10152 31385 10180 31418
rect 10138 31376 10194 31385
rect 10138 31311 10194 31320
rect 10244 30734 10272 31447
rect 10416 31408 10468 31414
rect 10416 31350 10468 31356
rect 10600 31408 10652 31414
rect 10600 31350 10652 31356
rect 10232 30728 10284 30734
rect 10232 30670 10284 30676
rect 10048 30252 10100 30258
rect 9968 30212 10048 30240
rect 9864 29776 9916 29782
rect 9864 29718 9916 29724
rect 9770 29472 9826 29481
rect 9770 29407 9826 29416
rect 9692 29294 9904 29322
rect 9772 29232 9824 29238
rect 9770 29200 9772 29209
rect 9824 29200 9826 29209
rect 9770 29135 9826 29144
rect 9402 28928 9458 28937
rect 9402 28863 9458 28872
rect 9140 28580 9352 28608
rect 9036 28552 9088 28558
rect 9036 28494 9088 28500
rect 9034 27976 9090 27985
rect 9034 27911 9090 27920
rect 9048 27878 9076 27911
rect 9036 27872 9088 27878
rect 9036 27814 9088 27820
rect 9140 27614 9168 28580
rect 9324 28490 9352 28580
rect 9220 28484 9272 28490
rect 9220 28426 9272 28432
rect 9312 28484 9364 28490
rect 9312 28426 9364 28432
rect 9232 28393 9260 28426
rect 9772 28416 9824 28422
rect 9218 28384 9274 28393
rect 9772 28358 9824 28364
rect 9218 28319 9274 28328
rect 9784 28218 9812 28358
rect 9772 28212 9824 28218
rect 9772 28154 9824 28160
rect 9048 27586 9168 27614
rect 9048 26382 9076 27586
rect 9876 27538 9904 29294
rect 9968 28422 9996 30212
rect 10048 30194 10100 30200
rect 10324 30252 10376 30258
rect 10324 30194 10376 30200
rect 10336 30054 10364 30194
rect 10324 30048 10376 30054
rect 10324 29990 10376 29996
rect 10138 29880 10194 29889
rect 10428 29832 10456 31350
rect 10612 30870 10640 31350
rect 10600 30864 10652 30870
rect 10600 30806 10652 30812
rect 10600 30728 10652 30734
rect 10600 30670 10652 30676
rect 10508 30660 10560 30666
rect 10508 30602 10560 30608
rect 10138 29815 10194 29824
rect 10152 29578 10180 29815
rect 10336 29804 10456 29832
rect 10140 29572 10192 29578
rect 10140 29514 10192 29520
rect 10232 29572 10284 29578
rect 10232 29514 10284 29520
rect 10244 29458 10272 29514
rect 10152 29430 10272 29458
rect 10152 29152 10180 29430
rect 10336 29152 10364 29804
rect 10414 29744 10470 29753
rect 10414 29679 10416 29688
rect 10468 29679 10470 29688
rect 10416 29650 10468 29656
rect 10416 29300 10468 29306
rect 10416 29242 10468 29248
rect 10428 29209 10456 29242
rect 10060 29124 10180 29152
rect 10244 29124 10364 29152
rect 10414 29200 10470 29209
rect 10414 29135 10470 29144
rect 9956 28416 10008 28422
rect 10060 28393 10088 29124
rect 10244 28694 10272 29124
rect 10520 29102 10548 30602
rect 10612 29152 10640 30670
rect 10704 29220 10732 34002
rect 10784 33992 10836 33998
rect 10784 33934 10836 33940
rect 10796 33862 10824 33934
rect 10784 33856 10836 33862
rect 10784 33798 10836 33804
rect 10784 33516 10836 33522
rect 10784 33458 10836 33464
rect 10796 33046 10824 33458
rect 10784 33040 10836 33046
rect 10784 32982 10836 32988
rect 10966 32736 11022 32745
rect 10966 32671 11022 32680
rect 10980 32230 11008 32671
rect 10968 32224 11020 32230
rect 10968 32166 11020 32172
rect 10874 31920 10930 31929
rect 10874 31855 10930 31864
rect 10968 31884 11020 31890
rect 10784 31272 10836 31278
rect 10784 31214 10836 31220
rect 10796 29753 10824 31214
rect 10888 30977 10916 31855
rect 10968 31826 11020 31832
rect 10980 31793 11008 31826
rect 10966 31784 11022 31793
rect 10966 31719 11022 31728
rect 10874 30968 10930 30977
rect 10874 30903 10930 30912
rect 10876 30864 10928 30870
rect 10876 30806 10928 30812
rect 10782 29744 10838 29753
rect 10782 29679 10838 29688
rect 10704 29192 10824 29220
rect 10612 29124 10732 29152
rect 10508 29096 10560 29102
rect 10414 29064 10470 29073
rect 10336 29022 10414 29050
rect 10232 28688 10284 28694
rect 10232 28630 10284 28636
rect 9956 28358 10008 28364
rect 10046 28384 10102 28393
rect 10046 28319 10102 28328
rect 10048 28144 10100 28150
rect 10048 28086 10100 28092
rect 10232 28144 10284 28150
rect 10232 28086 10284 28092
rect 9956 27872 10008 27878
rect 10060 27849 10088 28086
rect 9956 27814 10008 27820
rect 10046 27840 10102 27849
rect 9864 27532 9916 27538
rect 9864 27474 9916 27480
rect 9128 27328 9180 27334
rect 9128 27270 9180 27276
rect 9772 27328 9824 27334
rect 9772 27270 9824 27276
rect 9140 26790 9168 27270
rect 9496 27056 9548 27062
rect 9496 26998 9548 27004
rect 9128 26784 9180 26790
rect 9128 26726 9180 26732
rect 9036 26376 9088 26382
rect 9036 26318 9088 26324
rect 8944 26308 8996 26314
rect 8944 26250 8996 26256
rect 8668 24812 8720 24818
rect 8668 24754 8720 24760
rect 8852 24812 8904 24818
rect 8852 24754 8904 24760
rect 8680 24585 8708 24754
rect 8666 24576 8722 24585
rect 8666 24511 8722 24520
rect 8864 23186 8892 24754
rect 8956 24206 8984 26250
rect 8944 24200 8996 24206
rect 8944 24142 8996 24148
rect 8852 23180 8904 23186
rect 8852 23122 8904 23128
rect 8668 23044 8720 23050
rect 8668 22986 8720 22992
rect 8680 22778 8708 22986
rect 8668 22772 8720 22778
rect 8668 22714 8720 22720
rect 8576 22636 8628 22642
rect 8576 22578 8628 22584
rect 8208 21888 8260 21894
rect 8208 21830 8260 21836
rect 8588 21554 8616 22578
rect 8576 21548 8628 21554
rect 8576 21490 8628 21496
rect 8116 21140 8168 21146
rect 8116 21082 8168 21088
rect 7840 19848 7892 19854
rect 7840 19790 7892 19796
rect 9048 19334 9076 26318
rect 9220 26308 9272 26314
rect 9220 26250 9272 26256
rect 9312 26308 9364 26314
rect 9312 26250 9364 26256
rect 9128 26240 9180 26246
rect 9128 26182 9180 26188
rect 9140 25838 9168 26182
rect 9128 25832 9180 25838
rect 9128 25774 9180 25780
rect 9140 25498 9168 25774
rect 9232 25770 9260 26250
rect 9220 25764 9272 25770
rect 9220 25706 9272 25712
rect 9128 25492 9180 25498
rect 9128 25434 9180 25440
rect 9324 24750 9352 26250
rect 9404 25968 9456 25974
rect 9404 25910 9456 25916
rect 9416 25362 9444 25910
rect 9404 25356 9456 25362
rect 9404 25298 9456 25304
rect 9312 24744 9364 24750
rect 9312 24686 9364 24692
rect 9508 24614 9536 26998
rect 9784 25702 9812 27270
rect 9864 26920 9916 26926
rect 9864 26862 9916 26868
rect 9876 26314 9904 26862
rect 9968 26790 9996 27814
rect 10046 27775 10102 27784
rect 10138 27704 10194 27713
rect 10138 27639 10140 27648
rect 10192 27639 10194 27648
rect 10140 27610 10192 27616
rect 10048 27600 10100 27606
rect 10244 27554 10272 28086
rect 10100 27548 10272 27554
rect 10048 27542 10272 27548
rect 10060 27526 10272 27542
rect 10232 26988 10284 26994
rect 10232 26930 10284 26936
rect 10138 26888 10194 26897
rect 10138 26823 10194 26832
rect 9956 26784 10008 26790
rect 9956 26726 10008 26732
rect 9864 26308 9916 26314
rect 9864 26250 9916 26256
rect 9864 25832 9916 25838
rect 9864 25774 9916 25780
rect 9772 25696 9824 25702
rect 9772 25638 9824 25644
rect 9876 24954 9904 25774
rect 10152 25362 10180 26823
rect 10244 26761 10272 26930
rect 10230 26752 10286 26761
rect 10230 26687 10286 26696
rect 10232 26308 10284 26314
rect 10232 26250 10284 26256
rect 10140 25356 10192 25362
rect 10140 25298 10192 25304
rect 10152 25129 10180 25298
rect 10138 25120 10194 25129
rect 10138 25055 10194 25064
rect 9864 24948 9916 24954
rect 9864 24890 9916 24896
rect 10048 24744 10100 24750
rect 10048 24686 10100 24692
rect 9496 24608 9548 24614
rect 9496 24550 9548 24556
rect 9680 24268 9732 24274
rect 9680 24210 9732 24216
rect 9692 23769 9720 24210
rect 9956 24064 10008 24070
rect 9956 24006 10008 24012
rect 9678 23760 9734 23769
rect 9678 23695 9680 23704
rect 9732 23695 9734 23704
rect 9680 23666 9732 23672
rect 9404 23656 9456 23662
rect 9404 23598 9456 23604
rect 9416 23186 9444 23598
rect 9404 23180 9456 23186
rect 9404 23122 9456 23128
rect 9864 22976 9916 22982
rect 9864 22918 9916 22924
rect 9404 22636 9456 22642
rect 9404 22578 9456 22584
rect 9416 21554 9444 22578
rect 9680 22568 9732 22574
rect 9680 22510 9732 22516
rect 9692 21690 9720 22510
rect 9772 22024 9824 22030
rect 9772 21966 9824 21972
rect 9784 21690 9812 21966
rect 9680 21684 9732 21690
rect 9680 21626 9732 21632
rect 9772 21684 9824 21690
rect 9772 21626 9824 21632
rect 9404 21548 9456 21554
rect 9404 21490 9456 21496
rect 9416 20262 9444 21490
rect 9680 21480 9732 21486
rect 9680 21422 9732 21428
rect 9496 21140 9548 21146
rect 9496 21082 9548 21088
rect 9508 20942 9536 21082
rect 9496 20936 9548 20942
rect 9496 20878 9548 20884
rect 9404 20256 9456 20262
rect 9404 20198 9456 20204
rect 9416 19990 9444 20198
rect 9404 19984 9456 19990
rect 9404 19926 9456 19932
rect 9048 19306 9260 19334
rect 9232 18358 9260 19306
rect 9508 18834 9536 20878
rect 9496 18828 9548 18834
rect 9496 18770 9548 18776
rect 9220 18352 9272 18358
rect 9220 18294 9272 18300
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 7564 3188 7616 3194
rect 7564 3130 7616 3136
rect 2412 2848 2464 2854
rect 2412 2790 2464 2796
rect 1952 2440 2004 2446
rect 1952 2382 2004 2388
rect 2424 2378 2452 2790
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 5552 2446 5580 3130
rect 8588 3058 8616 9998
rect 9692 6866 9720 21422
rect 9876 20602 9904 22918
rect 9968 20806 9996 24006
rect 10060 23186 10088 24686
rect 10140 24132 10192 24138
rect 10140 24074 10192 24080
rect 10152 23866 10180 24074
rect 10140 23860 10192 23866
rect 10140 23802 10192 23808
rect 10048 23180 10100 23186
rect 10048 23122 10100 23128
rect 9956 20800 10008 20806
rect 9956 20742 10008 20748
rect 9864 20596 9916 20602
rect 9864 20538 9916 20544
rect 9772 20460 9824 20466
rect 9772 20402 9824 20408
rect 9784 20058 9812 20402
rect 9772 20052 9824 20058
rect 9772 19994 9824 20000
rect 10060 10266 10088 23122
rect 10138 22128 10194 22137
rect 10138 22063 10194 22072
rect 10152 22030 10180 22063
rect 10140 22024 10192 22030
rect 10140 21966 10192 21972
rect 10244 21486 10272 26250
rect 10336 25265 10364 29022
rect 10704 29050 10732 29124
rect 10508 29038 10560 29044
rect 10414 28999 10470 29008
rect 10612 29022 10732 29050
rect 10612 28994 10640 29022
rect 10796 28994 10824 29192
rect 10520 28966 10640 28994
rect 10704 28966 10824 28994
rect 10416 28008 10468 28014
rect 10416 27950 10468 27956
rect 10428 27674 10456 27950
rect 10416 27668 10468 27674
rect 10416 27610 10468 27616
rect 10428 26874 10456 27610
rect 10520 27520 10548 28966
rect 10520 27492 10640 27520
rect 10508 27396 10560 27402
rect 10508 27338 10560 27344
rect 10520 27130 10548 27338
rect 10508 27124 10560 27130
rect 10508 27066 10560 27072
rect 10428 26846 10548 26874
rect 10520 26450 10548 26846
rect 10508 26444 10560 26450
rect 10508 26386 10560 26392
rect 10508 25968 10560 25974
rect 10612 25956 10640 27492
rect 10704 26897 10732 28966
rect 10690 26888 10746 26897
rect 10690 26823 10746 26832
rect 10692 26784 10744 26790
rect 10692 26726 10744 26732
rect 10704 26466 10732 26726
rect 10704 26450 10824 26466
rect 10704 26444 10836 26450
rect 10704 26438 10784 26444
rect 10784 26386 10836 26392
rect 10560 25928 10640 25956
rect 10508 25910 10560 25916
rect 10416 25356 10468 25362
rect 10416 25298 10468 25304
rect 10322 25256 10378 25265
rect 10322 25191 10378 25200
rect 10336 24818 10364 25191
rect 10324 24812 10376 24818
rect 10324 24754 10376 24760
rect 10428 24274 10456 25298
rect 10600 25152 10652 25158
rect 10600 25094 10652 25100
rect 10508 24880 10560 24886
rect 10508 24822 10560 24828
rect 10520 24410 10548 24822
rect 10612 24682 10640 25094
rect 10600 24676 10652 24682
rect 10600 24618 10652 24624
rect 10508 24404 10560 24410
rect 10508 24346 10560 24352
rect 10416 24268 10468 24274
rect 10416 24210 10468 24216
rect 10324 22024 10376 22030
rect 10324 21966 10376 21972
rect 10232 21480 10284 21486
rect 10232 21422 10284 21428
rect 10336 21350 10364 21966
rect 10324 21344 10376 21350
rect 10324 21286 10376 21292
rect 10232 21072 10284 21078
rect 10428 21060 10456 24210
rect 10888 23730 10916 30806
rect 10966 30288 11022 30297
rect 11072 30258 11100 37046
rect 11242 36952 11298 36961
rect 11242 36887 11298 36896
rect 11152 36576 11204 36582
rect 11152 36518 11204 36524
rect 11164 36378 11192 36518
rect 11152 36372 11204 36378
rect 11152 36314 11204 36320
rect 11256 35136 11284 36887
rect 11348 36854 11376 37046
rect 11336 36848 11388 36854
rect 11336 36790 11388 36796
rect 11532 36718 11560 37198
rect 11704 37188 11756 37194
rect 11704 37130 11756 37136
rect 11520 36712 11572 36718
rect 11426 36680 11482 36689
rect 11520 36654 11572 36660
rect 11426 36615 11482 36624
rect 11336 36100 11388 36106
rect 11336 36042 11388 36048
rect 11348 36009 11376 36042
rect 11334 36000 11390 36009
rect 11334 35935 11390 35944
rect 11336 35828 11388 35834
rect 11336 35770 11388 35776
rect 11348 35630 11376 35770
rect 11336 35624 11388 35630
rect 11336 35566 11388 35572
rect 11164 35108 11284 35136
rect 11164 35018 11192 35108
rect 11152 35012 11204 35018
rect 11152 34954 11204 34960
rect 11244 35012 11296 35018
rect 11244 34954 11296 34960
rect 11164 33538 11192 34954
rect 11256 34921 11284 34954
rect 11242 34912 11298 34921
rect 11242 34847 11298 34856
rect 11440 34354 11468 36615
rect 11532 35834 11560 36654
rect 11520 35828 11572 35834
rect 11520 35770 11572 35776
rect 11532 35154 11560 35770
rect 11612 35488 11664 35494
rect 11612 35430 11664 35436
rect 11624 35154 11652 35430
rect 11520 35148 11572 35154
rect 11520 35090 11572 35096
rect 11612 35148 11664 35154
rect 11612 35090 11664 35096
rect 11532 34610 11560 35090
rect 11520 34604 11572 34610
rect 11572 34564 11652 34592
rect 11520 34546 11572 34552
rect 11440 34326 11560 34354
rect 11428 34128 11480 34134
rect 11428 34070 11480 34076
rect 11334 33824 11390 33833
rect 11334 33759 11390 33768
rect 11348 33658 11376 33759
rect 11336 33652 11388 33658
rect 11336 33594 11388 33600
rect 11164 33510 11376 33538
rect 11244 33448 11296 33454
rect 11244 33390 11296 33396
rect 11256 32978 11284 33390
rect 11244 32972 11296 32978
rect 11244 32914 11296 32920
rect 11150 32600 11206 32609
rect 11150 32535 11152 32544
rect 11204 32535 11206 32544
rect 11152 32506 11204 32512
rect 11256 32366 11284 32914
rect 11244 32360 11296 32366
rect 11244 32302 11296 32308
rect 11152 32224 11204 32230
rect 11152 32166 11204 32172
rect 10966 30223 10968 30232
rect 11020 30223 11022 30232
rect 11060 30252 11112 30258
rect 10968 30194 11020 30200
rect 11060 30194 11112 30200
rect 11164 30161 11192 32166
rect 11256 31890 11284 32302
rect 11244 31884 11296 31890
rect 11244 31826 11296 31832
rect 11256 31346 11284 31826
rect 11348 31822 11376 33510
rect 11440 31958 11468 34070
rect 11532 32978 11560 34326
rect 11624 34066 11652 34564
rect 11612 34060 11664 34066
rect 11612 34002 11664 34008
rect 11624 33522 11652 34002
rect 11612 33516 11664 33522
rect 11612 33458 11664 33464
rect 11520 32972 11572 32978
rect 11520 32914 11572 32920
rect 11520 32496 11572 32502
rect 11520 32438 11572 32444
rect 11532 32065 11560 32438
rect 11518 32056 11574 32065
rect 11518 31991 11574 32000
rect 11428 31952 11480 31958
rect 11428 31894 11480 31900
rect 11336 31816 11388 31822
rect 11336 31758 11388 31764
rect 11244 31340 11296 31346
rect 11296 31300 11376 31328
rect 11244 31282 11296 31288
rect 11244 31204 11296 31210
rect 11244 31146 11296 31152
rect 11150 30152 11206 30161
rect 11150 30087 11206 30096
rect 11060 30048 11112 30054
rect 11060 29990 11112 29996
rect 11072 29306 11100 29990
rect 11060 29300 11112 29306
rect 11060 29242 11112 29248
rect 11060 29028 11112 29034
rect 11060 28970 11112 28976
rect 11164 28994 11192 30087
rect 11256 29714 11284 31146
rect 11348 30190 11376 31300
rect 11520 30932 11572 30938
rect 11520 30874 11572 30880
rect 11532 30705 11560 30874
rect 11612 30796 11664 30802
rect 11612 30738 11664 30744
rect 11518 30696 11574 30705
rect 11518 30631 11574 30640
rect 11624 30598 11652 30738
rect 11612 30592 11664 30598
rect 11612 30534 11664 30540
rect 11716 30376 11744 37130
rect 11888 36848 11940 36854
rect 11888 36790 11940 36796
rect 11794 34096 11850 34105
rect 11794 34031 11850 34040
rect 11808 33318 11836 34031
rect 11900 33590 11928 36790
rect 12268 36378 12296 39200
rect 13556 39114 13584 39200
rect 13648 39114 13676 39222
rect 13556 39086 13676 39114
rect 13832 37330 13860 39222
rect 15474 39200 15530 39800
rect 16762 39200 16818 39800
rect 18694 39200 18750 39800
rect 20626 39200 20682 39800
rect 21914 39200 21970 39800
rect 23846 39200 23902 39800
rect 25134 39200 25190 39800
rect 27066 39200 27122 39800
rect 28998 39200 29054 39800
rect 30286 39200 30342 39800
rect 32218 39200 32274 39800
rect 33506 39200 33562 39800
rect 35438 39200 35494 39800
rect 37370 39200 37426 39800
rect 38658 39200 38714 39800
rect 12624 37324 12676 37330
rect 12624 37266 12676 37272
rect 13820 37324 13872 37330
rect 13820 37266 13872 37272
rect 12636 36922 12664 37266
rect 13728 37256 13780 37262
rect 13728 37198 13780 37204
rect 12900 37120 12952 37126
rect 12898 37088 12900 37097
rect 12952 37088 12954 37097
rect 12898 37023 12954 37032
rect 13450 37088 13506 37097
rect 13450 37023 13506 37032
rect 12532 36916 12584 36922
rect 12532 36858 12584 36864
rect 12624 36916 12676 36922
rect 12624 36858 12676 36864
rect 12440 36644 12492 36650
rect 12440 36586 12492 36592
rect 12164 36372 12216 36378
rect 12164 36314 12216 36320
rect 12256 36372 12308 36378
rect 12256 36314 12308 36320
rect 12176 36281 12204 36314
rect 12162 36272 12218 36281
rect 12162 36207 12218 36216
rect 12256 36236 12308 36242
rect 12256 36178 12308 36184
rect 12348 36236 12400 36242
rect 12348 36178 12400 36184
rect 12268 36038 12296 36178
rect 12360 36106 12388 36178
rect 12452 36106 12480 36586
rect 12544 36417 12572 36858
rect 13464 36854 13492 37023
rect 13452 36848 13504 36854
rect 13452 36790 13504 36796
rect 13740 36786 13768 37198
rect 14648 37188 14700 37194
rect 14648 37130 14700 37136
rect 13728 36780 13780 36786
rect 13728 36722 13780 36728
rect 12530 36408 12586 36417
rect 12530 36343 12586 36352
rect 13268 36372 13320 36378
rect 13268 36314 13320 36320
rect 13280 36281 13308 36314
rect 13266 36272 13322 36281
rect 13740 36242 13768 36722
rect 13266 36207 13322 36216
rect 13728 36236 13780 36242
rect 13728 36178 13780 36184
rect 12348 36100 12400 36106
rect 12348 36042 12400 36048
rect 12440 36100 12492 36106
rect 12440 36042 12492 36048
rect 13268 36100 13320 36106
rect 13268 36042 13320 36048
rect 12256 36032 12308 36038
rect 12256 35974 12308 35980
rect 13280 35986 13308 36042
rect 13280 35958 13400 35986
rect 12714 35864 12770 35873
rect 12714 35799 12770 35808
rect 12728 35630 12756 35799
rect 13176 35760 13228 35766
rect 13176 35702 13228 35708
rect 12716 35624 12768 35630
rect 12716 35566 12768 35572
rect 12808 35624 12860 35630
rect 12808 35566 12860 35572
rect 12820 35494 12848 35566
rect 12808 35488 12860 35494
rect 12808 35430 12860 35436
rect 12254 35320 12310 35329
rect 12254 35255 12256 35264
rect 12308 35255 12310 35264
rect 13082 35320 13138 35329
rect 13082 35255 13138 35264
rect 12256 35226 12308 35232
rect 12716 35148 12768 35154
rect 12716 35090 12768 35096
rect 12440 35012 12492 35018
rect 12176 34972 12440 35000
rect 12072 34536 12124 34542
rect 12072 34478 12124 34484
rect 11888 33584 11940 33590
rect 11888 33526 11940 33532
rect 11796 33312 11848 33318
rect 11796 33254 11848 33260
rect 11796 32768 11848 32774
rect 11796 32710 11848 32716
rect 11888 32768 11940 32774
rect 11888 32710 11940 32716
rect 11808 31890 11836 32710
rect 11900 32609 11928 32710
rect 11886 32600 11942 32609
rect 11886 32535 11942 32544
rect 11888 32292 11940 32298
rect 11888 32234 11940 32240
rect 11796 31884 11848 31890
rect 11796 31826 11848 31832
rect 11900 30410 11928 32234
rect 11980 31272 12032 31278
rect 11980 31214 12032 31220
rect 11992 30938 12020 31214
rect 12084 31090 12112 34478
rect 12176 31754 12204 34972
rect 12440 34954 12492 34960
rect 12728 34950 12756 35090
rect 12716 34944 12768 34950
rect 12716 34886 12768 34892
rect 12714 34776 12770 34785
rect 12714 34711 12716 34720
rect 12768 34711 12770 34720
rect 12808 34740 12860 34746
rect 12716 34682 12768 34688
rect 12808 34682 12860 34688
rect 12256 34672 12308 34678
rect 12256 34614 12308 34620
rect 12440 34672 12492 34678
rect 12820 34649 12848 34682
rect 12440 34614 12492 34620
rect 12806 34640 12862 34649
rect 12268 34513 12296 34614
rect 12348 34536 12400 34542
rect 12254 34504 12310 34513
rect 12348 34478 12400 34484
rect 12254 34439 12310 34448
rect 12360 34377 12388 34478
rect 12346 34368 12402 34377
rect 12346 34303 12402 34312
rect 12346 34232 12402 34241
rect 12256 34196 12308 34202
rect 12346 34167 12348 34176
rect 12256 34138 12308 34144
rect 12400 34167 12402 34176
rect 12348 34138 12400 34144
rect 12268 34066 12296 34138
rect 12256 34060 12308 34066
rect 12256 34002 12308 34008
rect 12452 33130 12480 34614
rect 12806 34575 12862 34584
rect 12530 34232 12586 34241
rect 12530 34167 12586 34176
rect 12544 34066 12572 34167
rect 12532 34060 12584 34066
rect 12532 34002 12584 34008
rect 12624 34060 12676 34066
rect 12624 34002 12676 34008
rect 12636 33561 12664 34002
rect 12728 33918 12940 33946
rect 12728 33862 12756 33918
rect 12716 33856 12768 33862
rect 12716 33798 12768 33804
rect 12912 33561 12940 33918
rect 12622 33552 12678 33561
rect 12622 33487 12678 33496
rect 12898 33552 12954 33561
rect 12898 33487 12954 33496
rect 12716 33448 12768 33454
rect 12716 33390 12768 33396
rect 12268 33114 12388 33130
rect 12268 33108 12400 33114
rect 12268 33102 12348 33108
rect 12268 32337 12296 33102
rect 12452 33102 12572 33130
rect 12348 33050 12400 33056
rect 12440 32836 12492 32842
rect 12440 32778 12492 32784
rect 12254 32328 12310 32337
rect 12254 32263 12310 32272
rect 12254 31920 12310 31929
rect 12254 31855 12310 31864
rect 12164 31748 12216 31754
rect 12164 31690 12216 31696
rect 12268 31686 12296 31855
rect 12256 31680 12308 31686
rect 12256 31622 12308 31628
rect 12164 31476 12216 31482
rect 12164 31418 12216 31424
rect 12176 31385 12204 31418
rect 12162 31376 12218 31385
rect 12162 31311 12218 31320
rect 12084 31062 12204 31090
rect 11980 30932 12032 30938
rect 11980 30874 12032 30880
rect 11900 30382 12020 30410
rect 11440 30348 11744 30376
rect 11336 30184 11388 30190
rect 11336 30126 11388 30132
rect 11334 30016 11390 30025
rect 11334 29951 11390 29960
rect 11348 29850 11376 29951
rect 11336 29844 11388 29850
rect 11336 29786 11388 29792
rect 11244 29708 11296 29714
rect 11244 29650 11296 29656
rect 11242 29608 11298 29617
rect 11242 29543 11298 29552
rect 11256 29238 11284 29543
rect 11244 29232 11296 29238
rect 11244 29174 11296 29180
rect 11336 29028 11388 29034
rect 10968 28416 11020 28422
rect 10968 28358 11020 28364
rect 10980 26994 11008 28358
rect 10968 26988 11020 26994
rect 10968 26930 11020 26936
rect 10980 24206 11008 26930
rect 11072 25809 11100 28970
rect 11164 28966 11284 28994
rect 11336 28970 11388 28976
rect 11150 28656 11206 28665
rect 11150 28591 11206 28600
rect 11164 28490 11192 28591
rect 11152 28484 11204 28490
rect 11152 28426 11204 28432
rect 11256 28014 11284 28966
rect 11348 28098 11376 28970
rect 11440 28626 11468 30348
rect 11992 30326 12020 30382
rect 11888 30320 11940 30326
rect 11888 30262 11940 30268
rect 11980 30320 12032 30326
rect 11980 30262 12032 30268
rect 11612 30252 11664 30258
rect 11612 30194 11664 30200
rect 11624 29578 11652 30194
rect 11704 30184 11756 30190
rect 11704 30126 11756 30132
rect 11716 29714 11744 30126
rect 11704 29708 11756 29714
rect 11704 29650 11756 29656
rect 11612 29572 11664 29578
rect 11612 29514 11664 29520
rect 11518 29336 11574 29345
rect 11518 29271 11574 29280
rect 11532 29170 11560 29271
rect 11520 29164 11572 29170
rect 11520 29106 11572 29112
rect 11624 28801 11652 29514
rect 11716 29102 11744 29650
rect 11796 29572 11848 29578
rect 11796 29514 11848 29520
rect 11704 29096 11756 29102
rect 11704 29038 11756 29044
rect 11610 28792 11666 28801
rect 11532 28750 11610 28778
rect 11428 28620 11480 28626
rect 11428 28562 11480 28568
rect 11348 28070 11468 28098
rect 11244 28008 11296 28014
rect 11244 27950 11296 27956
rect 11336 28008 11388 28014
rect 11336 27950 11388 27956
rect 11152 27940 11204 27946
rect 11152 27882 11204 27888
rect 11164 27062 11192 27882
rect 11152 27056 11204 27062
rect 11204 27016 11284 27044
rect 11152 26998 11204 27004
rect 11152 26920 11204 26926
rect 11152 26862 11204 26868
rect 11164 25974 11192 26862
rect 11152 25968 11204 25974
rect 11152 25910 11204 25916
rect 11058 25800 11114 25809
rect 11164 25770 11192 25910
rect 11058 25735 11114 25744
rect 11152 25764 11204 25770
rect 11152 25706 11204 25712
rect 10968 24200 11020 24206
rect 10968 24142 11020 24148
rect 10966 23896 11022 23905
rect 10966 23831 10968 23840
rect 11020 23831 11022 23840
rect 10968 23802 11020 23808
rect 10876 23724 10928 23730
rect 10876 23666 10928 23672
rect 11060 23724 11112 23730
rect 11060 23666 11112 23672
rect 10888 23594 10916 23666
rect 11072 23633 11100 23666
rect 11058 23624 11114 23633
rect 10876 23588 10928 23594
rect 11058 23559 11114 23568
rect 10876 23530 10928 23536
rect 11256 23322 11284 27016
rect 11348 26450 11376 27950
rect 11440 27690 11468 28070
rect 11532 27878 11560 28750
rect 11610 28727 11666 28736
rect 11716 28626 11744 29038
rect 11808 29034 11836 29514
rect 11796 29028 11848 29034
rect 11796 28970 11848 28976
rect 11796 28756 11848 28762
rect 11796 28698 11848 28704
rect 11704 28620 11756 28626
rect 11624 28580 11704 28608
rect 11624 28082 11652 28580
rect 11704 28562 11756 28568
rect 11702 28520 11758 28529
rect 11702 28455 11758 28464
rect 11716 28422 11744 28455
rect 11704 28416 11756 28422
rect 11808 28393 11836 28698
rect 11704 28358 11756 28364
rect 11794 28384 11850 28393
rect 11794 28319 11850 28328
rect 11612 28076 11664 28082
rect 11612 28018 11664 28024
rect 11520 27872 11572 27878
rect 11520 27814 11572 27820
rect 11440 27662 11560 27690
rect 11428 27532 11480 27538
rect 11428 27474 11480 27480
rect 11336 26444 11388 26450
rect 11336 26386 11388 26392
rect 11348 26246 11376 26386
rect 11336 26240 11388 26246
rect 11336 26182 11388 26188
rect 11440 24138 11468 27474
rect 11532 27402 11560 27662
rect 11520 27396 11572 27402
rect 11520 27338 11572 27344
rect 11336 24132 11388 24138
rect 11336 24074 11388 24080
rect 11428 24132 11480 24138
rect 11428 24074 11480 24080
rect 11244 23316 11296 23322
rect 11244 23258 11296 23264
rect 10876 23248 10928 23254
rect 10876 23190 10928 23196
rect 10784 22976 10836 22982
rect 10784 22918 10836 22924
rect 10692 22568 10744 22574
rect 10692 22510 10744 22516
rect 10704 21622 10732 22510
rect 10692 21616 10744 21622
rect 10692 21558 10744 21564
rect 10796 21146 10824 22918
rect 10888 22642 10916 23190
rect 10876 22636 10928 22642
rect 10876 22578 10928 22584
rect 10784 21140 10836 21146
rect 10784 21082 10836 21088
rect 10284 21032 10456 21060
rect 10232 21014 10284 21020
rect 10140 19848 10192 19854
rect 10140 19790 10192 19796
rect 10152 18970 10180 19790
rect 10140 18964 10192 18970
rect 10140 18906 10192 18912
rect 10244 18290 10272 21014
rect 10784 20868 10836 20874
rect 10784 20810 10836 20816
rect 10796 20398 10824 20810
rect 10888 20534 10916 22578
rect 11060 22432 11112 22438
rect 11060 22374 11112 22380
rect 10968 21888 11020 21894
rect 10968 21830 11020 21836
rect 10980 21622 11008 21830
rect 10968 21616 11020 21622
rect 10968 21558 11020 21564
rect 11072 21486 11100 22374
rect 11256 22166 11284 23258
rect 11244 22160 11296 22166
rect 11244 22102 11296 22108
rect 11152 21956 11204 21962
rect 11152 21898 11204 21904
rect 11060 21480 11112 21486
rect 11060 21422 11112 21428
rect 10876 20528 10928 20534
rect 10876 20470 10928 20476
rect 11060 20528 11112 20534
rect 11060 20470 11112 20476
rect 10784 20392 10836 20398
rect 10784 20334 10836 20340
rect 10888 19854 10916 20470
rect 10876 19848 10928 19854
rect 10876 19790 10928 19796
rect 10888 19514 10916 19790
rect 11072 19514 11100 20470
rect 11164 20058 11192 21898
rect 11244 21412 11296 21418
rect 11244 21354 11296 21360
rect 11256 20398 11284 21354
rect 11244 20392 11296 20398
rect 11244 20334 11296 20340
rect 11152 20052 11204 20058
rect 11152 19994 11204 20000
rect 10876 19508 10928 19514
rect 10876 19450 10928 19456
rect 11060 19508 11112 19514
rect 11060 19450 11112 19456
rect 11348 19174 11376 24074
rect 11440 19922 11468 24074
rect 11532 23186 11560 27338
rect 11796 26444 11848 26450
rect 11796 26386 11848 26392
rect 11808 26042 11836 26386
rect 11900 26042 11928 30262
rect 11992 29345 12020 30262
rect 12072 30184 12124 30190
rect 12072 30126 12124 30132
rect 11978 29336 12034 29345
rect 11978 29271 12034 29280
rect 11796 26036 11848 26042
rect 11796 25978 11848 25984
rect 11888 26036 11940 26042
rect 11888 25978 11940 25984
rect 11992 25514 12020 29271
rect 12084 27130 12112 30126
rect 12176 27606 12204 31062
rect 12346 30968 12402 30977
rect 12346 30903 12402 30912
rect 12360 30802 12388 30903
rect 12348 30796 12400 30802
rect 12348 30738 12400 30744
rect 12256 28552 12308 28558
rect 12256 28494 12308 28500
rect 12268 27713 12296 28494
rect 12360 28121 12388 30738
rect 12346 28112 12402 28121
rect 12346 28047 12402 28056
rect 12348 27872 12400 27878
rect 12348 27814 12400 27820
rect 12254 27704 12310 27713
rect 12254 27639 12310 27648
rect 12164 27600 12216 27606
rect 12164 27542 12216 27548
rect 12072 27124 12124 27130
rect 12072 27066 12124 27072
rect 12072 26852 12124 26858
rect 12072 26794 12124 26800
rect 11716 25486 12020 25514
rect 11612 25356 11664 25362
rect 11612 25298 11664 25304
rect 11624 24954 11652 25298
rect 11612 24948 11664 24954
rect 11612 24890 11664 24896
rect 11612 23520 11664 23526
rect 11612 23462 11664 23468
rect 11520 23180 11572 23186
rect 11520 23122 11572 23128
rect 11624 22710 11652 23462
rect 11612 22704 11664 22710
rect 11612 22646 11664 22652
rect 11716 22137 11744 25486
rect 11796 25220 11848 25226
rect 11796 25162 11848 25168
rect 11808 24614 11836 25162
rect 12084 25158 12112 26794
rect 12164 25764 12216 25770
rect 12164 25706 12216 25712
rect 12176 25430 12204 25706
rect 12164 25424 12216 25430
rect 12164 25366 12216 25372
rect 12072 25152 12124 25158
rect 12256 25152 12308 25158
rect 12072 25094 12124 25100
rect 12254 25120 12256 25129
rect 12308 25120 12310 25129
rect 11888 24880 11940 24886
rect 11888 24822 11940 24828
rect 11796 24608 11848 24614
rect 11796 24550 11848 24556
rect 11900 24342 11928 24822
rect 11888 24336 11940 24342
rect 11888 24278 11940 24284
rect 11978 23760 12034 23769
rect 11978 23695 11980 23704
rect 12032 23695 12034 23704
rect 11980 23666 12032 23672
rect 11886 23624 11942 23633
rect 11886 23559 11888 23568
rect 11940 23559 11942 23568
rect 11888 23530 11940 23536
rect 11980 23520 12032 23526
rect 11980 23462 12032 23468
rect 11888 23180 11940 23186
rect 11888 23122 11940 23128
rect 11796 23044 11848 23050
rect 11796 22986 11848 22992
rect 11702 22128 11758 22137
rect 11702 22063 11758 22072
rect 11808 21894 11836 22986
rect 11900 22574 11928 23122
rect 11888 22568 11940 22574
rect 11888 22510 11940 22516
rect 11992 21894 12020 23462
rect 11796 21888 11848 21894
rect 11796 21830 11848 21836
rect 11980 21888 12032 21894
rect 11980 21830 12032 21836
rect 11980 21480 12032 21486
rect 11980 21422 12032 21428
rect 11992 20806 12020 21422
rect 11980 20800 12032 20806
rect 11980 20742 12032 20748
rect 11428 19916 11480 19922
rect 11428 19858 11480 19864
rect 11428 19780 11480 19786
rect 11428 19722 11480 19728
rect 11440 19310 11468 19722
rect 11992 19514 12020 20742
rect 12084 20534 12112 25094
rect 12254 25055 12310 25064
rect 12164 24948 12216 24954
rect 12164 24890 12216 24896
rect 12176 24750 12204 24890
rect 12164 24744 12216 24750
rect 12164 24686 12216 24692
rect 12164 24268 12216 24274
rect 12164 24210 12216 24216
rect 12176 22710 12204 24210
rect 12256 24132 12308 24138
rect 12256 24074 12308 24080
rect 12268 23662 12296 24074
rect 12256 23656 12308 23662
rect 12256 23598 12308 23604
rect 12164 22704 12216 22710
rect 12164 22646 12216 22652
rect 12256 22500 12308 22506
rect 12256 22442 12308 22448
rect 12268 22137 12296 22442
rect 12254 22128 12310 22137
rect 12254 22063 12310 22072
rect 12360 20602 12388 27814
rect 12452 27538 12480 32778
rect 12544 28393 12572 33102
rect 12624 32496 12676 32502
rect 12624 32438 12676 32444
rect 12636 32337 12664 32438
rect 12622 32328 12678 32337
rect 12622 32263 12678 32272
rect 12624 32224 12676 32230
rect 12624 32166 12676 32172
rect 12636 31929 12664 32166
rect 12622 31920 12678 31929
rect 12622 31855 12678 31864
rect 12622 31784 12678 31793
rect 12622 31719 12678 31728
rect 12636 29866 12664 31719
rect 12728 30938 12756 33390
rect 12808 32904 12860 32910
rect 12808 32846 12860 32852
rect 12820 32201 12848 32846
rect 13096 32842 13124 35255
rect 13188 35222 13216 35702
rect 13176 35216 13228 35222
rect 13176 35158 13228 35164
rect 13188 34542 13216 35158
rect 13176 34536 13228 34542
rect 13176 34478 13228 34484
rect 13268 33856 13320 33862
rect 13188 33816 13268 33844
rect 13084 32836 13136 32842
rect 13084 32778 13136 32784
rect 13188 32502 13216 33816
rect 13268 33798 13320 33804
rect 13268 33040 13320 33046
rect 13268 32982 13320 32988
rect 13176 32496 13228 32502
rect 13174 32464 13176 32473
rect 13228 32464 13230 32473
rect 13174 32399 13230 32408
rect 13280 32280 13308 32982
rect 13372 32450 13400 35958
rect 13740 35698 13768 36178
rect 14660 36174 14688 37130
rect 15488 37126 15516 39200
rect 16672 37800 16724 37806
rect 16672 37742 16724 37748
rect 15844 37256 15896 37262
rect 15844 37198 15896 37204
rect 15200 37120 15252 37126
rect 15200 37062 15252 37068
rect 15476 37120 15528 37126
rect 15476 37062 15528 37068
rect 15752 37120 15804 37126
rect 15752 37062 15804 37068
rect 15016 36780 15068 36786
rect 15016 36722 15068 36728
rect 15028 36666 15056 36722
rect 14844 36638 15056 36666
rect 14648 36168 14700 36174
rect 14648 36110 14700 36116
rect 14464 36032 14516 36038
rect 14464 35974 14516 35980
rect 14740 36032 14792 36038
rect 14740 35974 14792 35980
rect 14476 35834 14504 35974
rect 14464 35828 14516 35834
rect 14464 35770 14516 35776
rect 13728 35692 13780 35698
rect 13728 35634 13780 35640
rect 14188 35692 14240 35698
rect 14188 35634 14240 35640
rect 14004 35556 14056 35562
rect 14004 35498 14056 35504
rect 14016 35465 14044 35498
rect 14200 35465 14228 35634
rect 14002 35456 14058 35465
rect 14002 35391 14058 35400
rect 14186 35456 14242 35465
rect 14186 35391 14242 35400
rect 13912 35080 13964 35086
rect 13912 35022 13964 35028
rect 13818 34504 13874 34513
rect 13818 34439 13874 34448
rect 13452 33856 13504 33862
rect 13452 33798 13504 33804
rect 13464 33318 13492 33798
rect 13726 33688 13782 33697
rect 13726 33623 13782 33632
rect 13740 33522 13768 33623
rect 13728 33516 13780 33522
rect 13728 33458 13780 33464
rect 13452 33312 13504 33318
rect 13452 33254 13504 33260
rect 13728 32972 13780 32978
rect 13728 32914 13780 32920
rect 13740 32858 13768 32914
rect 13464 32830 13768 32858
rect 13464 32774 13492 32830
rect 13452 32768 13504 32774
rect 13452 32710 13504 32716
rect 13636 32768 13688 32774
rect 13636 32710 13688 32716
rect 13648 32570 13676 32710
rect 13832 32609 13860 34439
rect 13924 33912 13952 35022
rect 14004 35012 14056 35018
rect 14004 34954 14056 34960
rect 14016 34649 14044 34954
rect 14096 34944 14148 34950
rect 14096 34886 14148 34892
rect 14002 34640 14058 34649
rect 14002 34575 14058 34584
rect 13924 33884 14044 33912
rect 13910 33824 13966 33833
rect 13910 33759 13966 33768
rect 13924 33522 13952 33759
rect 13912 33516 13964 33522
rect 13912 33458 13964 33464
rect 13912 33040 13964 33046
rect 13912 32982 13964 32988
rect 13818 32600 13874 32609
rect 13636 32564 13688 32570
rect 13818 32535 13874 32544
rect 13636 32506 13688 32512
rect 13372 32422 13676 32450
rect 13544 32292 13596 32298
rect 13280 32252 13544 32280
rect 12992 32224 13044 32230
rect 12806 32192 12862 32201
rect 12806 32127 12862 32136
rect 12912 32184 12992 32212
rect 12716 30932 12768 30938
rect 12716 30874 12768 30880
rect 12808 30864 12860 30870
rect 12808 30806 12860 30812
rect 12820 30734 12848 30806
rect 12808 30728 12860 30734
rect 12808 30670 12860 30676
rect 12716 30660 12768 30666
rect 12716 30602 12768 30608
rect 12728 30025 12756 30602
rect 12714 30016 12770 30025
rect 12714 29951 12770 29960
rect 12806 29880 12862 29889
rect 12636 29838 12756 29866
rect 12624 29776 12676 29782
rect 12624 29718 12676 29724
rect 12530 28384 12586 28393
rect 12530 28319 12586 28328
rect 12532 28212 12584 28218
rect 12532 28154 12584 28160
rect 12544 28121 12572 28154
rect 12530 28112 12586 28121
rect 12530 28047 12586 28056
rect 12440 27532 12492 27538
rect 12440 27474 12492 27480
rect 12532 27328 12584 27334
rect 12532 27270 12584 27276
rect 12440 27056 12492 27062
rect 12440 26998 12492 27004
rect 12452 26586 12480 26998
rect 12544 26897 12572 27270
rect 12530 26888 12586 26897
rect 12530 26823 12586 26832
rect 12532 26784 12584 26790
rect 12532 26726 12584 26732
rect 12544 26586 12572 26726
rect 12440 26580 12492 26586
rect 12440 26522 12492 26528
rect 12532 26580 12584 26586
rect 12532 26522 12584 26528
rect 12438 26480 12494 26489
rect 12438 26415 12494 26424
rect 12452 25378 12480 26415
rect 12544 26081 12572 26522
rect 12636 26234 12664 29718
rect 12728 27334 12756 29838
rect 12806 29815 12862 29824
rect 12820 28506 12848 29815
rect 12912 28642 12940 32184
rect 12992 32166 13044 32172
rect 13084 31816 13136 31822
rect 13084 31758 13136 31764
rect 13096 31385 13124 31758
rect 13176 31748 13228 31754
rect 13176 31690 13228 31696
rect 13188 31414 13216 31690
rect 13176 31408 13228 31414
rect 13082 31376 13138 31385
rect 13176 31350 13228 31356
rect 13082 31311 13138 31320
rect 13096 30734 13124 31311
rect 13084 30728 13136 30734
rect 13084 30670 13136 30676
rect 13084 30252 13136 30258
rect 13084 30194 13136 30200
rect 13096 29850 13124 30194
rect 13176 30048 13228 30054
rect 13176 29990 13228 29996
rect 13084 29844 13136 29850
rect 13084 29786 13136 29792
rect 13188 29578 13216 29990
rect 13280 29714 13308 32252
rect 13544 32234 13596 32240
rect 13648 32178 13676 32422
rect 13728 32360 13780 32366
rect 13728 32302 13780 32308
rect 13556 32150 13676 32178
rect 13360 31884 13412 31890
rect 13360 31826 13412 31832
rect 13372 31142 13400 31826
rect 13556 31754 13584 32150
rect 13636 32020 13688 32026
rect 13636 31962 13688 31968
rect 13544 31748 13596 31754
rect 13544 31690 13596 31696
rect 13452 31680 13504 31686
rect 13452 31622 13504 31628
rect 13464 31396 13492 31622
rect 13544 31408 13596 31414
rect 13464 31368 13544 31396
rect 13544 31350 13596 31356
rect 13360 31136 13412 31142
rect 13360 31078 13412 31084
rect 13452 30796 13504 30802
rect 13452 30738 13504 30744
rect 13464 30122 13492 30738
rect 13452 30116 13504 30122
rect 13452 30058 13504 30064
rect 13464 29782 13492 30058
rect 13452 29776 13504 29782
rect 13452 29718 13504 29724
rect 13268 29708 13320 29714
rect 13268 29650 13320 29656
rect 13176 29572 13228 29578
rect 13176 29514 13228 29520
rect 13544 29232 13596 29238
rect 13544 29174 13596 29180
rect 13176 29096 13228 29102
rect 13176 29038 13228 29044
rect 12912 28614 13032 28642
rect 13004 28558 13032 28614
rect 12992 28552 13044 28558
rect 12820 28478 12940 28506
rect 12992 28494 13044 28500
rect 13188 28490 13216 29038
rect 13268 28552 13320 28558
rect 13268 28494 13320 28500
rect 12808 28416 12860 28422
rect 12808 28358 12860 28364
rect 12820 28121 12848 28358
rect 12806 28112 12862 28121
rect 12806 28047 12862 28056
rect 12808 27532 12860 27538
rect 12808 27474 12860 27480
rect 12716 27328 12768 27334
rect 12716 27270 12768 27276
rect 12716 26580 12768 26586
rect 12716 26522 12768 26528
rect 12728 26382 12756 26522
rect 12716 26376 12768 26382
rect 12716 26318 12768 26324
rect 12636 26206 12756 26234
rect 12530 26072 12586 26081
rect 12530 26007 12586 26016
rect 12532 25968 12584 25974
rect 12532 25910 12584 25916
rect 12544 25498 12572 25910
rect 12728 25702 12756 26206
rect 12716 25696 12768 25702
rect 12716 25638 12768 25644
rect 12532 25492 12584 25498
rect 12532 25434 12584 25440
rect 12624 25492 12676 25498
rect 12624 25434 12676 25440
rect 12452 25350 12572 25378
rect 12440 25220 12492 25226
rect 12440 25162 12492 25168
rect 12452 23866 12480 25162
rect 12544 24970 12572 25350
rect 12636 25158 12664 25434
rect 12728 25158 12756 25638
rect 12624 25152 12676 25158
rect 12624 25094 12676 25100
rect 12716 25152 12768 25158
rect 12716 25094 12768 25100
rect 12544 24942 12756 24970
rect 12624 24880 12676 24886
rect 12624 24822 12676 24828
rect 12532 24812 12584 24818
rect 12532 24754 12584 24760
rect 12440 23860 12492 23866
rect 12440 23802 12492 23808
rect 12440 23656 12492 23662
rect 12440 23598 12492 23604
rect 12452 22234 12480 23598
rect 12544 22778 12572 24754
rect 12636 24342 12664 24822
rect 12624 24336 12676 24342
rect 12624 24278 12676 24284
rect 12728 23905 12756 24942
rect 12714 23896 12770 23905
rect 12714 23831 12770 23840
rect 12716 23792 12768 23798
rect 12716 23734 12768 23740
rect 12622 23624 12678 23633
rect 12622 23559 12678 23568
rect 12636 23526 12664 23559
rect 12624 23520 12676 23526
rect 12624 23462 12676 23468
rect 12624 22976 12676 22982
rect 12624 22918 12676 22924
rect 12532 22772 12584 22778
rect 12532 22714 12584 22720
rect 12440 22228 12492 22234
rect 12440 22170 12492 22176
rect 12636 22166 12664 22918
rect 12728 22778 12756 23734
rect 12820 23254 12848 27474
rect 12912 27470 12940 28478
rect 13176 28484 13228 28490
rect 13176 28426 13228 28432
rect 13280 28370 13308 28494
rect 13188 28342 13308 28370
rect 13360 28416 13412 28422
rect 13360 28358 13412 28364
rect 13084 27872 13136 27878
rect 13084 27814 13136 27820
rect 12992 27668 13044 27674
rect 12992 27610 13044 27616
rect 12900 27464 12952 27470
rect 12900 27406 12952 27412
rect 12808 23248 12860 23254
rect 12808 23190 12860 23196
rect 12912 23100 12940 27406
rect 13004 24154 13032 27610
rect 13096 27402 13124 27814
rect 13084 27396 13136 27402
rect 13084 27338 13136 27344
rect 13084 26784 13136 26790
rect 13084 26726 13136 26732
rect 13096 26518 13124 26726
rect 13084 26512 13136 26518
rect 13084 26454 13136 26460
rect 13096 26314 13124 26454
rect 13084 26308 13136 26314
rect 13084 26250 13136 26256
rect 13004 24138 13124 24154
rect 13004 24132 13136 24138
rect 13004 24126 13084 24132
rect 13084 24074 13136 24080
rect 12820 23072 12940 23100
rect 12716 22772 12768 22778
rect 12716 22714 12768 22720
rect 12624 22160 12676 22166
rect 12624 22102 12676 22108
rect 12820 21570 12848 23072
rect 12900 22432 12952 22438
rect 12900 22374 12952 22380
rect 12912 21978 12940 22374
rect 12912 21962 13032 21978
rect 12912 21956 13044 21962
rect 12912 21950 12992 21956
rect 12992 21898 13044 21904
rect 12820 21542 13032 21570
rect 12440 21480 12492 21486
rect 12440 21422 12492 21428
rect 12452 21010 12480 21422
rect 12808 21412 12860 21418
rect 12808 21354 12860 21360
rect 12820 21078 12848 21354
rect 12808 21072 12860 21078
rect 12808 21014 12860 21020
rect 12440 21004 12492 21010
rect 12440 20946 12492 20952
rect 12900 20936 12952 20942
rect 12900 20878 12952 20884
rect 12624 20868 12676 20874
rect 12624 20810 12676 20816
rect 12348 20596 12400 20602
rect 12348 20538 12400 20544
rect 12072 20528 12124 20534
rect 12072 20470 12124 20476
rect 12636 19922 12664 20810
rect 12808 20528 12860 20534
rect 12808 20470 12860 20476
rect 12624 19916 12676 19922
rect 12624 19858 12676 19864
rect 11980 19508 12032 19514
rect 11980 19450 12032 19456
rect 12636 19378 12664 19858
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 11428 19304 11480 19310
rect 11428 19246 11480 19252
rect 11336 19168 11388 19174
rect 11336 19110 11388 19116
rect 12636 18970 12664 19314
rect 12624 18964 12676 18970
rect 12624 18906 12676 18912
rect 11612 18828 11664 18834
rect 11612 18770 11664 18776
rect 11520 18760 11572 18766
rect 11520 18702 11572 18708
rect 11532 18630 11560 18702
rect 11624 18630 11652 18770
rect 11520 18624 11572 18630
rect 11520 18566 11572 18572
rect 11612 18624 11664 18630
rect 11612 18566 11664 18572
rect 10232 18284 10284 18290
rect 10232 18226 10284 18232
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 8312 2446 8340 2790
rect 8588 2514 8616 2994
rect 11532 2922 11560 18566
rect 12820 18426 12848 20470
rect 12912 18970 12940 20878
rect 13004 19242 13032 21542
rect 13188 21026 13216 28342
rect 13372 27402 13400 28358
rect 13268 27396 13320 27402
rect 13268 27338 13320 27344
rect 13360 27396 13412 27402
rect 13360 27338 13412 27344
rect 13280 24138 13308 27338
rect 13452 27328 13504 27334
rect 13452 27270 13504 27276
rect 13360 26308 13412 26314
rect 13360 26250 13412 26256
rect 13372 24721 13400 26250
rect 13464 25974 13492 27270
rect 13452 25968 13504 25974
rect 13452 25910 13504 25916
rect 13452 25764 13504 25770
rect 13452 25706 13504 25712
rect 13358 24712 13414 24721
rect 13358 24647 13414 24656
rect 13268 24132 13320 24138
rect 13320 24092 13400 24120
rect 13268 24074 13320 24080
rect 13268 22772 13320 22778
rect 13268 22714 13320 22720
rect 13280 21146 13308 22714
rect 13268 21140 13320 21146
rect 13268 21082 13320 21088
rect 13084 21004 13136 21010
rect 13188 20998 13308 21026
rect 13084 20946 13136 20952
rect 13096 19786 13124 20946
rect 13176 20868 13228 20874
rect 13176 20810 13228 20816
rect 13084 19780 13136 19786
rect 13084 19722 13136 19728
rect 12992 19236 13044 19242
rect 12992 19178 13044 19184
rect 12900 18964 12952 18970
rect 12900 18906 12952 18912
rect 12992 18624 13044 18630
rect 12992 18566 13044 18572
rect 12808 18420 12860 18426
rect 12808 18362 12860 18368
rect 13004 17882 13032 18566
rect 12992 17876 13044 17882
rect 12992 17818 13044 17824
rect 13096 10810 13124 19722
rect 13188 18426 13216 20810
rect 13280 20534 13308 20998
rect 13268 20528 13320 20534
rect 13268 20470 13320 20476
rect 13268 20324 13320 20330
rect 13268 20266 13320 20272
rect 13176 18420 13228 18426
rect 13176 18362 13228 18368
rect 13280 13530 13308 20266
rect 13372 19990 13400 24092
rect 13464 23798 13492 25706
rect 13556 24070 13584 29174
rect 13648 28665 13676 31962
rect 13740 31346 13768 32302
rect 13728 31340 13780 31346
rect 13728 31282 13780 31288
rect 13740 30870 13768 31282
rect 13728 30864 13780 30870
rect 13728 30806 13780 30812
rect 13728 30048 13780 30054
rect 13728 29990 13780 29996
rect 13740 29238 13768 29990
rect 13820 29708 13872 29714
rect 13820 29650 13872 29656
rect 13728 29232 13780 29238
rect 13728 29174 13780 29180
rect 13634 28656 13690 28665
rect 13634 28591 13690 28600
rect 13728 28416 13780 28422
rect 13728 28358 13780 28364
rect 13636 27940 13688 27946
rect 13636 27882 13688 27888
rect 13544 24064 13596 24070
rect 13544 24006 13596 24012
rect 13452 23792 13504 23798
rect 13452 23734 13504 23740
rect 13544 23792 13596 23798
rect 13544 23734 13596 23740
rect 13450 23216 13506 23225
rect 13450 23151 13506 23160
rect 13464 23118 13492 23151
rect 13452 23112 13504 23118
rect 13452 23054 13504 23060
rect 13464 22778 13492 23054
rect 13452 22772 13504 22778
rect 13452 22714 13504 22720
rect 13556 20602 13584 23734
rect 13648 22098 13676 27882
rect 13740 27062 13768 28358
rect 13728 27056 13780 27062
rect 13728 26998 13780 27004
rect 13728 26308 13780 26314
rect 13728 26250 13780 26256
rect 13740 25226 13768 26250
rect 13728 25220 13780 25226
rect 13728 25162 13780 25168
rect 13740 24410 13768 25162
rect 13832 24818 13860 29650
rect 13924 29646 13952 32982
rect 14016 30977 14044 33884
rect 14108 32502 14136 34886
rect 14096 32496 14148 32502
rect 14096 32438 14148 32444
rect 14096 31816 14148 31822
rect 14096 31758 14148 31764
rect 14002 30968 14058 30977
rect 14002 30903 14058 30912
rect 14002 30424 14058 30433
rect 14002 30359 14004 30368
rect 14056 30359 14058 30368
rect 14004 30330 14056 30336
rect 13912 29640 13964 29646
rect 13912 29582 13964 29588
rect 13912 29504 13964 29510
rect 13912 29446 13964 29452
rect 13924 24954 13952 29446
rect 14108 28937 14136 31758
rect 14094 28928 14150 28937
rect 14094 28863 14150 28872
rect 14200 28257 14228 35391
rect 14646 34912 14702 34921
rect 14646 34847 14702 34856
rect 14660 34626 14688 34847
rect 14292 34598 14688 34626
rect 14292 34542 14320 34598
rect 14280 34536 14332 34542
rect 14280 34478 14332 34484
rect 14464 34536 14516 34542
rect 14464 34478 14516 34484
rect 14476 34134 14504 34478
rect 14372 34128 14424 34134
rect 14370 34096 14372 34105
rect 14464 34128 14516 34134
rect 14424 34096 14426 34105
rect 14464 34070 14516 34076
rect 14370 34031 14426 34040
rect 14476 33930 14504 34070
rect 14556 33992 14608 33998
rect 14556 33934 14608 33940
rect 14464 33924 14516 33930
rect 14464 33866 14516 33872
rect 14372 33516 14424 33522
rect 14372 33458 14424 33464
rect 14280 31272 14332 31278
rect 14280 31214 14332 31220
rect 14292 30394 14320 31214
rect 14280 30388 14332 30394
rect 14280 30330 14332 30336
rect 14280 30252 14332 30258
rect 14280 30194 14332 30200
rect 14292 30161 14320 30194
rect 14278 30152 14334 30161
rect 14278 30087 14334 30096
rect 14278 29744 14334 29753
rect 14278 29679 14334 29688
rect 14292 29073 14320 29679
rect 14384 29322 14412 33458
rect 14568 33386 14596 33934
rect 14556 33380 14608 33386
rect 14556 33322 14608 33328
rect 14660 32434 14688 34598
rect 14648 32428 14700 32434
rect 14648 32370 14700 32376
rect 14660 32314 14688 32370
rect 14476 32286 14688 32314
rect 14476 29510 14504 32286
rect 14646 32056 14702 32065
rect 14646 31991 14702 32000
rect 14660 31754 14688 31991
rect 14648 31748 14700 31754
rect 14648 31690 14700 31696
rect 14556 30864 14608 30870
rect 14556 30806 14608 30812
rect 14568 30190 14596 30806
rect 14556 30184 14608 30190
rect 14556 30126 14608 30132
rect 14648 30116 14700 30122
rect 14648 30058 14700 30064
rect 14660 29714 14688 30058
rect 14648 29708 14700 29714
rect 14648 29650 14700 29656
rect 14752 29560 14780 35974
rect 14844 32978 14872 36638
rect 15016 36576 15068 36582
rect 15016 36518 15068 36524
rect 14924 36032 14976 36038
rect 14924 35974 14976 35980
rect 14832 32972 14884 32978
rect 14832 32914 14884 32920
rect 14832 32768 14884 32774
rect 14832 32710 14884 32716
rect 14844 30054 14872 32710
rect 14936 31770 14964 35974
rect 15028 34678 15056 36518
rect 15212 35766 15240 37062
rect 15568 36916 15620 36922
rect 15568 36858 15620 36864
rect 15292 36712 15344 36718
rect 15292 36654 15344 36660
rect 15304 36174 15332 36654
rect 15292 36168 15344 36174
rect 15292 36110 15344 36116
rect 15384 36032 15436 36038
rect 15384 35974 15436 35980
rect 15200 35760 15252 35766
rect 15200 35702 15252 35708
rect 15292 35692 15344 35698
rect 15292 35634 15344 35640
rect 15108 35284 15160 35290
rect 15108 35226 15160 35232
rect 15200 35284 15252 35290
rect 15200 35226 15252 35232
rect 15016 34672 15068 34678
rect 15016 34614 15068 34620
rect 15120 34610 15148 35226
rect 15212 35193 15240 35226
rect 15198 35184 15254 35193
rect 15198 35119 15254 35128
rect 15304 35034 15332 35634
rect 15212 35006 15332 35034
rect 15108 34604 15160 34610
rect 15108 34546 15160 34552
rect 15108 33652 15160 33658
rect 15108 33594 15160 33600
rect 15120 33114 15148 33594
rect 15108 33108 15160 33114
rect 15108 33050 15160 33056
rect 15212 33017 15240 35006
rect 15292 34944 15344 34950
rect 15292 34886 15344 34892
rect 15198 33008 15254 33017
rect 15198 32943 15254 32952
rect 15212 32910 15240 32943
rect 15200 32904 15252 32910
rect 15200 32846 15252 32852
rect 15304 31958 15332 34886
rect 15396 33930 15424 35974
rect 15474 35728 15530 35737
rect 15474 35663 15476 35672
rect 15528 35663 15530 35672
rect 15476 35634 15528 35640
rect 15476 35488 15528 35494
rect 15476 35430 15528 35436
rect 15384 33924 15436 33930
rect 15384 33866 15436 33872
rect 15384 33312 15436 33318
rect 15384 33254 15436 33260
rect 15292 31952 15344 31958
rect 15292 31894 15344 31900
rect 15108 31816 15160 31822
rect 15106 31784 15108 31793
rect 15160 31784 15162 31793
rect 14936 31742 15056 31770
rect 14924 31680 14976 31686
rect 14922 31648 14924 31657
rect 14976 31648 14978 31657
rect 14922 31583 14978 31592
rect 14924 31408 14976 31414
rect 14924 31350 14976 31356
rect 14936 30258 14964 31350
rect 15028 31260 15056 31742
rect 15106 31719 15162 31728
rect 15292 31748 15344 31754
rect 15292 31690 15344 31696
rect 15028 31232 15148 31260
rect 14924 30252 14976 30258
rect 14924 30194 14976 30200
rect 14832 30048 14884 30054
rect 14832 29990 14884 29996
rect 14924 29572 14976 29578
rect 14752 29532 14924 29560
rect 14924 29514 14976 29520
rect 14464 29504 14516 29510
rect 14464 29446 14516 29452
rect 14384 29294 14688 29322
rect 14556 29232 14608 29238
rect 14556 29174 14608 29180
rect 14464 29096 14516 29102
rect 14278 29064 14334 29073
rect 14334 29022 14412 29050
rect 14464 29038 14516 29044
rect 14278 28999 14334 29008
rect 14384 28762 14412 29022
rect 14372 28756 14424 28762
rect 14372 28698 14424 28704
rect 14476 28642 14504 29038
rect 14292 28614 14504 28642
rect 14186 28248 14242 28257
rect 14186 28183 14242 28192
rect 14188 27464 14240 27470
rect 14188 27406 14240 27412
rect 14004 26512 14056 26518
rect 14004 26454 14056 26460
rect 13912 24948 13964 24954
rect 13912 24890 13964 24896
rect 13820 24812 13872 24818
rect 13820 24754 13872 24760
rect 13728 24404 13780 24410
rect 13728 24346 13780 24352
rect 13832 24274 13860 24754
rect 13912 24676 13964 24682
rect 13912 24618 13964 24624
rect 13820 24268 13872 24274
rect 13820 24210 13872 24216
rect 13820 23656 13872 23662
rect 13820 23598 13872 23604
rect 13832 23186 13860 23598
rect 13820 23180 13872 23186
rect 13820 23122 13872 23128
rect 13924 23050 13952 24618
rect 14016 23769 14044 26454
rect 14200 24614 14228 27406
rect 14292 26926 14320 28614
rect 14568 27606 14596 29174
rect 14556 27600 14608 27606
rect 14556 27542 14608 27548
rect 14372 27532 14424 27538
rect 14372 27474 14424 27480
rect 14280 26920 14332 26926
rect 14280 26862 14332 26868
rect 14384 25974 14412 27474
rect 14556 27056 14608 27062
rect 14556 26998 14608 27004
rect 14660 27010 14688 29294
rect 14832 28756 14884 28762
rect 14832 28698 14884 28704
rect 14844 27946 14872 28698
rect 14936 28150 14964 29514
rect 15120 28626 15148 31232
rect 15304 28966 15332 31690
rect 15396 30172 15424 33254
rect 15488 32502 15516 35430
rect 15580 35018 15608 36858
rect 15764 36786 15792 37062
rect 15752 36780 15804 36786
rect 15752 36722 15804 36728
rect 15752 36304 15804 36310
rect 15752 36246 15804 36252
rect 15764 36174 15792 36246
rect 15752 36168 15804 36174
rect 15752 36110 15804 36116
rect 15856 36009 15884 37198
rect 15934 36408 15990 36417
rect 15934 36343 15990 36352
rect 15948 36310 15976 36343
rect 15936 36304 15988 36310
rect 15936 36246 15988 36252
rect 16028 36168 16080 36174
rect 16028 36110 16080 36116
rect 15842 36000 15898 36009
rect 15842 35935 15898 35944
rect 16040 35698 16068 36110
rect 16396 36032 16448 36038
rect 16396 35974 16448 35980
rect 16028 35692 16080 35698
rect 16028 35634 16080 35640
rect 15660 35624 15712 35630
rect 15660 35566 15712 35572
rect 15568 35012 15620 35018
rect 15568 34954 15620 34960
rect 15672 34610 15700 35566
rect 15660 34604 15712 34610
rect 15660 34546 15712 34552
rect 15752 34536 15804 34542
rect 15752 34478 15804 34484
rect 15658 34096 15714 34105
rect 15658 34031 15714 34040
rect 15672 33998 15700 34031
rect 15660 33992 15712 33998
rect 15660 33934 15712 33940
rect 15568 33652 15620 33658
rect 15568 33594 15620 33600
rect 15476 32496 15528 32502
rect 15476 32438 15528 32444
rect 15476 32360 15528 32366
rect 15476 32302 15528 32308
rect 15488 32065 15516 32302
rect 15474 32056 15530 32065
rect 15474 31991 15530 32000
rect 15476 31884 15528 31890
rect 15476 31826 15528 31832
rect 15488 30666 15516 31826
rect 15580 31686 15608 33594
rect 15660 33448 15712 33454
rect 15660 33390 15712 33396
rect 15568 31680 15620 31686
rect 15568 31622 15620 31628
rect 15568 31340 15620 31346
rect 15568 31282 15620 31288
rect 15580 30870 15608 31282
rect 15672 30938 15700 33390
rect 15764 31226 15792 34478
rect 15936 33924 15988 33930
rect 15936 33866 15988 33872
rect 15948 33046 15976 33866
rect 15936 33040 15988 33046
rect 15936 32982 15988 32988
rect 15842 32056 15898 32065
rect 15842 31991 15898 32000
rect 15856 31346 15884 31991
rect 15844 31340 15896 31346
rect 15844 31282 15896 31288
rect 16040 31278 16068 35634
rect 16120 35624 16172 35630
rect 16120 35566 16172 35572
rect 16132 35494 16160 35566
rect 16120 35488 16172 35494
rect 16120 35430 16172 35436
rect 16120 35080 16172 35086
rect 16120 35022 16172 35028
rect 16212 35080 16264 35086
rect 16212 35022 16264 35028
rect 16132 34785 16160 35022
rect 16118 34776 16174 34785
rect 16118 34711 16174 34720
rect 16224 34202 16252 35022
rect 16212 34196 16264 34202
rect 16212 34138 16264 34144
rect 16408 33658 16436 35974
rect 16488 35488 16540 35494
rect 16488 35430 16540 35436
rect 16396 33652 16448 33658
rect 16396 33594 16448 33600
rect 16500 32978 16528 35430
rect 16580 34536 16632 34542
rect 16580 34478 16632 34484
rect 16212 32972 16264 32978
rect 16212 32914 16264 32920
rect 16488 32972 16540 32978
rect 16488 32914 16540 32920
rect 16120 31884 16172 31890
rect 16120 31826 16172 31832
rect 16028 31272 16080 31278
rect 15764 31198 15884 31226
rect 16028 31214 16080 31220
rect 15752 31136 15804 31142
rect 15752 31078 15804 31084
rect 15660 30932 15712 30938
rect 15660 30874 15712 30880
rect 15568 30864 15620 30870
rect 15568 30806 15620 30812
rect 15476 30660 15528 30666
rect 15476 30602 15528 30608
rect 15660 30592 15712 30598
rect 15660 30534 15712 30540
rect 15568 30184 15620 30190
rect 15396 30144 15568 30172
rect 15568 30126 15620 30132
rect 15476 29776 15528 29782
rect 15476 29718 15528 29724
rect 15292 28960 15344 28966
rect 15292 28902 15344 28908
rect 15384 28960 15436 28966
rect 15384 28902 15436 28908
rect 15108 28620 15160 28626
rect 15108 28562 15160 28568
rect 14924 28144 14976 28150
rect 14924 28086 14976 28092
rect 14832 27940 14884 27946
rect 14832 27882 14884 27888
rect 15120 27130 15148 28562
rect 15200 28484 15252 28490
rect 15200 28426 15252 28432
rect 15212 27878 15240 28426
rect 15200 27872 15252 27878
rect 15200 27814 15252 27820
rect 15304 27334 15332 28902
rect 15396 28014 15424 28902
rect 15384 28008 15436 28014
rect 15384 27950 15436 27956
rect 15396 27606 15424 27950
rect 15384 27600 15436 27606
rect 15384 27542 15436 27548
rect 15292 27328 15344 27334
rect 15292 27270 15344 27276
rect 15108 27124 15160 27130
rect 15108 27066 15160 27072
rect 14462 26752 14518 26761
rect 14462 26687 14518 26696
rect 14476 25974 14504 26687
rect 14372 25968 14424 25974
rect 14372 25910 14424 25916
rect 14464 25968 14516 25974
rect 14464 25910 14516 25916
rect 14370 25800 14426 25809
rect 14476 25770 14504 25910
rect 14370 25735 14426 25744
rect 14464 25764 14516 25770
rect 14280 25288 14332 25294
rect 14278 25256 14280 25265
rect 14332 25256 14334 25265
rect 14278 25191 14334 25200
rect 14384 24886 14412 25735
rect 14464 25706 14516 25712
rect 14464 25152 14516 25158
rect 14464 25094 14516 25100
rect 14372 24880 14424 24886
rect 14372 24822 14424 24828
rect 14372 24744 14424 24750
rect 14372 24686 14424 24692
rect 14188 24608 14240 24614
rect 14188 24550 14240 24556
rect 14280 24268 14332 24274
rect 14280 24210 14332 24216
rect 14002 23760 14058 23769
rect 14002 23695 14058 23704
rect 13912 23044 13964 23050
rect 13912 22986 13964 22992
rect 13636 22092 13688 22098
rect 13636 22034 13688 22040
rect 13648 21978 13676 22034
rect 13648 21950 13768 21978
rect 13740 21010 13768 21950
rect 14292 21486 14320 24210
rect 14384 23594 14412 24686
rect 14372 23588 14424 23594
rect 14372 23530 14424 23536
rect 14280 21480 14332 21486
rect 14280 21422 14332 21428
rect 14384 21010 14412 23530
rect 13728 21004 13780 21010
rect 13728 20946 13780 20952
rect 14372 21004 14424 21010
rect 14372 20946 14424 20952
rect 13544 20596 13596 20602
rect 13544 20538 13596 20544
rect 13728 20528 13780 20534
rect 13728 20470 13780 20476
rect 14280 20528 14332 20534
rect 14280 20470 14332 20476
rect 13740 20058 13768 20470
rect 14188 20392 14240 20398
rect 14188 20334 14240 20340
rect 13728 20052 13780 20058
rect 13728 19994 13780 20000
rect 13360 19984 13412 19990
rect 13360 19926 13412 19932
rect 13544 19780 13596 19786
rect 13544 19722 13596 19728
rect 13556 19514 13584 19722
rect 13636 19712 13688 19718
rect 13636 19654 13688 19660
rect 13544 19508 13596 19514
rect 13544 19450 13596 19456
rect 13648 19378 13676 19654
rect 13740 19446 13768 19994
rect 14200 19446 14228 20334
rect 13728 19440 13780 19446
rect 13728 19382 13780 19388
rect 14188 19440 14240 19446
rect 14188 19382 14240 19388
rect 13636 19372 13688 19378
rect 13636 19314 13688 19320
rect 13648 18902 13676 19314
rect 14200 18970 14228 19382
rect 14188 18964 14240 18970
rect 14188 18906 14240 18912
rect 13636 18896 13688 18902
rect 13636 18838 13688 18844
rect 13912 18828 13964 18834
rect 13912 18770 13964 18776
rect 13544 18760 13596 18766
rect 13544 18702 13596 18708
rect 13556 18358 13584 18702
rect 13728 18624 13780 18630
rect 13728 18566 13780 18572
rect 13544 18352 13596 18358
rect 13544 18294 13596 18300
rect 13740 18290 13768 18566
rect 13728 18284 13780 18290
rect 13728 18226 13780 18232
rect 13924 18222 13952 18770
rect 14292 18426 14320 20470
rect 14384 20398 14412 20946
rect 14372 20392 14424 20398
rect 14372 20334 14424 20340
rect 14280 18420 14332 18426
rect 14280 18362 14332 18368
rect 13912 18216 13964 18222
rect 13912 18158 13964 18164
rect 13924 17338 13952 18158
rect 13912 17332 13964 17338
rect 13912 17274 13964 17280
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13084 10804 13136 10810
rect 13084 10746 13136 10752
rect 12714 10296 12770 10305
rect 12714 10231 12716 10240
rect 12768 10231 12770 10240
rect 12716 10202 12768 10208
rect 12728 10062 12756 10202
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 13268 9920 13320 9926
rect 13268 9862 13320 9868
rect 12716 3052 12768 3058
rect 12716 2994 12768 3000
rect 11520 2916 11572 2922
rect 11520 2858 11572 2864
rect 11886 2680 11942 2689
rect 11886 2615 11888 2624
rect 11940 2615 11942 2624
rect 11888 2586 11940 2592
rect 8576 2508 8628 2514
rect 8576 2450 8628 2456
rect 12728 2446 12756 2994
rect 13280 2446 13308 9862
rect 13464 3058 13492 13262
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13832 9722 13860 10406
rect 13820 9716 13872 9722
rect 13820 9658 13872 9664
rect 13452 3052 13504 3058
rect 13452 2994 13504 3000
rect 14476 2650 14504 25094
rect 14568 23254 14596 26998
rect 14660 26982 15148 27010
rect 14740 26784 14792 26790
rect 14740 26726 14792 26732
rect 14752 26382 14780 26726
rect 14740 26376 14792 26382
rect 14740 26318 14792 26324
rect 14832 26308 14884 26314
rect 14832 26250 14884 26256
rect 14648 25900 14700 25906
rect 14844 25888 14872 26250
rect 14700 25860 14872 25888
rect 14648 25842 14700 25848
rect 14740 25764 14792 25770
rect 14740 25706 14792 25712
rect 14648 25696 14700 25702
rect 14648 25638 14700 25644
rect 14556 23248 14608 23254
rect 14556 23190 14608 23196
rect 14556 22976 14608 22982
rect 14556 22918 14608 22924
rect 14568 22506 14596 22918
rect 14556 22500 14608 22506
rect 14556 22442 14608 22448
rect 14660 22094 14688 25638
rect 14752 25498 14780 25706
rect 14740 25492 14792 25498
rect 14740 25434 14792 25440
rect 15016 25492 15068 25498
rect 15016 25434 15068 25440
rect 15028 25226 15056 25434
rect 15016 25220 15068 25226
rect 15016 25162 15068 25168
rect 14924 24336 14976 24342
rect 14924 24278 14976 24284
rect 14740 24132 14792 24138
rect 14740 24074 14792 24080
rect 14832 24132 14884 24138
rect 14832 24074 14884 24080
rect 14752 23322 14780 24074
rect 14844 23866 14872 24074
rect 14832 23860 14884 23866
rect 14832 23802 14884 23808
rect 14740 23316 14792 23322
rect 14740 23258 14792 23264
rect 14936 22710 14964 24278
rect 15016 23656 15068 23662
rect 15016 23598 15068 23604
rect 15028 23050 15056 23598
rect 15016 23044 15068 23050
rect 15016 22986 15068 22992
rect 14924 22704 14976 22710
rect 14924 22646 14976 22652
rect 14568 22066 14688 22094
rect 14568 22030 14596 22066
rect 14556 22024 14608 22030
rect 14556 21966 14608 21972
rect 14568 19922 14596 21966
rect 14936 20330 14964 22646
rect 15028 21486 15056 22986
rect 15016 21480 15068 21486
rect 15016 21422 15068 21428
rect 14924 20324 14976 20330
rect 14924 20266 14976 20272
rect 14832 20256 14884 20262
rect 14832 20198 14884 20204
rect 14556 19916 14608 19922
rect 14556 19858 14608 19864
rect 14844 19786 14872 20198
rect 14832 19780 14884 19786
rect 14832 19722 14884 19728
rect 14648 19168 14700 19174
rect 14648 19110 14700 19116
rect 14660 18766 14688 19110
rect 14648 18760 14700 18766
rect 14648 18702 14700 18708
rect 14844 17746 14872 19722
rect 15028 19310 15056 21422
rect 15016 19304 15068 19310
rect 15016 19246 15068 19252
rect 15120 19122 15148 26982
rect 15304 26790 15332 27270
rect 15292 26784 15344 26790
rect 15292 26726 15344 26732
rect 15384 26512 15436 26518
rect 15384 26454 15436 26460
rect 15396 26314 15424 26454
rect 15384 26308 15436 26314
rect 15384 26250 15436 26256
rect 15292 25968 15344 25974
rect 15292 25910 15344 25916
rect 15304 23322 15332 25910
rect 15384 25696 15436 25702
rect 15384 25638 15436 25644
rect 15396 25226 15424 25638
rect 15384 25220 15436 25226
rect 15384 25162 15436 25168
rect 15488 23798 15516 29718
rect 15580 28422 15608 30126
rect 15672 29753 15700 30534
rect 15658 29744 15714 29753
rect 15658 29679 15714 29688
rect 15568 28416 15620 28422
rect 15568 28358 15620 28364
rect 15672 27946 15700 29679
rect 15764 29238 15792 31078
rect 15856 30326 15884 31198
rect 16028 30932 16080 30938
rect 16028 30874 16080 30880
rect 15936 30388 15988 30394
rect 15936 30330 15988 30336
rect 15844 30320 15896 30326
rect 15844 30262 15896 30268
rect 15948 29578 15976 30330
rect 15936 29572 15988 29578
rect 15936 29514 15988 29520
rect 15752 29232 15804 29238
rect 15752 29174 15804 29180
rect 15936 29232 15988 29238
rect 15936 29174 15988 29180
rect 15752 28620 15804 28626
rect 15752 28562 15804 28568
rect 15660 27940 15712 27946
rect 15660 27882 15712 27888
rect 15568 27396 15620 27402
rect 15568 27338 15620 27344
rect 15580 24750 15608 27338
rect 15764 26518 15792 28562
rect 15844 26852 15896 26858
rect 15844 26794 15896 26800
rect 15752 26512 15804 26518
rect 15752 26454 15804 26460
rect 15752 25968 15804 25974
rect 15752 25910 15804 25916
rect 15658 24848 15714 24857
rect 15658 24783 15660 24792
rect 15712 24783 15714 24792
rect 15660 24754 15712 24760
rect 15568 24744 15620 24750
rect 15568 24686 15620 24692
rect 15568 24608 15620 24614
rect 15568 24550 15620 24556
rect 15476 23792 15528 23798
rect 15476 23734 15528 23740
rect 15292 23316 15344 23322
rect 15292 23258 15344 23264
rect 15580 23118 15608 24550
rect 15568 23112 15620 23118
rect 15568 23054 15620 23060
rect 15200 22772 15252 22778
rect 15200 22714 15252 22720
rect 15028 19094 15148 19122
rect 14832 17740 14884 17746
rect 14832 17682 14884 17688
rect 14556 17604 14608 17610
rect 14556 17546 14608 17552
rect 14568 17338 14596 17546
rect 14556 17332 14608 17338
rect 14556 17274 14608 17280
rect 15028 17202 15056 19094
rect 15212 18970 15240 22714
rect 15384 22568 15436 22574
rect 15384 22510 15436 22516
rect 15292 22432 15344 22438
rect 15292 22374 15344 22380
rect 15304 19786 15332 22374
rect 15396 22030 15424 22510
rect 15580 22234 15608 23054
rect 15568 22228 15620 22234
rect 15568 22170 15620 22176
rect 15384 22024 15436 22030
rect 15672 22001 15700 24754
rect 15764 24614 15792 25910
rect 15752 24608 15804 24614
rect 15752 24550 15804 24556
rect 15856 24410 15884 26794
rect 15948 24954 15976 29174
rect 16040 25770 16068 30874
rect 16132 29050 16160 31826
rect 16224 29782 16252 32914
rect 16304 32292 16356 32298
rect 16304 32234 16356 32240
rect 16316 31958 16344 32234
rect 16304 31952 16356 31958
rect 16304 31894 16356 31900
rect 16396 31952 16448 31958
rect 16396 31894 16448 31900
rect 16304 31340 16356 31346
rect 16304 31282 16356 31288
rect 16212 29776 16264 29782
rect 16212 29718 16264 29724
rect 16316 29238 16344 31282
rect 16408 29889 16436 31894
rect 16592 31482 16620 34478
rect 16684 33289 16712 37742
rect 16776 37262 16804 39200
rect 16856 37324 16908 37330
rect 16856 37266 16908 37272
rect 18604 37324 18656 37330
rect 18604 37266 18656 37272
rect 16764 37256 16816 37262
rect 16764 37198 16816 37204
rect 16868 36666 16896 37266
rect 18512 37120 18564 37126
rect 18616 37097 18644 37266
rect 18708 37108 18736 39200
rect 20536 37460 20588 37466
rect 20536 37402 20588 37408
rect 19432 37256 19484 37262
rect 19432 37198 19484 37204
rect 18788 37120 18840 37126
rect 18512 37062 18564 37068
rect 18602 37088 18658 37097
rect 17868 36848 17920 36854
rect 17868 36790 17920 36796
rect 18524 36802 18552 37062
rect 18708 37080 18788 37108
rect 18788 37062 18840 37068
rect 18602 37023 18658 37032
rect 17500 36780 17552 36786
rect 17500 36722 17552 36728
rect 16776 36638 16896 36666
rect 16670 33280 16726 33289
rect 16670 33215 16726 33224
rect 16684 32366 16712 33215
rect 16672 32360 16724 32366
rect 16672 32302 16724 32308
rect 16672 31816 16724 31822
rect 16672 31758 16724 31764
rect 16580 31476 16632 31482
rect 16580 31418 16632 31424
rect 16684 31385 16712 31758
rect 16670 31376 16726 31385
rect 16670 31311 16726 31320
rect 16672 30728 16724 30734
rect 16670 30696 16672 30705
rect 16724 30696 16726 30705
rect 16670 30631 16726 30640
rect 16580 30592 16632 30598
rect 16776 30546 16804 36638
rect 16856 36576 16908 36582
rect 16856 36518 16908 36524
rect 16868 36106 16896 36518
rect 16856 36100 16908 36106
rect 16856 36042 16908 36048
rect 16948 35760 17000 35766
rect 16946 35728 16948 35737
rect 17000 35728 17002 35737
rect 16946 35663 17002 35672
rect 16948 35488 17000 35494
rect 16948 35430 17000 35436
rect 16856 34944 16908 34950
rect 16856 34886 16908 34892
rect 16868 31482 16896 34886
rect 16960 33590 16988 35430
rect 17316 35012 17368 35018
rect 17316 34954 17368 34960
rect 17040 34944 17092 34950
rect 17038 34912 17040 34921
rect 17092 34912 17094 34921
rect 17038 34847 17094 34856
rect 17132 34536 17184 34542
rect 17132 34478 17184 34484
rect 17040 34060 17092 34066
rect 17040 34002 17092 34008
rect 16948 33584 17000 33590
rect 16948 33526 17000 33532
rect 17052 32910 17080 34002
rect 17040 32904 17092 32910
rect 17040 32846 17092 32852
rect 17144 32842 17172 34478
rect 17224 34196 17276 34202
rect 17224 34138 17276 34144
rect 17236 33454 17264 34138
rect 17328 33998 17356 34954
rect 17316 33992 17368 33998
rect 17316 33934 17368 33940
rect 17328 33522 17356 33934
rect 17406 33688 17462 33697
rect 17406 33623 17408 33632
rect 17460 33623 17462 33632
rect 17408 33594 17460 33600
rect 17316 33516 17368 33522
rect 17316 33458 17368 33464
rect 17224 33448 17276 33454
rect 17224 33390 17276 33396
rect 17236 32910 17264 33390
rect 17316 32972 17368 32978
rect 17316 32914 17368 32920
rect 17224 32904 17276 32910
rect 17224 32846 17276 32852
rect 17132 32836 17184 32842
rect 17132 32778 17184 32784
rect 16948 32224 17000 32230
rect 16948 32166 17000 32172
rect 16960 32026 16988 32166
rect 16948 32020 17000 32026
rect 16948 31962 17000 31968
rect 17236 31822 17264 32846
rect 17328 32842 17356 32914
rect 17316 32836 17368 32842
rect 17316 32778 17368 32784
rect 17328 32745 17356 32778
rect 17512 32774 17540 36722
rect 17776 36032 17828 36038
rect 17776 35974 17828 35980
rect 17788 35698 17816 35974
rect 17776 35692 17828 35698
rect 17776 35634 17828 35640
rect 17788 35494 17816 35634
rect 17776 35488 17828 35494
rect 17776 35430 17828 35436
rect 17880 35018 17908 36790
rect 18052 36780 18104 36786
rect 18524 36774 19012 36802
rect 18052 36722 18104 36728
rect 17958 35864 18014 35873
rect 17958 35799 17960 35808
rect 18012 35799 18014 35808
rect 17960 35770 18012 35776
rect 17958 35320 18014 35329
rect 18064 35290 18092 36722
rect 18788 36576 18840 36582
rect 18788 36518 18840 36524
rect 18694 36136 18750 36145
rect 18694 36071 18750 36080
rect 18512 36032 18564 36038
rect 18512 35974 18564 35980
rect 18420 35692 18472 35698
rect 18420 35634 18472 35640
rect 17958 35255 18014 35264
rect 18052 35284 18104 35290
rect 17972 35018 18000 35255
rect 18052 35226 18104 35232
rect 17868 35012 17920 35018
rect 17868 34954 17920 34960
rect 17960 35012 18012 35018
rect 17960 34954 18012 34960
rect 18064 34678 18092 35226
rect 18236 34740 18288 34746
rect 18236 34682 18288 34688
rect 17592 34672 17644 34678
rect 18052 34672 18104 34678
rect 17592 34614 17644 34620
rect 17958 34640 18014 34649
rect 17500 32768 17552 32774
rect 17314 32736 17370 32745
rect 17500 32710 17552 32716
rect 17314 32671 17370 32680
rect 17408 32428 17460 32434
rect 17512 32416 17540 32710
rect 17460 32388 17540 32416
rect 17408 32370 17460 32376
rect 17406 32328 17462 32337
rect 17406 32263 17462 32272
rect 17420 32230 17448 32263
rect 17316 32224 17368 32230
rect 17316 32166 17368 32172
rect 17408 32224 17460 32230
rect 17408 32166 17460 32172
rect 17224 31816 17276 31822
rect 17224 31758 17276 31764
rect 16946 31648 17002 31657
rect 16946 31583 17002 31592
rect 16960 31482 16988 31583
rect 16856 31476 16908 31482
rect 16856 31418 16908 31424
rect 16948 31476 17000 31482
rect 16948 31418 17000 31424
rect 17328 30666 17356 32166
rect 17604 31754 17632 34614
rect 18052 34614 18104 34620
rect 17958 34575 17960 34584
rect 18012 34575 18014 34584
rect 17960 34546 18012 34552
rect 18064 33998 18092 34614
rect 18248 34610 18276 34682
rect 18236 34604 18288 34610
rect 18236 34546 18288 34552
rect 17960 33992 18012 33998
rect 17960 33934 18012 33940
rect 18052 33992 18104 33998
rect 18052 33934 18104 33940
rect 17684 33040 17736 33046
rect 17684 32982 17736 32988
rect 17696 31890 17724 32982
rect 17972 32722 18000 33934
rect 18064 32842 18092 33934
rect 18432 33590 18460 35634
rect 18524 35465 18552 35974
rect 18510 35456 18566 35465
rect 18510 35391 18566 35400
rect 18708 35290 18736 36071
rect 18696 35284 18748 35290
rect 18696 35226 18748 35232
rect 18696 35080 18748 35086
rect 18800 35057 18828 36518
rect 18880 36168 18932 36174
rect 18880 36110 18932 36116
rect 18696 35022 18748 35028
rect 18786 35048 18842 35057
rect 18604 34060 18656 34066
rect 18604 34002 18656 34008
rect 18420 33584 18472 33590
rect 18420 33526 18472 33532
rect 18510 33552 18566 33561
rect 18144 33040 18196 33046
rect 18144 32982 18196 32988
rect 18156 32910 18184 32982
rect 18144 32904 18196 32910
rect 18144 32846 18196 32852
rect 18236 32904 18288 32910
rect 18236 32846 18288 32852
rect 18052 32836 18104 32842
rect 18052 32778 18104 32784
rect 18248 32722 18276 32846
rect 17972 32694 18276 32722
rect 17684 31884 17736 31890
rect 17684 31826 17736 31832
rect 17592 31748 17644 31754
rect 17592 31690 17644 31696
rect 17406 30968 17462 30977
rect 17406 30903 17462 30912
rect 17040 30660 17092 30666
rect 17040 30602 17092 30608
rect 17316 30660 17368 30666
rect 17316 30602 17368 30608
rect 16580 30534 16632 30540
rect 16394 29880 16450 29889
rect 16394 29815 16450 29824
rect 16396 29572 16448 29578
rect 16396 29514 16448 29520
rect 16304 29232 16356 29238
rect 16304 29174 16356 29180
rect 16408 29186 16436 29514
rect 16592 29510 16620 30534
rect 16684 30518 16804 30546
rect 17052 30546 17080 30602
rect 17052 30518 17264 30546
rect 16684 30258 16712 30518
rect 16856 30388 16908 30394
rect 16856 30330 16908 30336
rect 16672 30252 16724 30258
rect 16672 30194 16724 30200
rect 16684 29782 16712 30194
rect 16764 30184 16816 30190
rect 16764 30126 16816 30132
rect 16672 29776 16724 29782
rect 16672 29718 16724 29724
rect 16580 29504 16632 29510
rect 16580 29446 16632 29452
rect 16672 29504 16724 29510
rect 16672 29446 16724 29452
rect 16408 29158 16528 29186
rect 16684 29170 16712 29446
rect 16132 29034 16252 29050
rect 16132 29028 16264 29034
rect 16132 29022 16212 29028
rect 16212 28970 16264 28976
rect 16120 28688 16172 28694
rect 16120 28630 16172 28636
rect 16132 28218 16160 28630
rect 16120 28212 16172 28218
rect 16120 28154 16172 28160
rect 16118 28112 16174 28121
rect 16118 28047 16174 28056
rect 16132 27470 16160 28047
rect 16120 27464 16172 27470
rect 16120 27406 16172 27412
rect 16132 26926 16160 27406
rect 16224 27010 16252 28970
rect 16396 28484 16448 28490
rect 16396 28426 16448 28432
rect 16408 27606 16436 28426
rect 16500 27946 16528 29158
rect 16672 29164 16724 29170
rect 16672 29106 16724 29112
rect 16580 29096 16632 29102
rect 16580 29038 16632 29044
rect 16592 28626 16620 29038
rect 16684 28801 16712 29106
rect 16670 28792 16726 28801
rect 16670 28727 16726 28736
rect 16580 28620 16632 28626
rect 16580 28562 16632 28568
rect 16488 27940 16540 27946
rect 16488 27882 16540 27888
rect 16396 27600 16448 27606
rect 16396 27542 16448 27548
rect 16396 27396 16448 27402
rect 16396 27338 16448 27344
rect 16224 26982 16344 27010
rect 16408 26994 16436 27338
rect 16120 26920 16172 26926
rect 16120 26862 16172 26868
rect 16210 26480 16266 26489
rect 16210 26415 16266 26424
rect 16224 25906 16252 26415
rect 16316 26382 16344 26982
rect 16396 26988 16448 26994
rect 16396 26930 16448 26936
rect 16500 26874 16528 27882
rect 16408 26846 16528 26874
rect 16304 26376 16356 26382
rect 16304 26318 16356 26324
rect 16212 25900 16264 25906
rect 16212 25842 16264 25848
rect 16028 25764 16080 25770
rect 16028 25706 16080 25712
rect 16316 25362 16344 26318
rect 16304 25356 16356 25362
rect 16304 25298 16356 25304
rect 16408 25242 16436 26846
rect 16488 26444 16540 26450
rect 16488 26386 16540 26392
rect 16500 25362 16528 26386
rect 16776 25362 16804 30126
rect 16868 28626 16896 30330
rect 17132 30048 17184 30054
rect 17132 29990 17184 29996
rect 17144 29578 17172 29990
rect 17040 29572 17092 29578
rect 17040 29514 17092 29520
rect 17132 29572 17184 29578
rect 17132 29514 17184 29520
rect 16948 29028 17000 29034
rect 16948 28970 17000 28976
rect 16856 28620 16908 28626
rect 16856 28562 16908 28568
rect 16854 27840 16910 27849
rect 16854 27775 16910 27784
rect 16868 27674 16896 27775
rect 16856 27668 16908 27674
rect 16856 27610 16908 27616
rect 16960 27062 16988 28970
rect 16948 27056 17000 27062
rect 16948 26998 17000 27004
rect 16946 26072 17002 26081
rect 16946 26007 17002 26016
rect 16856 25900 16908 25906
rect 16856 25842 16908 25848
rect 16488 25356 16540 25362
rect 16488 25298 16540 25304
rect 16764 25356 16816 25362
rect 16764 25298 16816 25304
rect 16316 25214 16436 25242
rect 16672 25220 16724 25226
rect 15936 24948 15988 24954
rect 15936 24890 15988 24896
rect 16316 24682 16344 25214
rect 16500 25180 16672 25208
rect 16500 24954 16528 25180
rect 16672 25162 16724 25168
rect 16488 24948 16540 24954
rect 16488 24890 16540 24896
rect 16396 24812 16448 24818
rect 16396 24754 16448 24760
rect 16304 24676 16356 24682
rect 16304 24618 16356 24624
rect 16212 24608 16264 24614
rect 16212 24550 16264 24556
rect 15844 24404 15896 24410
rect 15844 24346 15896 24352
rect 15856 24138 15884 24346
rect 15844 24132 15896 24138
rect 15844 24074 15896 24080
rect 15752 23520 15804 23526
rect 15752 23462 15804 23468
rect 15384 21966 15436 21972
rect 15658 21992 15714 22001
rect 15658 21927 15714 21936
rect 15384 21888 15436 21894
rect 15384 21830 15436 21836
rect 15396 20602 15424 21830
rect 15476 21616 15528 21622
rect 15476 21558 15528 21564
rect 15488 20602 15516 21558
rect 15660 21480 15712 21486
rect 15660 21422 15712 21428
rect 15568 21140 15620 21146
rect 15568 21082 15620 21088
rect 15384 20596 15436 20602
rect 15384 20538 15436 20544
rect 15476 20596 15528 20602
rect 15476 20538 15528 20544
rect 15292 19780 15344 19786
rect 15292 19722 15344 19728
rect 15292 19236 15344 19242
rect 15292 19178 15344 19184
rect 15200 18964 15252 18970
rect 15200 18906 15252 18912
rect 15108 18828 15160 18834
rect 15108 18770 15160 18776
rect 15120 18426 15148 18770
rect 15200 18760 15252 18766
rect 15200 18702 15252 18708
rect 15108 18420 15160 18426
rect 15108 18362 15160 18368
rect 15212 17882 15240 18702
rect 15304 18358 15332 19178
rect 15292 18352 15344 18358
rect 15292 18294 15344 18300
rect 15200 17876 15252 17882
rect 15200 17818 15252 17824
rect 15016 17196 15068 17202
rect 15016 17138 15068 17144
rect 14464 2644 14516 2650
rect 14464 2586 14516 2592
rect 15212 2582 15240 17818
rect 15304 17338 15332 18294
rect 15292 17332 15344 17338
rect 15292 17274 15344 17280
rect 15580 12238 15608 21082
rect 15672 21010 15700 21422
rect 15660 21004 15712 21010
rect 15660 20946 15712 20952
rect 15764 19854 15792 23462
rect 16028 23180 16080 23186
rect 16028 23122 16080 23128
rect 16040 22642 16068 23122
rect 16120 23044 16172 23050
rect 16120 22986 16172 22992
rect 16028 22636 16080 22642
rect 16028 22578 16080 22584
rect 16040 22094 16068 22578
rect 15856 22066 16068 22094
rect 15856 20466 15884 22066
rect 15936 21956 15988 21962
rect 15936 21898 15988 21904
rect 15948 21350 15976 21898
rect 16028 21888 16080 21894
rect 16028 21830 16080 21836
rect 16040 21486 16068 21830
rect 16028 21480 16080 21486
rect 16028 21422 16080 21428
rect 15936 21344 15988 21350
rect 15936 21286 15988 21292
rect 15948 21146 15976 21286
rect 15936 21140 15988 21146
rect 15936 21082 15988 21088
rect 16132 20534 16160 22986
rect 16224 22030 16252 24550
rect 16408 24410 16436 24754
rect 16396 24404 16448 24410
rect 16396 24346 16448 24352
rect 16776 24342 16804 25298
rect 16764 24336 16816 24342
rect 16764 24278 16816 24284
rect 16396 24268 16448 24274
rect 16396 24210 16448 24216
rect 16408 23798 16436 24210
rect 16580 24064 16632 24070
rect 16500 24012 16580 24018
rect 16500 24006 16632 24012
rect 16500 23990 16620 24006
rect 16396 23792 16448 23798
rect 16396 23734 16448 23740
rect 16500 23662 16528 23990
rect 16488 23656 16540 23662
rect 16488 23598 16540 23604
rect 16304 22704 16356 22710
rect 16304 22646 16356 22652
rect 16212 22024 16264 22030
rect 16212 21966 16264 21972
rect 16212 20800 16264 20806
rect 16212 20742 16264 20748
rect 16120 20528 16172 20534
rect 16120 20470 16172 20476
rect 15844 20460 15896 20466
rect 15844 20402 15896 20408
rect 15752 19848 15804 19854
rect 15752 19790 15804 19796
rect 15764 19378 15792 19790
rect 15752 19372 15804 19378
rect 15752 19314 15804 19320
rect 16224 18970 16252 20742
rect 16316 20058 16344 22646
rect 16394 21992 16450 22001
rect 16394 21927 16450 21936
rect 16304 20052 16356 20058
rect 16304 19994 16356 20000
rect 16304 19712 16356 19718
rect 16304 19654 16356 19660
rect 16316 19514 16344 19654
rect 16304 19508 16356 19514
rect 16304 19450 16356 19456
rect 16212 18964 16264 18970
rect 16212 18906 16264 18912
rect 16408 16574 16436 21927
rect 16500 19922 16528 23598
rect 16868 23322 16896 25842
rect 16856 23316 16908 23322
rect 16856 23258 16908 23264
rect 16764 23112 16816 23118
rect 16868 23100 16896 23258
rect 16816 23072 16896 23100
rect 16764 23054 16816 23060
rect 16856 22568 16908 22574
rect 16856 22510 16908 22516
rect 16868 20942 16896 22510
rect 16856 20936 16908 20942
rect 16856 20878 16908 20884
rect 16868 19922 16896 20878
rect 16960 20874 16988 26007
rect 17052 23594 17080 29514
rect 17130 28928 17186 28937
rect 17130 28863 17186 28872
rect 17144 25906 17172 28863
rect 17236 28762 17264 30518
rect 17314 30424 17370 30433
rect 17314 30359 17370 30368
rect 17224 28756 17276 28762
rect 17224 28698 17276 28704
rect 17328 26466 17356 30359
rect 17420 28937 17448 30903
rect 17406 28928 17462 28937
rect 17406 28863 17462 28872
rect 17696 28762 17724 31826
rect 17972 31793 18000 32694
rect 18432 32502 18460 33526
rect 18510 33487 18566 33496
rect 18524 33114 18552 33487
rect 18616 33454 18644 34002
rect 18708 33590 18736 35022
rect 18786 34983 18842 34992
rect 18696 33584 18748 33590
rect 18696 33526 18748 33532
rect 18604 33448 18656 33454
rect 18604 33390 18656 33396
rect 18512 33108 18564 33114
rect 18512 33050 18564 33056
rect 18420 32496 18472 32502
rect 18142 32464 18198 32473
rect 18420 32438 18472 32444
rect 18142 32399 18198 32408
rect 17958 31784 18014 31793
rect 17868 31748 17920 31754
rect 17958 31719 18014 31728
rect 17868 31690 17920 31696
rect 17880 31278 17908 31690
rect 17972 31346 18000 31719
rect 17960 31340 18012 31346
rect 17960 31282 18012 31288
rect 17868 31272 17920 31278
rect 17868 31214 17920 31220
rect 17776 31204 17828 31210
rect 17776 31146 17828 31152
rect 17788 30326 17816 31146
rect 17776 30320 17828 30326
rect 17776 30262 17828 30268
rect 17880 30190 17908 31214
rect 17868 30184 17920 30190
rect 17868 30126 17920 30132
rect 18052 30184 18104 30190
rect 18052 30126 18104 30132
rect 18064 29753 18092 30126
rect 18050 29744 18106 29753
rect 18050 29679 18052 29688
rect 18104 29679 18106 29688
rect 18052 29650 18104 29656
rect 17776 29572 17828 29578
rect 17776 29514 17828 29520
rect 17788 29034 17816 29514
rect 17776 29028 17828 29034
rect 17776 28970 17828 28976
rect 17684 28756 17736 28762
rect 17684 28698 17736 28704
rect 17776 28688 17828 28694
rect 17960 28688 18012 28694
rect 17828 28636 17960 28642
rect 17776 28630 18012 28636
rect 17788 28614 18000 28630
rect 17684 28484 17736 28490
rect 17684 28426 17736 28432
rect 17408 28144 17460 28150
rect 17408 28086 17460 28092
rect 17420 26586 17448 28086
rect 17592 27872 17644 27878
rect 17592 27814 17644 27820
rect 17604 27538 17632 27814
rect 17592 27532 17644 27538
rect 17592 27474 17644 27480
rect 17500 27396 17552 27402
rect 17500 27338 17552 27344
rect 17408 26580 17460 26586
rect 17408 26522 17460 26528
rect 17328 26438 17448 26466
rect 17316 26308 17368 26314
rect 17316 26250 17368 26256
rect 17328 26042 17356 26250
rect 17316 26036 17368 26042
rect 17316 25978 17368 25984
rect 17132 25900 17184 25906
rect 17132 25842 17184 25848
rect 17420 25702 17448 26438
rect 17512 26042 17540 27338
rect 17604 26926 17632 27474
rect 17592 26920 17644 26926
rect 17592 26862 17644 26868
rect 17604 26450 17632 26862
rect 17696 26489 17724 28426
rect 17868 27056 17920 27062
rect 17868 26998 17920 27004
rect 17682 26480 17738 26489
rect 17592 26444 17644 26450
rect 17682 26415 17738 26424
rect 17592 26386 17644 26392
rect 17500 26036 17552 26042
rect 17500 25978 17552 25984
rect 17408 25696 17460 25702
rect 17408 25638 17460 25644
rect 17592 24812 17644 24818
rect 17592 24754 17644 24760
rect 17316 24744 17368 24750
rect 17316 24686 17368 24692
rect 17224 24676 17276 24682
rect 17224 24618 17276 24624
rect 17040 23588 17092 23594
rect 17040 23530 17092 23536
rect 17132 23520 17184 23526
rect 17132 23462 17184 23468
rect 17144 22030 17172 23462
rect 17236 23186 17264 24618
rect 17328 23798 17356 24686
rect 17604 24614 17632 24754
rect 17682 24712 17738 24721
rect 17682 24647 17738 24656
rect 17592 24608 17644 24614
rect 17590 24576 17592 24585
rect 17644 24576 17646 24585
rect 17590 24511 17646 24520
rect 17316 23792 17368 23798
rect 17316 23734 17368 23740
rect 17500 23588 17552 23594
rect 17500 23530 17552 23536
rect 17224 23180 17276 23186
rect 17224 23122 17276 23128
rect 17132 22024 17184 22030
rect 17132 21966 17184 21972
rect 17040 21888 17092 21894
rect 17040 21830 17092 21836
rect 17052 21690 17080 21830
rect 17040 21684 17092 21690
rect 17040 21626 17092 21632
rect 16948 20868 17000 20874
rect 16948 20810 17000 20816
rect 17144 20602 17172 21966
rect 17224 21956 17276 21962
rect 17224 21898 17276 21904
rect 17132 20596 17184 20602
rect 17132 20538 17184 20544
rect 16488 19916 16540 19922
rect 16488 19858 16540 19864
rect 16856 19916 16908 19922
rect 16856 19858 16908 19864
rect 16500 18970 16528 19858
rect 17236 19378 17264 21898
rect 17512 21078 17540 23530
rect 17604 22642 17632 24511
rect 17696 23050 17724 24647
rect 17776 23316 17828 23322
rect 17776 23258 17828 23264
rect 17788 23118 17816 23258
rect 17880 23254 17908 26998
rect 17958 26072 18014 26081
rect 17958 26007 18014 26016
rect 17972 25906 18000 26007
rect 18156 25906 18184 32399
rect 18236 31476 18288 31482
rect 18236 31418 18288 31424
rect 18248 26586 18276 31418
rect 18432 31210 18460 32438
rect 18892 31754 18920 36110
rect 18984 34490 19012 36774
rect 19340 36576 19392 36582
rect 19340 36518 19392 36524
rect 19076 36366 19288 36394
rect 19076 36038 19104 36366
rect 19260 36310 19288 36366
rect 19156 36304 19208 36310
rect 19156 36246 19208 36252
rect 19248 36304 19300 36310
rect 19248 36246 19300 36252
rect 19064 36032 19116 36038
rect 19064 35974 19116 35980
rect 19168 34746 19196 36246
rect 19352 36106 19380 36518
rect 19340 36100 19392 36106
rect 19340 36042 19392 36048
rect 19352 35578 19380 36042
rect 19444 35714 19472 37198
rect 19984 37188 20036 37194
rect 19984 37130 20036 37136
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19996 36786 20024 37130
rect 19984 36780 20036 36786
rect 19984 36722 20036 36728
rect 20548 36582 20576 37402
rect 20640 37346 20668 39200
rect 20640 37318 20760 37346
rect 20732 37262 20760 37318
rect 20720 37256 20772 37262
rect 20720 37198 20772 37204
rect 21456 37256 21508 37262
rect 21456 37198 21508 37204
rect 20720 37120 20772 37126
rect 20720 37062 20772 37068
rect 20732 36718 20760 37062
rect 21468 36922 21496 37198
rect 21928 37108 21956 39200
rect 22744 37732 22796 37738
rect 22744 37674 22796 37680
rect 22756 37466 22784 37674
rect 23860 37466 23888 39200
rect 22744 37460 22796 37466
rect 22744 37402 22796 37408
rect 23848 37460 23900 37466
rect 23848 37402 23900 37408
rect 22100 37120 22152 37126
rect 21928 37080 22100 37108
rect 22100 37062 22152 37068
rect 21456 36916 21508 36922
rect 21456 36858 21508 36864
rect 20720 36712 20772 36718
rect 20720 36654 20772 36660
rect 20812 36712 20864 36718
rect 20812 36654 20864 36660
rect 19984 36576 20036 36582
rect 19984 36518 20036 36524
rect 20536 36576 20588 36582
rect 20536 36518 20588 36524
rect 19996 36242 20024 36518
rect 19984 36236 20036 36242
rect 19984 36178 20036 36184
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19996 35834 20024 36178
rect 19984 35828 20036 35834
rect 19984 35770 20036 35776
rect 19444 35686 19564 35714
rect 19536 35630 19564 35686
rect 19524 35624 19576 35630
rect 19352 35550 19472 35578
rect 19524 35566 19576 35572
rect 19248 35488 19300 35494
rect 19248 35430 19300 35436
rect 19260 35086 19288 35430
rect 19248 35080 19300 35086
rect 19248 35022 19300 35028
rect 19156 34740 19208 34746
rect 19156 34682 19208 34688
rect 19260 34610 19288 35022
rect 19248 34604 19300 34610
rect 19248 34546 19300 34552
rect 18984 34462 19196 34490
rect 19168 34406 19196 34462
rect 19064 34400 19116 34406
rect 19064 34342 19116 34348
rect 19156 34400 19208 34406
rect 19156 34342 19208 34348
rect 19076 34202 19104 34342
rect 19064 34196 19116 34202
rect 19064 34138 19116 34144
rect 19156 34128 19208 34134
rect 19156 34070 19208 34076
rect 19064 33856 19116 33862
rect 19064 33798 19116 33804
rect 19076 33590 19104 33798
rect 19064 33584 19116 33590
rect 19064 33526 19116 33532
rect 19168 33046 19196 34070
rect 19156 33040 19208 33046
rect 19156 32982 19208 32988
rect 19260 32910 19288 34546
rect 19444 33969 19472 35550
rect 19524 35488 19576 35494
rect 19524 35430 19576 35436
rect 20168 35488 20220 35494
rect 20168 35430 20220 35436
rect 19536 35057 19564 35430
rect 19522 35048 19578 35057
rect 19522 34983 19578 34992
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19984 34536 20036 34542
rect 19984 34478 20036 34484
rect 20076 34536 20128 34542
rect 20076 34478 20128 34484
rect 19522 34232 19578 34241
rect 19522 34167 19578 34176
rect 19430 33960 19486 33969
rect 19430 33895 19486 33904
rect 19536 33862 19564 34167
rect 19890 34096 19946 34105
rect 19890 34031 19892 34040
rect 19944 34031 19946 34040
rect 19892 34002 19944 34008
rect 19524 33856 19576 33862
rect 19524 33798 19576 33804
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19996 33590 20024 34478
rect 20088 33658 20116 34478
rect 20180 33998 20208 35430
rect 20352 35148 20404 35154
rect 20352 35090 20404 35096
rect 20168 33992 20220 33998
rect 20168 33934 20220 33940
rect 20076 33652 20128 33658
rect 20076 33594 20128 33600
rect 19984 33584 20036 33590
rect 19984 33526 20036 33532
rect 19800 33448 19852 33454
rect 19800 33390 19852 33396
rect 19340 33380 19392 33386
rect 19340 33322 19392 33328
rect 19248 32904 19300 32910
rect 19248 32846 19300 32852
rect 19156 32836 19208 32842
rect 19156 32778 19208 32784
rect 19168 32434 19196 32778
rect 19246 32600 19302 32609
rect 19246 32535 19302 32544
rect 19260 32502 19288 32535
rect 19248 32496 19300 32502
rect 19248 32438 19300 32444
rect 19156 32428 19208 32434
rect 19156 32370 19208 32376
rect 19062 32192 19118 32201
rect 19062 32127 19118 32136
rect 18880 31748 18932 31754
rect 18880 31690 18932 31696
rect 18604 31476 18656 31482
rect 18604 31418 18656 31424
rect 18420 31204 18472 31210
rect 18420 31146 18472 31152
rect 18616 31142 18644 31418
rect 18880 31272 18932 31278
rect 18880 31214 18932 31220
rect 18512 31136 18564 31142
rect 18512 31078 18564 31084
rect 18604 31136 18656 31142
rect 18604 31078 18656 31084
rect 18420 30932 18472 30938
rect 18420 30874 18472 30880
rect 18432 30841 18460 30874
rect 18418 30832 18474 30841
rect 18418 30767 18474 30776
rect 18432 30734 18460 30767
rect 18420 30728 18472 30734
rect 18420 30670 18472 30676
rect 18420 30592 18472 30598
rect 18420 30534 18472 30540
rect 18328 30048 18380 30054
rect 18328 29990 18380 29996
rect 18340 28966 18368 29990
rect 18432 29238 18460 30534
rect 18524 29850 18552 31078
rect 18892 30705 18920 31214
rect 18878 30696 18934 30705
rect 18788 30660 18840 30666
rect 18878 30631 18934 30640
rect 18788 30602 18840 30608
rect 18800 30394 18828 30602
rect 19076 30394 19104 32127
rect 19352 30598 19380 33322
rect 19524 33312 19576 33318
rect 19616 33312 19668 33318
rect 19524 33254 19576 33260
rect 19614 33280 19616 33289
rect 19668 33280 19670 33289
rect 19536 33114 19564 33254
rect 19614 33215 19670 33224
rect 19524 33108 19576 33114
rect 19524 33050 19576 33056
rect 19812 32774 19840 33390
rect 20166 33144 20222 33153
rect 20166 33079 20168 33088
rect 20220 33079 20222 33088
rect 20168 33050 20220 33056
rect 19800 32768 19852 32774
rect 19800 32710 19852 32716
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 20076 32360 20128 32366
rect 20076 32302 20128 32308
rect 20088 31890 20116 32302
rect 20168 32224 20220 32230
rect 20168 32166 20220 32172
rect 20076 31884 20128 31890
rect 20076 31826 20128 31832
rect 19430 31784 19486 31793
rect 19430 31719 19486 31728
rect 19984 31748 20036 31754
rect 19444 31521 19472 31719
rect 19984 31690 20036 31696
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19430 31512 19486 31521
rect 19574 31515 19882 31524
rect 19996 31482 20024 31690
rect 19430 31447 19486 31456
rect 19984 31476 20036 31482
rect 19984 31418 20036 31424
rect 20180 30784 20208 32166
rect 20364 30920 20392 35090
rect 20444 34944 20496 34950
rect 20444 34886 20496 34892
rect 20088 30756 20208 30784
rect 20272 30892 20392 30920
rect 19984 30660 20036 30666
rect 19984 30602 20036 30608
rect 19340 30592 19392 30598
rect 19392 30552 19472 30580
rect 19340 30534 19392 30540
rect 18788 30388 18840 30394
rect 18788 30330 18840 30336
rect 19064 30388 19116 30394
rect 19064 30330 19116 30336
rect 18512 29844 18564 29850
rect 18512 29786 18564 29792
rect 18800 29714 18828 30330
rect 19340 30320 19392 30326
rect 19340 30262 19392 30268
rect 19156 30184 19208 30190
rect 19156 30126 19208 30132
rect 18788 29708 18840 29714
rect 18788 29650 18840 29656
rect 18972 29708 19024 29714
rect 18972 29650 19024 29656
rect 18696 29572 18748 29578
rect 18696 29514 18748 29520
rect 18420 29232 18472 29238
rect 18420 29174 18472 29180
rect 18708 29102 18736 29514
rect 18696 29096 18748 29102
rect 18696 29038 18748 29044
rect 18328 28960 18380 28966
rect 18328 28902 18380 28908
rect 18340 28014 18368 28902
rect 18602 28656 18658 28665
rect 18602 28591 18658 28600
rect 18616 28014 18644 28591
rect 18328 28008 18380 28014
rect 18328 27950 18380 27956
rect 18512 28008 18564 28014
rect 18512 27950 18564 27956
rect 18604 28008 18656 28014
rect 18604 27950 18656 27956
rect 18420 26920 18472 26926
rect 18420 26862 18472 26868
rect 18432 26761 18460 26862
rect 18418 26752 18474 26761
rect 18418 26687 18474 26696
rect 18236 26580 18288 26586
rect 18236 26522 18288 26528
rect 18420 26580 18472 26586
rect 18420 26522 18472 26528
rect 18248 26246 18276 26522
rect 18236 26240 18288 26246
rect 18236 26182 18288 26188
rect 17960 25900 18012 25906
rect 17960 25842 18012 25848
rect 18144 25900 18196 25906
rect 18144 25842 18196 25848
rect 18156 24818 18184 25842
rect 18432 25362 18460 26522
rect 18524 25922 18552 27950
rect 18880 27940 18932 27946
rect 18880 27882 18932 27888
rect 18788 27600 18840 27606
rect 18788 27542 18840 27548
rect 18696 27396 18748 27402
rect 18696 27338 18748 27344
rect 18708 26042 18736 27338
rect 18800 26382 18828 27542
rect 18788 26376 18840 26382
rect 18788 26318 18840 26324
rect 18696 26036 18748 26042
rect 18696 25978 18748 25984
rect 18524 25894 18736 25922
rect 18420 25356 18472 25362
rect 18420 25298 18472 25304
rect 18144 24812 18196 24818
rect 18144 24754 18196 24760
rect 18052 23792 18104 23798
rect 18052 23734 18104 23740
rect 18064 23322 18092 23734
rect 18052 23316 18104 23322
rect 18052 23258 18104 23264
rect 17868 23248 17920 23254
rect 17868 23190 17920 23196
rect 17776 23112 17828 23118
rect 17776 23054 17828 23060
rect 18236 23112 18288 23118
rect 18236 23054 18288 23060
rect 17684 23044 17736 23050
rect 17684 22986 17736 22992
rect 18050 22808 18106 22817
rect 18050 22743 18052 22752
rect 18104 22743 18106 22752
rect 18052 22714 18104 22720
rect 17592 22636 17644 22642
rect 17592 22578 17644 22584
rect 17604 21418 17632 22578
rect 17960 21616 18012 21622
rect 17960 21558 18012 21564
rect 17684 21548 17736 21554
rect 17684 21490 17736 21496
rect 17592 21412 17644 21418
rect 17592 21354 17644 21360
rect 17696 21350 17724 21490
rect 17972 21418 18000 21558
rect 17960 21412 18012 21418
rect 17960 21354 18012 21360
rect 17684 21344 17736 21350
rect 17684 21286 17736 21292
rect 17500 21072 17552 21078
rect 17500 21014 17552 21020
rect 17500 20936 17552 20942
rect 17500 20878 17552 20884
rect 17316 20800 17368 20806
rect 17316 20742 17368 20748
rect 17224 19372 17276 19378
rect 17224 19314 17276 19320
rect 16488 18964 16540 18970
rect 16488 18906 16540 18912
rect 16500 17542 16528 18906
rect 17328 18698 17356 20742
rect 17512 20466 17540 20878
rect 17500 20460 17552 20466
rect 17500 20402 17552 20408
rect 17316 18692 17368 18698
rect 17316 18634 17368 18640
rect 16488 17536 16540 17542
rect 16488 17478 16540 17484
rect 16408 16546 16528 16574
rect 16120 12640 16172 12646
rect 16120 12582 16172 12588
rect 15568 12232 15620 12238
rect 15568 12174 15620 12180
rect 15200 2576 15252 2582
rect 15200 2518 15252 2524
rect 16132 2446 16160 12582
rect 16500 2650 16528 16546
rect 16856 12368 16908 12374
rect 16856 12310 16908 12316
rect 16488 2644 16540 2650
rect 16488 2586 16540 2592
rect 16868 2446 16896 12310
rect 17696 8838 17724 21286
rect 17868 20460 17920 20466
rect 17868 20402 17920 20408
rect 17880 20262 17908 20402
rect 17868 20256 17920 20262
rect 17868 20198 17920 20204
rect 17880 19786 17908 20198
rect 17972 20058 18000 21354
rect 18248 21078 18276 23054
rect 18432 22982 18460 25298
rect 18512 25220 18564 25226
rect 18708 25208 18736 25894
rect 18800 25276 18828 26318
rect 18892 25498 18920 27882
rect 18984 26926 19012 29650
rect 19064 29504 19116 29510
rect 19064 29446 19116 29452
rect 18972 26920 19024 26926
rect 18972 26862 19024 26868
rect 18880 25492 18932 25498
rect 18880 25434 18932 25440
rect 18800 25248 18920 25276
rect 18708 25180 18828 25208
rect 18512 25162 18564 25168
rect 18524 24954 18552 25162
rect 18512 24948 18564 24954
rect 18512 24890 18564 24896
rect 18604 24132 18656 24138
rect 18604 24074 18656 24080
rect 18512 24064 18564 24070
rect 18512 24006 18564 24012
rect 18420 22976 18472 22982
rect 18420 22918 18472 22924
rect 18328 22568 18380 22574
rect 18328 22510 18380 22516
rect 18340 22098 18368 22510
rect 18328 22092 18380 22098
rect 18328 22034 18380 22040
rect 18340 21690 18368 22034
rect 18328 21684 18380 21690
rect 18328 21626 18380 21632
rect 18236 21072 18288 21078
rect 18236 21014 18288 21020
rect 17960 20052 18012 20058
rect 17960 19994 18012 20000
rect 17868 19780 17920 19786
rect 17868 19722 17920 19728
rect 18524 10742 18552 24006
rect 18616 23866 18644 24074
rect 18604 23860 18656 23866
rect 18604 23802 18656 23808
rect 18604 22976 18656 22982
rect 18604 22918 18656 22924
rect 18616 16590 18644 22918
rect 18696 20800 18748 20806
rect 18696 20742 18748 20748
rect 18604 16584 18656 16590
rect 18604 16526 18656 16532
rect 18512 10736 18564 10742
rect 18512 10678 18564 10684
rect 17684 8832 17736 8838
rect 17684 8774 17736 8780
rect 18708 3466 18736 20742
rect 18800 11898 18828 25180
rect 18892 20942 18920 25248
rect 19076 24206 19104 29446
rect 19168 29306 19196 30126
rect 19156 29300 19208 29306
rect 19156 29242 19208 29248
rect 19248 29232 19300 29238
rect 19248 29174 19300 29180
rect 19260 28762 19288 29174
rect 19352 29034 19380 30262
rect 19444 29220 19472 30552
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19524 30320 19576 30326
rect 19524 30262 19576 30268
rect 19800 30320 19852 30326
rect 19800 30262 19852 30268
rect 19536 29850 19564 30262
rect 19812 30122 19840 30262
rect 19800 30116 19852 30122
rect 19800 30058 19852 30064
rect 19892 30048 19944 30054
rect 19892 29990 19944 29996
rect 19524 29844 19576 29850
rect 19524 29786 19576 29792
rect 19904 29510 19932 29990
rect 19892 29504 19944 29510
rect 19892 29446 19944 29452
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19524 29232 19576 29238
rect 19444 29192 19524 29220
rect 19340 29028 19392 29034
rect 19340 28970 19392 28976
rect 19248 28756 19300 28762
rect 19248 28698 19300 28704
rect 19352 27962 19380 28970
rect 19444 28150 19472 29192
rect 19524 29174 19576 29180
rect 19614 29200 19670 29209
rect 19614 29135 19670 29144
rect 19628 28558 19656 29135
rect 19996 28626 20024 30602
rect 20088 30569 20116 30756
rect 20074 30560 20130 30569
rect 20074 30495 20130 30504
rect 20076 30184 20128 30190
rect 20076 30126 20128 30132
rect 20088 29714 20116 30126
rect 20076 29708 20128 29714
rect 20076 29650 20128 29656
rect 20272 29578 20300 30892
rect 20350 30560 20406 30569
rect 20350 30495 20406 30504
rect 20076 29572 20128 29578
rect 20076 29514 20128 29520
rect 20260 29572 20312 29578
rect 20260 29514 20312 29520
rect 19892 28620 19944 28626
rect 19892 28562 19944 28568
rect 19984 28620 20036 28626
rect 19984 28562 20036 28568
rect 19524 28552 19576 28558
rect 19524 28494 19576 28500
rect 19616 28552 19668 28558
rect 19616 28494 19668 28500
rect 19536 28422 19564 28494
rect 19904 28472 19932 28562
rect 19904 28444 20024 28472
rect 19524 28416 19576 28422
rect 19524 28358 19576 28364
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19432 28144 19484 28150
rect 19432 28086 19484 28092
rect 19352 27934 19472 27962
rect 19340 27328 19392 27334
rect 19340 27270 19392 27276
rect 19352 27062 19380 27270
rect 19340 27056 19392 27062
rect 19340 26998 19392 27004
rect 19444 27010 19472 27934
rect 19996 27878 20024 28444
rect 19524 27872 19576 27878
rect 19524 27814 19576 27820
rect 19984 27872 20036 27878
rect 19984 27814 20036 27820
rect 19536 27538 19564 27814
rect 19524 27532 19576 27538
rect 19524 27474 19576 27480
rect 19984 27464 20036 27470
rect 19984 27406 20036 27412
rect 19996 27334 20024 27406
rect 19984 27328 20036 27334
rect 19984 27270 20036 27276
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19800 27056 19852 27062
rect 19706 27024 19762 27033
rect 19444 26982 19564 27010
rect 19432 26920 19484 26926
rect 19432 26862 19484 26868
rect 19444 26602 19472 26862
rect 19536 26790 19564 26982
rect 19800 26998 19852 27004
rect 19706 26959 19762 26968
rect 19524 26784 19576 26790
rect 19524 26726 19576 26732
rect 19444 26574 19656 26602
rect 19340 26376 19392 26382
rect 19338 26344 19340 26353
rect 19628 26364 19656 26574
rect 19392 26344 19394 26353
rect 19338 26279 19394 26288
rect 19444 26336 19656 26364
rect 19156 26240 19208 26246
rect 19156 26182 19208 26188
rect 19168 25294 19196 26182
rect 19340 25968 19392 25974
rect 19340 25910 19392 25916
rect 19352 25770 19380 25910
rect 19340 25764 19392 25770
rect 19340 25706 19392 25712
rect 19156 25288 19208 25294
rect 19156 25230 19208 25236
rect 19340 25288 19392 25294
rect 19340 25230 19392 25236
rect 19248 25152 19300 25158
rect 19248 25094 19300 25100
rect 19260 24274 19288 25094
rect 19248 24268 19300 24274
rect 19248 24210 19300 24216
rect 19064 24200 19116 24206
rect 19064 24142 19116 24148
rect 19156 23316 19208 23322
rect 19156 23258 19208 23264
rect 18972 23112 19024 23118
rect 18972 23054 19024 23060
rect 18984 22030 19012 23054
rect 18972 22024 19024 22030
rect 18972 21966 19024 21972
rect 18984 21418 19012 21966
rect 19064 21548 19116 21554
rect 19064 21490 19116 21496
rect 18972 21412 19024 21418
rect 18972 21354 19024 21360
rect 18880 20936 18932 20942
rect 18880 20878 18932 20884
rect 19076 20874 19104 21490
rect 19064 20868 19116 20874
rect 19064 20810 19116 20816
rect 19168 20602 19196 23258
rect 19352 23118 19380 25230
rect 19444 25140 19472 26336
rect 19524 26240 19576 26246
rect 19720 26228 19748 26959
rect 19812 26246 19840 26998
rect 19576 26200 19748 26228
rect 19800 26240 19852 26246
rect 19524 26182 19576 26188
rect 19800 26182 19852 26188
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19524 25356 19576 25362
rect 19524 25298 19576 25304
rect 19536 25140 19564 25298
rect 19444 25112 19564 25140
rect 19444 24750 19472 25112
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19892 24812 19944 24818
rect 19892 24754 19944 24760
rect 19432 24744 19484 24750
rect 19432 24686 19484 24692
rect 19904 24138 19932 24754
rect 19892 24132 19944 24138
rect 19892 24074 19944 24080
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19996 23322 20024 27270
rect 20088 25974 20116 29514
rect 20258 29336 20314 29345
rect 20258 29271 20314 29280
rect 20168 28552 20220 28558
rect 20168 28494 20220 28500
rect 20076 25968 20128 25974
rect 20076 25910 20128 25916
rect 20180 25922 20208 28494
rect 20272 26926 20300 29271
rect 20364 27674 20392 30495
rect 20456 29714 20484 34886
rect 20548 31793 20576 36518
rect 20824 36038 20852 36654
rect 22192 36644 22244 36650
rect 22192 36586 22244 36592
rect 22204 36378 22232 36586
rect 22192 36372 22244 36378
rect 22192 36314 22244 36320
rect 20812 36032 20864 36038
rect 20812 35974 20864 35980
rect 21640 36032 21692 36038
rect 21640 35974 21692 35980
rect 21088 35828 21140 35834
rect 21088 35770 21140 35776
rect 21100 35290 21128 35770
rect 21652 35766 21680 35974
rect 21640 35760 21692 35766
rect 21640 35702 21692 35708
rect 21088 35284 21140 35290
rect 21088 35226 21140 35232
rect 21100 34746 21128 35226
rect 21364 34944 21416 34950
rect 21364 34886 21416 34892
rect 21088 34740 21140 34746
rect 21088 34682 21140 34688
rect 20720 34604 20772 34610
rect 20720 34546 20772 34552
rect 20812 34604 20864 34610
rect 20812 34546 20864 34552
rect 20626 34096 20682 34105
rect 20626 34031 20628 34040
rect 20680 34031 20682 34040
rect 20628 34002 20680 34008
rect 20732 33658 20760 34546
rect 20720 33652 20772 33658
rect 20720 33594 20772 33600
rect 20732 32910 20760 33594
rect 20720 32904 20772 32910
rect 20720 32846 20772 32852
rect 20720 32496 20772 32502
rect 20720 32438 20772 32444
rect 20732 31958 20760 32438
rect 20720 31952 20772 31958
rect 20720 31894 20772 31900
rect 20534 31784 20590 31793
rect 20534 31719 20590 31728
rect 20548 31346 20576 31719
rect 20628 31408 20680 31414
rect 20628 31350 20680 31356
rect 20536 31340 20588 31346
rect 20536 31282 20588 31288
rect 20548 30802 20576 31282
rect 20536 30796 20588 30802
rect 20536 30738 20588 30744
rect 20444 29708 20496 29714
rect 20444 29650 20496 29656
rect 20444 29572 20496 29578
rect 20444 29514 20496 29520
rect 20456 29345 20484 29514
rect 20442 29336 20498 29345
rect 20442 29271 20498 29280
rect 20444 29232 20496 29238
rect 20444 29174 20496 29180
rect 20456 28762 20484 29174
rect 20444 28756 20496 28762
rect 20444 28698 20496 28704
rect 20548 28422 20576 30738
rect 20536 28416 20588 28422
rect 20536 28358 20588 28364
rect 20444 28076 20496 28082
rect 20444 28018 20496 28024
rect 20456 27946 20484 28018
rect 20444 27940 20496 27946
rect 20444 27882 20496 27888
rect 20352 27668 20404 27674
rect 20352 27610 20404 27616
rect 20260 26920 20312 26926
rect 20260 26862 20312 26868
rect 20272 26790 20300 26862
rect 20260 26784 20312 26790
rect 20260 26726 20312 26732
rect 20456 26234 20484 27882
rect 20640 27538 20668 31350
rect 20720 30592 20772 30598
rect 20720 30534 20772 30540
rect 20732 30394 20760 30534
rect 20720 30388 20772 30394
rect 20720 30330 20772 30336
rect 20720 30116 20772 30122
rect 20720 30058 20772 30064
rect 20732 28082 20760 30058
rect 20824 29170 20852 34546
rect 21100 34202 21128 34682
rect 21088 34196 21140 34202
rect 21088 34138 21140 34144
rect 20904 33040 20956 33046
rect 20904 32982 20956 32988
rect 20916 32434 20944 32982
rect 20996 32904 21048 32910
rect 20996 32846 21048 32852
rect 21086 32872 21142 32881
rect 20904 32428 20956 32434
rect 20904 32370 20956 32376
rect 20916 31346 20944 32370
rect 21008 31822 21036 32846
rect 21086 32807 21088 32816
rect 21140 32807 21142 32816
rect 21088 32778 21140 32784
rect 20996 31816 21048 31822
rect 20996 31758 21048 31764
rect 21272 31816 21324 31822
rect 21272 31758 21324 31764
rect 20996 31680 21048 31686
rect 20996 31622 21048 31628
rect 21008 31482 21036 31622
rect 21284 31482 21312 31758
rect 20996 31476 21048 31482
rect 20996 31418 21048 31424
rect 21272 31476 21324 31482
rect 21272 31418 21324 31424
rect 20904 31340 20956 31346
rect 20904 31282 20956 31288
rect 20916 30734 20944 31282
rect 21376 30977 21404 34886
rect 21652 32570 21680 35702
rect 21916 34400 21968 34406
rect 21916 34342 21968 34348
rect 21824 33856 21876 33862
rect 21824 33798 21876 33804
rect 21836 32978 21864 33798
rect 21928 33658 21956 34342
rect 22008 33924 22060 33930
rect 22008 33866 22060 33872
rect 21916 33652 21968 33658
rect 21916 33594 21968 33600
rect 21824 32972 21876 32978
rect 21824 32914 21876 32920
rect 21640 32564 21692 32570
rect 21640 32506 21692 32512
rect 21362 30968 21418 30977
rect 21362 30903 21418 30912
rect 20904 30728 20956 30734
rect 20904 30670 20956 30676
rect 21548 30252 21600 30258
rect 21548 30194 21600 30200
rect 20904 30116 20956 30122
rect 20904 30058 20956 30064
rect 20916 29782 20944 30058
rect 20904 29776 20956 29782
rect 20904 29718 20956 29724
rect 20996 29504 21048 29510
rect 20996 29446 21048 29452
rect 21008 29306 21036 29446
rect 20996 29300 21048 29306
rect 20996 29242 21048 29248
rect 20812 29164 20864 29170
rect 20812 29106 20864 29112
rect 20824 28558 20852 29106
rect 21560 29034 21588 30194
rect 21916 29640 21968 29646
rect 21916 29582 21968 29588
rect 21732 29504 21784 29510
rect 21732 29446 21784 29452
rect 21744 29238 21772 29446
rect 21732 29232 21784 29238
rect 21732 29174 21784 29180
rect 21548 29028 21600 29034
rect 21548 28970 21600 28976
rect 20812 28552 20864 28558
rect 20812 28494 20864 28500
rect 20720 28076 20772 28082
rect 20720 28018 20772 28024
rect 21364 28008 21416 28014
rect 21364 27950 21416 27956
rect 21272 27600 21324 27606
rect 21272 27542 21324 27548
rect 20628 27532 20680 27538
rect 20628 27474 20680 27480
rect 20536 27396 20588 27402
rect 20536 27338 20588 27344
rect 20548 26450 20576 27338
rect 20640 26926 20668 27474
rect 20996 27396 21048 27402
rect 20996 27338 21048 27344
rect 20720 27124 20772 27130
rect 20720 27066 20772 27072
rect 20628 26920 20680 26926
rect 20628 26862 20680 26868
rect 20640 26518 20668 26862
rect 20628 26512 20680 26518
rect 20628 26454 20680 26460
rect 20536 26444 20588 26450
rect 20536 26386 20588 26392
rect 20456 26206 20576 26234
rect 20180 25894 20392 25922
rect 20076 25832 20128 25838
rect 20076 25774 20128 25780
rect 20168 25832 20220 25838
rect 20168 25774 20220 25780
rect 20088 24682 20116 25774
rect 20180 24954 20208 25774
rect 20260 25220 20312 25226
rect 20260 25162 20312 25168
rect 20168 24948 20220 24954
rect 20168 24890 20220 24896
rect 20076 24676 20128 24682
rect 20076 24618 20128 24624
rect 20180 24290 20208 24890
rect 20272 24750 20300 25162
rect 20260 24744 20312 24750
rect 20260 24686 20312 24692
rect 20180 24262 20300 24290
rect 19984 23316 20036 23322
rect 19984 23258 20036 23264
rect 19340 23112 19392 23118
rect 19340 23054 19392 23060
rect 19352 22094 19380 23054
rect 20076 22976 20128 22982
rect 20076 22918 20128 22924
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 20088 22574 20116 22918
rect 20168 22704 20220 22710
rect 20168 22646 20220 22652
rect 20076 22568 20128 22574
rect 20076 22510 20128 22516
rect 19352 22066 19472 22094
rect 19444 21894 19472 22066
rect 19432 21888 19484 21894
rect 19432 21830 19484 21836
rect 19984 21888 20036 21894
rect 19984 21830 20036 21836
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19996 21146 20024 21830
rect 20180 21690 20208 22646
rect 20168 21684 20220 21690
rect 20168 21626 20220 21632
rect 19984 21140 20036 21146
rect 19984 21082 20036 21088
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19156 20596 19208 20602
rect 19156 20538 19208 20544
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 20076 13184 20128 13190
rect 20076 13126 20128 13132
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 18788 11892 18840 11898
rect 18788 11834 18840 11840
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19984 9716 20036 9722
rect 19984 9658 20036 9664
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 18696 3460 18748 3466
rect 18696 3402 18748 3408
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19996 3058 20024 9658
rect 19984 3052 20036 3058
rect 19984 2994 20036 3000
rect 19996 2514 20024 2994
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 20088 2446 20116 13126
rect 20272 9654 20300 24262
rect 20364 24206 20392 25894
rect 20352 24200 20404 24206
rect 20352 24142 20404 24148
rect 20364 23798 20392 24142
rect 20352 23792 20404 23798
rect 20352 23734 20404 23740
rect 20364 22658 20392 23734
rect 20364 22630 20484 22658
rect 20352 22568 20404 22574
rect 20352 22510 20404 22516
rect 20364 22098 20392 22510
rect 20456 22234 20484 22630
rect 20444 22228 20496 22234
rect 20444 22170 20496 22176
rect 20352 22092 20404 22098
rect 20548 22094 20576 26206
rect 20732 26042 20760 27066
rect 20904 26376 20956 26382
rect 20902 26344 20904 26353
rect 20956 26344 20958 26353
rect 20902 26279 20958 26288
rect 21008 26042 21036 27338
rect 21284 27334 21312 27542
rect 21272 27328 21324 27334
rect 21272 27270 21324 27276
rect 21376 26994 21404 27950
rect 21364 26988 21416 26994
rect 21364 26930 21416 26936
rect 21376 26466 21404 26930
rect 21284 26438 21404 26466
rect 20720 26036 20772 26042
rect 20720 25978 20772 25984
rect 20996 26036 21048 26042
rect 20996 25978 21048 25984
rect 20628 25900 20680 25906
rect 20628 25842 20680 25848
rect 20640 25430 20668 25842
rect 20628 25424 20680 25430
rect 20628 25366 20680 25372
rect 20640 23730 20668 25366
rect 21284 24818 21312 26438
rect 21364 26308 21416 26314
rect 21364 26250 21416 26256
rect 21376 24818 21404 26250
rect 21560 24818 21588 28970
rect 21732 28620 21784 28626
rect 21732 28562 21784 28568
rect 21744 28082 21772 28562
rect 21732 28076 21784 28082
rect 21732 28018 21784 28024
rect 21640 27464 21692 27470
rect 21640 27406 21692 27412
rect 21652 26858 21680 27406
rect 21640 26852 21692 26858
rect 21640 26794 21692 26800
rect 21272 24812 21324 24818
rect 21272 24754 21324 24760
rect 21364 24812 21416 24818
rect 21364 24754 21416 24760
rect 21548 24812 21600 24818
rect 21548 24754 21600 24760
rect 20720 24676 20772 24682
rect 20772 24636 20852 24664
rect 20720 24618 20772 24624
rect 20628 23724 20680 23730
rect 20628 23666 20680 23672
rect 20720 23520 20772 23526
rect 20720 23462 20772 23468
rect 20732 23118 20760 23462
rect 20720 23112 20772 23118
rect 20720 23054 20772 23060
rect 20824 22710 20852 24636
rect 21284 24274 21312 24754
rect 21272 24268 21324 24274
rect 21272 24210 21324 24216
rect 21180 24132 21232 24138
rect 21180 24074 21232 24080
rect 20904 23112 20956 23118
rect 20904 23054 20956 23060
rect 20812 22704 20864 22710
rect 20812 22646 20864 22652
rect 20352 22034 20404 22040
rect 20456 22066 20576 22094
rect 20456 13530 20484 22066
rect 20916 18834 20944 23054
rect 21192 22098 21220 24074
rect 21284 23594 21312 24210
rect 21744 23866 21772 28018
rect 21824 27328 21876 27334
rect 21824 27270 21876 27276
rect 21836 26858 21864 27270
rect 21824 26852 21876 26858
rect 21824 26794 21876 26800
rect 21928 26738 21956 29582
rect 22020 27606 22048 33866
rect 22468 32224 22520 32230
rect 22468 32166 22520 32172
rect 22480 31278 22508 32166
rect 22100 31272 22152 31278
rect 22100 31214 22152 31220
rect 22468 31272 22520 31278
rect 22468 31214 22520 31220
rect 22112 30598 22140 31214
rect 22100 30592 22152 30598
rect 22100 30534 22152 30540
rect 22112 30326 22140 30534
rect 22100 30320 22152 30326
rect 22100 30262 22152 30268
rect 22112 29714 22140 30262
rect 22100 29708 22152 29714
rect 22100 29650 22152 29656
rect 22008 27600 22060 27606
rect 22008 27542 22060 27548
rect 21836 26710 21956 26738
rect 21732 23860 21784 23866
rect 21732 23802 21784 23808
rect 21272 23588 21324 23594
rect 21272 23530 21324 23536
rect 21180 22092 21232 22098
rect 21180 22034 21232 22040
rect 21456 21616 21508 21622
rect 21456 21558 21508 21564
rect 21468 20058 21496 21558
rect 21456 20052 21508 20058
rect 21456 19994 21508 20000
rect 21468 19854 21496 19994
rect 21456 19848 21508 19854
rect 21456 19790 21508 19796
rect 20904 18828 20956 18834
rect 20904 18770 20956 18776
rect 20444 13524 20496 13530
rect 20444 13466 20496 13472
rect 20456 13326 20484 13466
rect 20444 13320 20496 13326
rect 20444 13262 20496 13268
rect 21836 12986 21864 26710
rect 22112 25294 22140 29650
rect 22560 28756 22612 28762
rect 22560 28698 22612 28704
rect 22572 27878 22600 28698
rect 22560 27872 22612 27878
rect 22560 27814 22612 27820
rect 22652 27056 22704 27062
rect 22652 26998 22704 27004
rect 22468 26852 22520 26858
rect 22468 26794 22520 26800
rect 22480 26586 22508 26794
rect 22664 26586 22692 26998
rect 22468 26580 22520 26586
rect 22468 26522 22520 26528
rect 22652 26580 22704 26586
rect 22652 26522 22704 26528
rect 22756 26382 22784 37402
rect 23860 37262 23888 37402
rect 23848 37256 23900 37262
rect 23848 37198 23900 37204
rect 23204 37188 23256 37194
rect 23204 37130 23256 37136
rect 23112 36100 23164 36106
rect 23112 36042 23164 36048
rect 23020 35012 23072 35018
rect 23020 34954 23072 34960
rect 22928 34740 22980 34746
rect 22928 34682 22980 34688
rect 22940 34202 22968 34682
rect 22928 34196 22980 34202
rect 22928 34138 22980 34144
rect 22940 33658 22968 34138
rect 22928 33652 22980 33658
rect 22928 33594 22980 33600
rect 22940 33114 22968 33594
rect 22928 33108 22980 33114
rect 22928 33050 22980 33056
rect 22940 32570 22968 33050
rect 22928 32564 22980 32570
rect 22928 32506 22980 32512
rect 22940 32026 22968 32506
rect 22928 32020 22980 32026
rect 22928 31962 22980 31968
rect 22940 31482 22968 31962
rect 22928 31476 22980 31482
rect 22928 31418 22980 31424
rect 23032 30938 23060 34954
rect 23124 34678 23152 36042
rect 23112 34672 23164 34678
rect 23112 34614 23164 34620
rect 23020 30932 23072 30938
rect 23020 30874 23072 30880
rect 23032 30666 23060 30874
rect 23020 30660 23072 30666
rect 23020 30602 23072 30608
rect 22928 30048 22980 30054
rect 22928 29990 22980 29996
rect 22744 26376 22796 26382
rect 22744 26318 22796 26324
rect 22756 26194 22784 26318
rect 22756 26166 22876 26194
rect 22744 26036 22796 26042
rect 22744 25978 22796 25984
rect 22652 25832 22704 25838
rect 22652 25774 22704 25780
rect 22664 25498 22692 25774
rect 22652 25492 22704 25498
rect 22652 25434 22704 25440
rect 22100 25288 22152 25294
rect 22100 25230 22152 25236
rect 22192 25220 22244 25226
rect 22192 25162 22244 25168
rect 21916 24744 21968 24750
rect 21916 24686 21968 24692
rect 21928 24274 21956 24686
rect 22204 24274 22232 25162
rect 22756 24954 22784 25978
rect 22848 25906 22876 26166
rect 22836 25900 22888 25906
rect 22836 25842 22888 25848
rect 22744 24948 22796 24954
rect 22744 24890 22796 24896
rect 21916 24268 21968 24274
rect 21916 24210 21968 24216
rect 22192 24268 22244 24274
rect 22192 24210 22244 24216
rect 22204 22778 22232 24210
rect 22192 22772 22244 22778
rect 22192 22714 22244 22720
rect 22848 22094 22876 25842
rect 22940 23118 22968 29990
rect 23216 29306 23244 37130
rect 25148 37126 25176 39200
rect 27080 37126 27108 39200
rect 28908 37256 28960 37262
rect 28908 37198 28960 37204
rect 23296 37120 23348 37126
rect 23296 37062 23348 37068
rect 24676 37120 24728 37126
rect 24676 37062 24728 37068
rect 25136 37120 25188 37126
rect 25136 37062 25188 37068
rect 26516 37120 26568 37126
rect 26516 37062 26568 37068
rect 27068 37120 27120 37126
rect 27068 37062 27120 37068
rect 23308 36650 23336 37062
rect 23296 36644 23348 36650
rect 23296 36586 23348 36592
rect 23308 36378 23336 36586
rect 23296 36372 23348 36378
rect 23296 36314 23348 36320
rect 24584 36032 24636 36038
rect 24584 35974 24636 35980
rect 23388 34944 23440 34950
rect 23388 34886 23440 34892
rect 23400 34746 23428 34886
rect 23388 34740 23440 34746
rect 23388 34682 23440 34688
rect 24596 33590 24624 35974
rect 24584 33584 24636 33590
rect 24584 33526 24636 33532
rect 23662 33416 23718 33425
rect 23662 33351 23664 33360
rect 23716 33351 23718 33360
rect 23664 33322 23716 33328
rect 23296 32768 23348 32774
rect 23296 32710 23348 32716
rect 23204 29300 23256 29306
rect 23204 29242 23256 29248
rect 23204 29028 23256 29034
rect 23204 28970 23256 28976
rect 23216 27316 23244 28970
rect 23308 28762 23336 32710
rect 23572 32292 23624 32298
rect 23572 32234 23624 32240
rect 23388 29028 23440 29034
rect 23388 28970 23440 28976
rect 23296 28756 23348 28762
rect 23296 28698 23348 28704
rect 23400 28150 23428 28970
rect 23388 28144 23440 28150
rect 23388 28086 23440 28092
rect 23400 27946 23428 28086
rect 23388 27940 23440 27946
rect 23388 27882 23440 27888
rect 23388 27328 23440 27334
rect 23216 27288 23388 27316
rect 23388 27270 23440 27276
rect 23296 27056 23348 27062
rect 23400 27033 23428 27270
rect 23296 26998 23348 27004
rect 23386 27024 23442 27033
rect 23308 26586 23336 26998
rect 23386 26959 23442 26968
rect 23584 26926 23612 32234
rect 24124 30728 24176 30734
rect 24124 30670 24176 30676
rect 24136 29170 24164 30670
rect 24124 29164 24176 29170
rect 24124 29106 24176 29112
rect 23756 28688 23808 28694
rect 23756 28630 23808 28636
rect 23768 28218 23796 28630
rect 23756 28212 23808 28218
rect 23756 28154 23808 28160
rect 24688 28082 24716 37062
rect 24768 36304 24820 36310
rect 24768 36246 24820 36252
rect 24780 33658 24808 36246
rect 25688 36032 25740 36038
rect 25688 35974 25740 35980
rect 25320 35624 25372 35630
rect 25318 35592 25320 35601
rect 25372 35592 25374 35601
rect 25318 35527 25374 35536
rect 24768 33652 24820 33658
rect 24768 33594 24820 33600
rect 25700 30802 25728 35974
rect 25688 30796 25740 30802
rect 25688 30738 25740 30744
rect 24676 28076 24728 28082
rect 24676 28018 24728 28024
rect 23572 26920 23624 26926
rect 23572 26862 23624 26868
rect 23296 26580 23348 26586
rect 23296 26522 23348 26528
rect 23204 26376 23256 26382
rect 23204 26318 23256 26324
rect 23216 26042 23244 26318
rect 23204 26036 23256 26042
rect 23204 25978 23256 25984
rect 23584 25770 23612 26862
rect 26240 26444 26292 26450
rect 26240 26386 26292 26392
rect 23572 25764 23624 25770
rect 23572 25706 23624 25712
rect 23112 25696 23164 25702
rect 23112 25638 23164 25644
rect 23124 25226 23152 25638
rect 23112 25220 23164 25226
rect 23112 25162 23164 25168
rect 23124 24954 23152 25162
rect 23112 24948 23164 24954
rect 23112 24890 23164 24896
rect 22928 23112 22980 23118
rect 22928 23054 22980 23060
rect 23584 22438 23612 25706
rect 24032 25220 24084 25226
rect 24032 25162 24084 25168
rect 24044 24342 24072 25162
rect 24032 24336 24084 24342
rect 24032 24278 24084 24284
rect 26252 23866 26280 26386
rect 26240 23860 26292 23866
rect 26240 23802 26292 23808
rect 23572 22432 23624 22438
rect 23572 22374 23624 22380
rect 22756 22066 22876 22094
rect 22756 19514 22784 22066
rect 26528 21486 26556 37062
rect 27620 36848 27672 36854
rect 27620 36790 27672 36796
rect 27632 35834 27660 36790
rect 28920 36650 28948 37198
rect 29012 37126 29040 39200
rect 30300 37330 30328 39200
rect 30288 37324 30340 37330
rect 30288 37266 30340 37272
rect 30656 37256 30708 37262
rect 30656 37198 30708 37204
rect 29000 37120 29052 37126
rect 29000 37062 29052 37068
rect 30668 36922 30696 37198
rect 31852 37188 31904 37194
rect 31852 37130 31904 37136
rect 31760 37120 31812 37126
rect 31760 37062 31812 37068
rect 30656 36916 30708 36922
rect 30656 36858 30708 36864
rect 31668 36780 31720 36786
rect 31668 36722 31720 36728
rect 28908 36644 28960 36650
rect 28908 36586 28960 36592
rect 27620 35828 27672 35834
rect 27620 35770 27672 35776
rect 31680 34066 31708 36722
rect 31668 34060 31720 34066
rect 31668 34002 31720 34008
rect 29828 26784 29880 26790
rect 29828 26726 29880 26732
rect 29840 26586 29868 26726
rect 29828 26580 29880 26586
rect 29828 26522 29880 26528
rect 30012 24744 30064 24750
rect 30012 24686 30064 24692
rect 27252 24200 27304 24206
rect 27252 24142 27304 24148
rect 27264 23866 27292 24142
rect 30024 23866 30052 24686
rect 27252 23860 27304 23866
rect 27252 23802 27304 23808
rect 30012 23860 30064 23866
rect 30012 23802 30064 23808
rect 31772 23186 31800 37062
rect 31864 36718 31892 37130
rect 32232 37126 32260 39200
rect 32404 37392 32456 37398
rect 32404 37334 32456 37340
rect 32220 37120 32272 37126
rect 32220 37062 32272 37068
rect 31852 36712 31904 36718
rect 31852 36654 31904 36660
rect 31760 23180 31812 23186
rect 31760 23122 31812 23128
rect 26516 21480 26568 21486
rect 26516 21422 26568 21428
rect 23296 19984 23348 19990
rect 23296 19926 23348 19932
rect 22744 19508 22796 19514
rect 22744 19450 22796 19456
rect 21824 12980 21876 12986
rect 21824 12922 21876 12928
rect 20260 9648 20312 9654
rect 20260 9590 20312 9596
rect 23308 2582 23336 19926
rect 24584 16652 24636 16658
rect 24584 16594 24636 16600
rect 24596 6914 24624 16594
rect 24952 11756 25004 11762
rect 24952 11698 25004 11704
rect 24964 11558 24992 11698
rect 24952 11552 25004 11558
rect 24952 11494 25004 11500
rect 24768 9376 24820 9382
rect 24768 9318 24820 9324
rect 24596 6886 24716 6914
rect 24688 6798 24716 6886
rect 24676 6792 24728 6798
rect 24676 6734 24728 6740
rect 24688 6662 24716 6734
rect 24676 6656 24728 6662
rect 24676 6598 24728 6604
rect 23296 2576 23348 2582
rect 23296 2518 23348 2524
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 12716 2440 12768 2446
rect 12716 2382 12768 2388
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 20076 2440 20128 2446
rect 20076 2382 20128 2388
rect 2412 2372 2464 2378
rect 2412 2314 2464 2320
rect 1674 1456 1730 1465
rect 1674 1391 1730 1400
rect 2424 1358 2452 2314
rect 3240 2304 3292 2310
rect 3240 2246 3292 2252
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 2412 1352 2464 1358
rect 2412 1294 2464 1300
rect 3252 800 3280 2246
rect 4540 800 4568 2246
rect 6472 800 6500 2246
rect 8404 800 8432 2246
rect 9692 800 9720 2382
rect 24780 2378 24808 9318
rect 24964 2514 24992 11494
rect 25228 6724 25280 6730
rect 25228 6666 25280 6672
rect 24952 2508 25004 2514
rect 24952 2450 25004 2456
rect 25240 2446 25268 6666
rect 27344 2916 27396 2922
rect 27344 2858 27396 2864
rect 27356 2446 27384 2858
rect 29644 2848 29696 2854
rect 29644 2790 29696 2796
rect 29656 2446 29684 2790
rect 32416 2650 32444 37334
rect 33520 37126 33548 39200
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 33600 37256 33652 37262
rect 33600 37198 33652 37204
rect 33508 37120 33560 37126
rect 33508 37062 33560 37068
rect 32956 25220 33008 25226
rect 32956 25162 33008 25168
rect 32968 6458 32996 25162
rect 33612 24410 33640 37198
rect 35452 37126 35480 39200
rect 36726 38856 36782 38865
rect 36726 38791 36782 38800
rect 36740 37466 36768 38791
rect 36728 37460 36780 37466
rect 36728 37402 36780 37408
rect 37384 37346 37412 39200
rect 38198 37496 38254 37505
rect 38198 37431 38254 37440
rect 37384 37318 37504 37346
rect 35532 37256 35584 37262
rect 35532 37198 35584 37204
rect 37372 37256 37424 37262
rect 37372 37198 37424 37204
rect 35440 37120 35492 37126
rect 35440 37062 35492 37068
rect 35544 36854 35572 37198
rect 35532 36848 35584 36854
rect 35532 36790 35584 36796
rect 34336 36780 34388 36786
rect 34336 36722 34388 36728
rect 34348 36242 34376 36722
rect 34428 36576 34480 36582
rect 34428 36518 34480 36524
rect 34336 36236 34388 36242
rect 34336 36178 34388 36184
rect 34440 36174 34468 36518
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34428 36168 34480 36174
rect 34428 36110 34480 36116
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34520 33380 34572 33386
rect 34520 33322 34572 33328
rect 34532 27402 34560 33322
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 36636 29028 36688 29034
rect 36636 28970 36688 28976
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34520 27396 34572 27402
rect 34520 27338 34572 27344
rect 36648 26994 36676 28970
rect 36636 26988 36688 26994
rect 36636 26930 36688 26936
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 36544 24608 36596 24614
rect 36544 24550 36596 24556
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 33600 24404 33652 24410
rect 33600 24346 33652 24352
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 36556 19854 36584 24550
rect 37384 21894 37412 37198
rect 37476 37126 37504 37318
rect 37464 37120 37516 37126
rect 37464 37062 37516 37068
rect 38212 36922 38240 37431
rect 38200 36916 38252 36922
rect 38200 36858 38252 36864
rect 38672 36378 38700 39200
rect 38660 36372 38712 36378
rect 38660 36314 38712 36320
rect 37464 35692 37516 35698
rect 37464 35634 37516 35640
rect 37476 35494 37504 35634
rect 37464 35488 37516 35494
rect 38200 35488 38252 35494
rect 37464 35430 37516 35436
rect 38198 35456 38200 35465
rect 38252 35456 38254 35465
rect 37372 21888 37424 21894
rect 37372 21830 37424 21836
rect 37476 19922 37504 35430
rect 38198 35391 38254 35400
rect 38200 33516 38252 33522
rect 38200 33458 38252 33464
rect 38212 33425 38240 33458
rect 38198 33416 38254 33425
rect 38198 33351 38254 33360
rect 38200 32428 38252 32434
rect 38200 32370 38252 32376
rect 38016 32292 38068 32298
rect 38016 32234 38068 32240
rect 37832 30184 37884 30190
rect 37832 30126 37884 30132
rect 37740 27940 37792 27946
rect 37740 27882 37792 27888
rect 37556 24064 37608 24070
rect 37556 24006 37608 24012
rect 37464 19916 37516 19922
rect 37464 19858 37516 19864
rect 36544 19848 36596 19854
rect 36544 19790 36596 19796
rect 33692 19780 33744 19786
rect 33692 19722 33744 19728
rect 32956 6452 33008 6458
rect 32956 6394 33008 6400
rect 33704 2650 33732 19722
rect 36728 19712 36780 19718
rect 36728 19654 36780 19660
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34796 16992 34848 16998
rect 34796 16934 34848 16940
rect 34520 6180 34572 6186
rect 34520 6122 34572 6128
rect 34532 3058 34560 6122
rect 34808 3194 34836 16934
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34796 3188 34848 3194
rect 34796 3130 34848 3136
rect 33876 3052 33928 3058
rect 33876 2994 33928 3000
rect 34520 3052 34572 3058
rect 34520 2994 34572 3000
rect 32404 2644 32456 2650
rect 32404 2586 32456 2592
rect 33692 2644 33744 2650
rect 33692 2586 33744 2592
rect 33888 2514 33916 2994
rect 33876 2508 33928 2514
rect 33876 2450 33928 2456
rect 34808 2446 34836 3130
rect 35900 2916 35952 2922
rect 35900 2858 35952 2864
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35912 2446 35940 2858
rect 36740 2650 36768 19654
rect 37464 12776 37516 12782
rect 37462 12744 37464 12753
rect 37516 12744 37518 12753
rect 37462 12679 37518 12688
rect 37464 3392 37516 3398
rect 37464 3334 37516 3340
rect 37476 2990 37504 3334
rect 37464 2984 37516 2990
rect 37464 2926 37516 2932
rect 36820 2848 36872 2854
rect 36820 2790 36872 2796
rect 36728 2644 36780 2650
rect 36728 2586 36780 2592
rect 25228 2440 25280 2446
rect 25228 2382 25280 2388
rect 27344 2440 27396 2446
rect 27344 2382 27396 2388
rect 29644 2440 29696 2446
rect 29644 2382 29696 2388
rect 34796 2440 34848 2446
rect 34796 2382 34848 2388
rect 35900 2440 35952 2446
rect 35900 2382 35952 2388
rect 11612 2372 11664 2378
rect 11612 2314 11664 2320
rect 14832 2372 14884 2378
rect 14832 2314 14884 2320
rect 18052 2372 18104 2378
rect 18052 2314 18104 2320
rect 23204 2372 23256 2378
rect 23204 2314 23256 2320
rect 24768 2372 24820 2378
rect 24768 2314 24820 2320
rect 11624 800 11652 2314
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 12912 800 12940 2246
rect 14844 800 14872 2314
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 16776 800 16804 2246
rect 18064 800 18092 2314
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 21640 2304 21692 2310
rect 21640 2246 21692 2252
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19996 800 20024 2246
rect 21284 870 21404 898
rect 21284 800 21312 870
rect 18 200 74 800
rect 1306 200 1362 800
rect 3238 200 3294 800
rect 4526 200 4582 800
rect 6458 200 6514 800
rect 8390 200 8446 800
rect 9678 200 9734 800
rect 11610 200 11666 800
rect 12898 200 12954 800
rect 14830 200 14886 800
rect 16762 200 16818 800
rect 18050 200 18106 800
rect 19982 200 20038 800
rect 21270 200 21326 800
rect 21376 762 21404 870
rect 21652 762 21680 2246
rect 23216 800 23244 2314
rect 25136 2304 25188 2310
rect 25136 2246 25188 2252
rect 26424 2304 26476 2310
rect 26424 2246 26476 2252
rect 28356 2304 28408 2310
rect 28356 2246 28408 2252
rect 25148 800 25176 2246
rect 26436 800 26464 2246
rect 28368 800 28396 2246
rect 29656 800 29684 2382
rect 36832 2378 36860 2790
rect 37568 2650 37596 24006
rect 37752 7478 37780 27882
rect 37844 25294 37872 30126
rect 38028 29510 38056 32234
rect 38212 32065 38240 32370
rect 38198 32056 38254 32065
rect 38198 31991 38254 32000
rect 38292 30184 38344 30190
rect 38292 30126 38344 30132
rect 38304 30025 38332 30126
rect 38290 30016 38346 30025
rect 38290 29951 38346 29960
rect 38304 29850 38332 29951
rect 38292 29844 38344 29850
rect 38292 29786 38344 29792
rect 38016 29504 38068 29510
rect 38016 29446 38068 29452
rect 38016 29096 38068 29102
rect 38016 29038 38068 29044
rect 38292 29096 38344 29102
rect 38292 29038 38344 29044
rect 38028 28490 38056 29038
rect 38304 28694 38332 29038
rect 38292 28688 38344 28694
rect 38290 28656 38292 28665
rect 38344 28656 38346 28665
rect 38290 28591 38346 28600
rect 38016 28484 38068 28490
rect 38016 28426 38068 28432
rect 38200 26784 38252 26790
rect 38200 26726 38252 26732
rect 38212 26625 38240 26726
rect 38198 26616 38254 26625
rect 38198 26551 38254 26560
rect 37924 26376 37976 26382
rect 37924 26318 37976 26324
rect 37832 25288 37884 25294
rect 37832 25230 37884 25236
rect 37844 24206 37872 25230
rect 37936 24750 37964 26318
rect 38292 25152 38344 25158
rect 38292 25094 38344 25100
rect 38304 24750 38332 25094
rect 37924 24744 37976 24750
rect 37924 24686 37976 24692
rect 38292 24744 38344 24750
rect 38292 24686 38344 24692
rect 37832 24200 37884 24206
rect 37832 24142 37884 24148
rect 37832 23724 37884 23730
rect 37832 23666 37884 23672
rect 37844 22438 37872 23666
rect 37832 22432 37884 22438
rect 37832 22374 37884 22380
rect 37844 22030 37872 22374
rect 37832 22024 37884 22030
rect 37832 21966 37884 21972
rect 37844 16574 37872 21966
rect 37936 20466 37964 24686
rect 38304 24585 38332 24686
rect 38290 24576 38346 24585
rect 38290 24511 38346 24520
rect 38016 24064 38068 24070
rect 38016 24006 38068 24012
rect 38028 23730 38056 24006
rect 38016 23724 38068 23730
rect 38016 23666 38068 23672
rect 38200 23520 38252 23526
rect 38200 23462 38252 23468
rect 38212 23225 38240 23462
rect 38198 23216 38254 23225
rect 38198 23151 38254 23160
rect 38016 22976 38068 22982
rect 38016 22918 38068 22924
rect 38028 21554 38056 22918
rect 38016 21548 38068 21554
rect 38016 21490 38068 21496
rect 38200 21344 38252 21350
rect 38200 21286 38252 21292
rect 38212 21185 38240 21286
rect 38198 21176 38254 21185
rect 38198 21111 38254 21120
rect 37924 20460 37976 20466
rect 37924 20402 37976 20408
rect 38108 20256 38160 20262
rect 38108 20198 38160 20204
rect 38016 17672 38068 17678
rect 38016 17614 38068 17620
rect 37844 16546 37964 16574
rect 37740 7472 37792 7478
rect 37740 7414 37792 7420
rect 37936 5846 37964 16546
rect 38028 14482 38056 17614
rect 38120 16114 38148 20198
rect 38198 19816 38254 19825
rect 38198 19751 38254 19760
rect 38212 19718 38240 19751
rect 38200 19712 38252 19718
rect 38200 19654 38252 19660
rect 38108 16108 38160 16114
rect 38108 16050 38160 16056
rect 38200 15904 38252 15910
rect 38200 15846 38252 15852
rect 38212 15745 38240 15846
rect 38198 15736 38254 15745
rect 38198 15671 38254 15680
rect 38016 14476 38068 14482
rect 38016 14418 38068 14424
rect 38028 12238 38056 14418
rect 38292 14408 38344 14414
rect 38290 14376 38292 14385
rect 38344 14376 38346 14385
rect 38290 14311 38346 14320
rect 38304 14074 38332 14311
rect 38292 14068 38344 14074
rect 38292 14010 38344 14016
rect 38200 12640 38252 12646
rect 38200 12582 38252 12588
rect 38212 12345 38240 12582
rect 38198 12336 38254 12345
rect 38198 12271 38254 12280
rect 38016 12232 38068 12238
rect 38016 12174 38068 12180
rect 38016 12096 38068 12102
rect 38016 12038 38068 12044
rect 38028 8974 38056 12038
rect 38108 11076 38160 11082
rect 38108 11018 38160 11024
rect 38200 11076 38252 11082
rect 38200 11018 38252 11024
rect 38016 8968 38068 8974
rect 38016 8910 38068 8916
rect 38120 6662 38148 11018
rect 38212 10985 38240 11018
rect 38198 10976 38254 10985
rect 38198 10911 38254 10920
rect 38198 8936 38254 8945
rect 38198 8871 38254 8880
rect 38212 8838 38240 8871
rect 38200 8832 38252 8838
rect 38200 8774 38252 8780
rect 38200 7404 38252 7410
rect 38200 7346 38252 7352
rect 38212 6905 38240 7346
rect 38198 6896 38254 6905
rect 38198 6831 38254 6840
rect 38108 6656 38160 6662
rect 38108 6598 38160 6604
rect 37924 5840 37976 5846
rect 37924 5782 37976 5788
rect 38200 5636 38252 5642
rect 38200 5578 38252 5584
rect 38212 5545 38240 5578
rect 38198 5536 38254 5545
rect 38198 5471 38254 5480
rect 38198 3496 38254 3505
rect 38198 3431 38254 3440
rect 38212 3398 38240 3431
rect 38200 3392 38252 3398
rect 38200 3334 38252 3340
rect 37648 2848 37700 2854
rect 37648 2790 37700 2796
rect 38016 2848 38068 2854
rect 38016 2790 38068 2796
rect 37556 2644 37608 2650
rect 37556 2586 37608 2592
rect 37280 2440 37332 2446
rect 37280 2382 37332 2388
rect 33508 2372 33560 2378
rect 33508 2314 33560 2320
rect 36820 2372 36872 2378
rect 36820 2314 36872 2320
rect 31760 2304 31812 2310
rect 31760 2246 31812 2252
rect 31772 1714 31800 2246
rect 31588 1686 31800 1714
rect 31588 800 31616 1686
rect 33520 800 33548 2314
rect 34796 2304 34848 2310
rect 34796 2246 34848 2252
rect 35808 2304 35860 2310
rect 37292 2292 37320 2382
rect 35808 2246 35860 2252
rect 37200 2264 37320 2292
rect 34808 800 34836 2246
rect 35820 2145 35848 2246
rect 35806 2136 35862 2145
rect 35806 2071 35862 2080
rect 36740 870 36860 898
rect 36740 800 36768 870
rect 21376 734 21680 762
rect 23202 200 23258 800
rect 25134 200 25190 800
rect 26422 200 26478 800
rect 28354 200 28410 800
rect 29642 200 29698 800
rect 31574 200 31630 800
rect 33506 200 33562 800
rect 34794 200 34850 800
rect 36726 200 36782 800
rect 36832 762 36860 870
rect 37200 762 37228 2264
rect 36832 734 37228 762
rect 37660 105 37688 2790
rect 38028 800 38056 2790
rect 38014 200 38070 800
rect 37646 96 37702 105
rect 37646 31 37702 40
<< via2 >>
rect 2410 38800 2466 38856
rect 1674 31320 1730 31376
rect 1582 30776 1638 30832
rect 1674 29960 1730 30016
rect 1766 27920 1822 27976
rect 1674 26560 1730 26616
rect 1582 24520 1638 24576
rect 1674 22500 1730 22536
rect 1674 22480 1676 22500
rect 1676 22480 1728 22500
rect 1728 22480 1730 22500
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 2870 36760 2926 36816
rect 2410 29552 2466 29608
rect 2686 33532 2688 33552
rect 2688 33532 2740 33552
rect 2740 33532 2742 33552
rect 2686 33496 2742 33532
rect 3238 33224 3294 33280
rect 3054 32408 3110 32464
rect 1674 21120 1730 21176
rect 1674 19116 1676 19136
rect 1676 19116 1728 19136
rect 1728 19116 1730 19136
rect 1674 19080 1730 19116
rect 1674 17720 1730 17776
rect 1674 15680 1730 15736
rect 1674 13676 1676 13696
rect 1676 13676 1728 13696
rect 1728 13676 1730 13696
rect 1674 13640 1730 13676
rect 1674 12280 1730 12336
rect 1674 10240 1730 10296
rect 1674 8900 1730 8936
rect 1674 8880 1676 8900
rect 1676 8880 1728 8900
rect 1728 8880 1730 8900
rect 3422 31764 3424 31784
rect 3424 31764 3476 31784
rect 3476 31764 3478 31784
rect 3422 31728 3478 31764
rect 3422 30368 3478 30424
rect 3606 29708 3662 29744
rect 3606 29688 3608 29708
rect 3608 29688 3660 29708
rect 3660 29688 3662 29708
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 3882 35672 3938 35728
rect 3790 35536 3846 35592
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4066 35012 4122 35048
rect 4066 34992 4068 35012
rect 4068 34992 4120 35012
rect 4120 34992 4122 35012
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4250 33768 4306 33824
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4066 33088 4122 33144
rect 4250 32272 4306 32328
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 5354 35692 5410 35728
rect 5354 35672 5356 35692
rect 5356 35672 5408 35692
rect 5408 35672 5410 35692
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4066 30676 4068 30696
rect 4068 30676 4120 30696
rect 4120 30676 4122 30696
rect 4066 30640 4122 30676
rect 4618 30096 4674 30152
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4710 28464 4766 28520
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4066 27548 4068 27568
rect 4068 27548 4120 27568
rect 4120 27548 4122 27568
rect 4066 27512 4122 27548
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 6734 36896 6790 36952
rect 5262 29008 5318 29064
rect 5354 28736 5410 28792
rect 5722 30368 5778 30424
rect 5906 30096 5962 30152
rect 5630 29300 5686 29336
rect 5630 29280 5632 29300
rect 5632 29280 5684 29300
rect 5684 29280 5686 29300
rect 6366 31592 6422 31648
rect 6274 29416 6330 29472
rect 6182 29280 6238 29336
rect 6182 29144 6238 29200
rect 6274 29028 6330 29064
rect 6274 29008 6276 29028
rect 6276 29008 6328 29028
rect 6328 29008 6330 29028
rect 6274 28872 6330 28928
rect 6826 34312 6882 34368
rect 7470 35400 7526 35456
rect 6642 30640 6698 30696
rect 6642 30096 6698 30152
rect 6642 29844 6698 29880
rect 6642 29824 6644 29844
rect 6644 29824 6696 29844
rect 6696 29824 6698 29844
rect 6642 29416 6698 29472
rect 6550 29144 6606 29200
rect 6734 29008 6790 29064
rect 6642 28464 6698 28520
rect 9034 36644 9090 36680
rect 9034 36624 9036 36644
rect 9036 36624 9088 36644
rect 9088 36624 9090 36644
rect 7746 34856 7802 34912
rect 7378 29280 7434 29336
rect 7838 33632 7894 33688
rect 7470 26696 7526 26752
rect 8206 34196 8262 34232
rect 8206 34176 8208 34196
rect 8208 34176 8260 34196
rect 8260 34176 8262 34196
rect 8206 33496 8262 33552
rect 8114 33088 8170 33144
rect 8022 32816 8078 32872
rect 8298 29552 8354 29608
rect 8022 29280 8078 29336
rect 8298 29280 8354 29336
rect 7930 29008 7986 29064
rect 8390 28464 8446 28520
rect 7286 24792 7342 24848
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 1582 6840 1638 6896
rect 1582 4820 1638 4856
rect 1582 4800 1584 4820
rect 1584 4800 1636 4820
rect 1636 4800 1638 4820
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 1674 3440 1730 3496
rect 8666 29824 8722 29880
rect 8390 23604 8392 23624
rect 8392 23604 8444 23624
rect 8444 23604 8446 23624
rect 8390 23568 8446 23604
rect 9034 29008 9090 29064
rect 9310 34040 9366 34096
rect 9310 32292 9366 32328
rect 9310 32272 9312 32292
rect 9312 32272 9364 32292
rect 9364 32272 9366 32292
rect 9310 29688 9366 29744
rect 9770 34584 9826 34640
rect 10966 37032 11022 37088
rect 10690 36080 10746 36136
rect 10782 35128 10838 35184
rect 10874 34584 10930 34640
rect 9586 32408 9642 32464
rect 9494 31900 9496 31920
rect 9496 31900 9548 31920
rect 9548 31900 9550 31920
rect 9494 31864 9550 31900
rect 9586 29416 9642 29472
rect 9862 33224 9918 33280
rect 9954 32716 9956 32736
rect 9956 32716 10008 32736
rect 10008 32716 10010 32736
rect 9954 32680 10010 32716
rect 10230 31456 10286 31512
rect 10138 31320 10194 31376
rect 9770 29416 9826 29472
rect 9770 29180 9772 29200
rect 9772 29180 9824 29200
rect 9824 29180 9826 29200
rect 9770 29144 9826 29180
rect 9402 28872 9458 28928
rect 9034 27920 9090 27976
rect 9218 28328 9274 28384
rect 10138 29824 10194 29880
rect 10414 29708 10470 29744
rect 10414 29688 10416 29708
rect 10416 29688 10468 29708
rect 10468 29688 10470 29708
rect 10414 29144 10470 29200
rect 10966 32680 11022 32736
rect 10874 31864 10930 31920
rect 10966 31728 11022 31784
rect 10874 30912 10930 30968
rect 10782 29688 10838 29744
rect 10046 28328 10102 28384
rect 8666 24520 8722 24576
rect 10046 27784 10102 27840
rect 10138 27668 10194 27704
rect 10138 27648 10140 27668
rect 10140 27648 10192 27668
rect 10192 27648 10194 27668
rect 10138 26832 10194 26888
rect 10230 26696 10286 26752
rect 10138 25064 10194 25120
rect 9678 23724 9734 23760
rect 9678 23704 9680 23724
rect 9680 23704 9732 23724
rect 9732 23704 9734 23724
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 10138 22072 10194 22128
rect 10414 29008 10470 29064
rect 10690 26832 10746 26888
rect 10322 25200 10378 25256
rect 10966 30252 11022 30288
rect 11242 36896 11298 36952
rect 11426 36624 11482 36680
rect 11334 35944 11390 36000
rect 11242 34856 11298 34912
rect 11334 33768 11390 33824
rect 11150 32564 11206 32600
rect 11150 32544 11152 32564
rect 11152 32544 11204 32564
rect 11204 32544 11206 32564
rect 10966 30232 10968 30252
rect 10968 30232 11020 30252
rect 11020 30232 11022 30252
rect 11518 32000 11574 32056
rect 11150 30096 11206 30152
rect 11518 30640 11574 30696
rect 11794 34040 11850 34096
rect 12898 37068 12900 37088
rect 12900 37068 12952 37088
rect 12952 37068 12954 37088
rect 12898 37032 12954 37068
rect 13450 37032 13506 37088
rect 12162 36216 12218 36272
rect 12530 36352 12586 36408
rect 13266 36216 13322 36272
rect 12714 35808 12770 35864
rect 12254 35284 12310 35320
rect 12254 35264 12256 35284
rect 12256 35264 12308 35284
rect 12308 35264 12310 35284
rect 13082 35264 13138 35320
rect 11886 32544 11942 32600
rect 12714 34740 12770 34776
rect 12714 34720 12716 34740
rect 12716 34720 12768 34740
rect 12768 34720 12770 34740
rect 12254 34448 12310 34504
rect 12346 34312 12402 34368
rect 12346 34196 12402 34232
rect 12346 34176 12348 34196
rect 12348 34176 12400 34196
rect 12400 34176 12402 34196
rect 12806 34584 12862 34640
rect 12530 34176 12586 34232
rect 12622 33496 12678 33552
rect 12898 33496 12954 33552
rect 12254 32272 12310 32328
rect 12254 31864 12310 31920
rect 12162 31320 12218 31376
rect 11334 29960 11390 30016
rect 11242 29552 11298 29608
rect 11150 28600 11206 28656
rect 11518 29280 11574 29336
rect 11058 25744 11114 25800
rect 10966 23860 11022 23896
rect 10966 23840 10968 23860
rect 10968 23840 11020 23860
rect 11020 23840 11022 23860
rect 11058 23568 11114 23624
rect 11610 28736 11666 28792
rect 11702 28464 11758 28520
rect 11794 28328 11850 28384
rect 11978 29280 12034 29336
rect 12346 30912 12402 30968
rect 12346 28056 12402 28112
rect 12254 27648 12310 27704
rect 12254 25100 12256 25120
rect 12256 25100 12308 25120
rect 12308 25100 12310 25120
rect 11978 23724 12034 23760
rect 11978 23704 11980 23724
rect 11980 23704 12032 23724
rect 12032 23704 12034 23724
rect 11886 23588 11942 23624
rect 11886 23568 11888 23588
rect 11888 23568 11940 23588
rect 11940 23568 11942 23588
rect 11702 22072 11758 22128
rect 12254 25064 12310 25100
rect 12254 22072 12310 22128
rect 12622 32272 12678 32328
rect 12622 31864 12678 31920
rect 12622 31728 12678 31784
rect 13174 32444 13176 32464
rect 13176 32444 13228 32464
rect 13228 32444 13230 32464
rect 13174 32408 13230 32444
rect 14002 35400 14058 35456
rect 14186 35400 14242 35456
rect 13818 34448 13874 34504
rect 13726 33632 13782 33688
rect 14002 34584 14058 34640
rect 13910 33768 13966 33824
rect 13818 32544 13874 32600
rect 12806 32136 12862 32192
rect 12714 29960 12770 30016
rect 12530 28328 12586 28384
rect 12530 28056 12586 28112
rect 12530 26832 12586 26888
rect 12438 26424 12494 26480
rect 12806 29824 12862 29880
rect 13082 31320 13138 31376
rect 12806 28056 12862 28112
rect 12530 26016 12586 26072
rect 12714 23840 12770 23896
rect 12622 23568 12678 23624
rect 13358 24656 13414 24712
rect 13634 28600 13690 28656
rect 13450 23160 13506 23216
rect 14002 30912 14058 30968
rect 14002 30388 14058 30424
rect 14002 30368 14004 30388
rect 14004 30368 14056 30388
rect 14056 30368 14058 30388
rect 14094 28872 14150 28928
rect 14646 34856 14702 34912
rect 14370 34076 14372 34096
rect 14372 34076 14424 34096
rect 14424 34076 14426 34096
rect 14370 34040 14426 34076
rect 14278 30096 14334 30152
rect 14278 29688 14334 29744
rect 14646 32000 14702 32056
rect 15198 35128 15254 35184
rect 15198 32952 15254 33008
rect 15474 35692 15530 35728
rect 15474 35672 15476 35692
rect 15476 35672 15528 35692
rect 15528 35672 15530 35692
rect 14922 31628 14924 31648
rect 14924 31628 14976 31648
rect 14976 31628 14978 31648
rect 14922 31592 14978 31628
rect 15106 31764 15108 31784
rect 15108 31764 15160 31784
rect 15160 31764 15162 31784
rect 15106 31728 15162 31764
rect 14278 29008 14334 29064
rect 14186 28192 14242 28248
rect 15934 36352 15990 36408
rect 15842 35944 15898 36000
rect 15658 34040 15714 34096
rect 15474 32000 15530 32056
rect 15842 32000 15898 32056
rect 16118 34720 16174 34776
rect 14462 26696 14518 26752
rect 14370 25744 14426 25800
rect 14278 25236 14280 25256
rect 14280 25236 14332 25256
rect 14332 25236 14334 25256
rect 14278 25200 14334 25236
rect 14002 23704 14058 23760
rect 12714 10260 12770 10296
rect 12714 10240 12716 10260
rect 12716 10240 12768 10260
rect 12768 10240 12770 10260
rect 11886 2644 11942 2680
rect 11886 2624 11888 2644
rect 11888 2624 11940 2644
rect 11940 2624 11942 2644
rect 15658 29688 15714 29744
rect 15658 24812 15714 24848
rect 15658 24792 15660 24812
rect 15660 24792 15712 24812
rect 15712 24792 15714 24812
rect 18602 37032 18658 37088
rect 16670 33224 16726 33280
rect 16670 31320 16726 31376
rect 16670 30676 16672 30696
rect 16672 30676 16724 30696
rect 16724 30676 16726 30696
rect 16670 30640 16726 30676
rect 16946 35708 16948 35728
rect 16948 35708 17000 35728
rect 17000 35708 17002 35728
rect 16946 35672 17002 35708
rect 17038 34892 17040 34912
rect 17040 34892 17092 34912
rect 17092 34892 17094 34912
rect 17038 34856 17094 34892
rect 17406 33652 17462 33688
rect 17406 33632 17408 33652
rect 17408 33632 17460 33652
rect 17460 33632 17462 33652
rect 17958 35828 18014 35864
rect 17958 35808 17960 35828
rect 17960 35808 18012 35828
rect 18012 35808 18014 35828
rect 17958 35264 18014 35320
rect 18694 36080 18750 36136
rect 17314 32680 17370 32736
rect 17406 32272 17462 32328
rect 16946 31592 17002 31648
rect 17958 34604 18014 34640
rect 17958 34584 17960 34604
rect 17960 34584 18012 34604
rect 18012 34584 18014 34604
rect 18510 35400 18566 35456
rect 17406 30912 17462 30968
rect 16394 29824 16450 29880
rect 16118 28056 16174 28112
rect 16670 28736 16726 28792
rect 16210 26424 16266 26480
rect 16854 27784 16910 27840
rect 16946 26016 17002 26072
rect 15658 21936 15714 21992
rect 16394 21936 16450 21992
rect 17130 28872 17186 28928
rect 17314 30368 17370 30424
rect 17406 28872 17462 28928
rect 18510 33496 18566 33552
rect 18786 34992 18842 35048
rect 18142 32408 18198 32464
rect 17958 31728 18014 31784
rect 18050 29708 18106 29744
rect 18050 29688 18052 29708
rect 18052 29688 18104 29708
rect 18104 29688 18106 29708
rect 17682 26424 17738 26480
rect 17682 24656 17738 24712
rect 17590 24556 17592 24576
rect 17592 24556 17644 24576
rect 17644 24556 17646 24576
rect 17590 24520 17646 24556
rect 17958 26016 18014 26072
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19522 34992 19578 35048
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19522 34176 19578 34232
rect 19430 33904 19486 33960
rect 19890 34060 19946 34096
rect 19890 34040 19892 34060
rect 19892 34040 19944 34060
rect 19944 34040 19946 34060
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19246 32544 19302 32600
rect 19062 32136 19118 32192
rect 18418 30776 18474 30832
rect 18878 30640 18934 30696
rect 19614 33260 19616 33280
rect 19616 33260 19668 33280
rect 19668 33260 19670 33280
rect 19614 33224 19670 33260
rect 20166 33108 20222 33144
rect 20166 33088 20168 33108
rect 20168 33088 20220 33108
rect 20220 33088 20222 33108
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19430 31728 19486 31784
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19430 31456 19486 31512
rect 18602 28600 18658 28656
rect 18418 26696 18474 26752
rect 18050 22772 18106 22808
rect 18050 22752 18052 22772
rect 18052 22752 18104 22772
rect 18104 22752 18106 22772
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19614 29144 19670 29200
rect 20074 30504 20130 30560
rect 20350 30504 20406 30560
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19706 26968 19762 27024
rect 19338 26324 19340 26344
rect 19340 26324 19392 26344
rect 19392 26324 19394 26344
rect 19338 26288 19394 26324
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 20258 29280 20314 29336
rect 20626 34060 20682 34096
rect 20626 34040 20628 34060
rect 20628 34040 20680 34060
rect 20680 34040 20682 34060
rect 20534 31728 20590 31784
rect 20442 29280 20498 29336
rect 21086 32836 21142 32872
rect 21086 32816 21088 32836
rect 21088 32816 21140 32836
rect 21140 32816 21142 32836
rect 21362 30912 21418 30968
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 20902 26324 20904 26344
rect 20904 26324 20956 26344
rect 20956 26324 20958 26344
rect 20902 26288 20958 26324
rect 23662 33380 23718 33416
rect 23662 33360 23664 33380
rect 23664 33360 23716 33380
rect 23716 33360 23718 33380
rect 23386 26968 23442 27024
rect 25318 35572 25320 35592
rect 25320 35572 25372 35592
rect 25372 35572 25374 35592
rect 25318 35536 25374 35572
rect 1674 1400 1730 1456
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 36726 38800 36782 38856
rect 38198 37440 38254 37496
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 38198 35436 38200 35456
rect 38200 35436 38252 35456
rect 38252 35436 38254 35456
rect 38198 35400 38254 35436
rect 38198 33360 38254 33416
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 37462 12724 37464 12744
rect 37464 12724 37516 12744
rect 37516 12724 37518 12744
rect 37462 12688 37518 12724
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 38198 32000 38254 32056
rect 38290 29960 38346 30016
rect 38290 28636 38292 28656
rect 38292 28636 38344 28656
rect 38344 28636 38346 28656
rect 38290 28600 38346 28636
rect 38198 26560 38254 26616
rect 38290 24520 38346 24576
rect 38198 23160 38254 23216
rect 38198 21120 38254 21176
rect 38198 19760 38254 19816
rect 38198 15680 38254 15736
rect 38290 14356 38292 14376
rect 38292 14356 38344 14376
rect 38344 14356 38346 14376
rect 38290 14320 38346 14356
rect 38198 12280 38254 12336
rect 38198 10920 38254 10976
rect 38198 8880 38254 8936
rect 38198 6840 38254 6896
rect 38198 5480 38254 5536
rect 38198 3440 38254 3496
rect 35806 2080 35862 2136
rect 37646 40 37702 96
<< metal3 >>
rect 200 38858 800 38888
rect 2405 38858 2471 38861
rect 200 38856 2471 38858
rect 200 38800 2410 38856
rect 2466 38800 2471 38856
rect 200 38798 2471 38800
rect 200 38768 800 38798
rect 2405 38795 2471 38798
rect 36721 38858 36787 38861
rect 39200 38858 39800 38888
rect 36721 38856 39800 38858
rect 36721 38800 36726 38856
rect 36782 38800 39800 38856
rect 36721 38798 39800 38800
rect 36721 38795 36787 38798
rect 39200 38768 39800 38798
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 38193 37498 38259 37501
rect 39200 37498 39800 37528
rect 38193 37496 39800 37498
rect 38193 37440 38198 37496
rect 38254 37440 39800 37496
rect 38193 37438 39800 37440
rect 38193 37435 38259 37438
rect 39200 37408 39800 37438
rect 10961 37090 11027 37093
rect 12893 37090 12959 37093
rect 10961 37088 12959 37090
rect 10961 37032 10966 37088
rect 11022 37032 12898 37088
rect 12954 37032 12959 37088
rect 10961 37030 12959 37032
rect 10961 37027 11027 37030
rect 12893 37027 12959 37030
rect 13445 37090 13511 37093
rect 18597 37090 18663 37093
rect 13445 37088 18663 37090
rect 13445 37032 13450 37088
rect 13506 37032 18602 37088
rect 18658 37032 18663 37088
rect 13445 37030 18663 37032
rect 13445 37027 13511 37030
rect 18597 37027 18663 37030
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 6729 36954 6795 36957
rect 11237 36954 11303 36957
rect 6729 36952 11303 36954
rect 6729 36896 6734 36952
rect 6790 36896 11242 36952
rect 11298 36896 11303 36952
rect 6729 36894 11303 36896
rect 6729 36891 6795 36894
rect 11237 36891 11303 36894
rect 200 36818 800 36848
rect 2865 36818 2931 36821
rect 200 36816 2931 36818
rect 200 36760 2870 36816
rect 2926 36760 2931 36816
rect 200 36758 2931 36760
rect 200 36728 800 36758
rect 2865 36755 2931 36758
rect 9029 36682 9095 36685
rect 11421 36682 11487 36685
rect 9029 36680 11487 36682
rect 9029 36624 9034 36680
rect 9090 36624 11426 36680
rect 11482 36624 11487 36680
rect 9029 36622 11487 36624
rect 9029 36619 9095 36622
rect 11421 36619 11487 36622
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 12525 36410 12591 36413
rect 15929 36410 15995 36413
rect 12525 36408 15995 36410
rect 12525 36352 12530 36408
rect 12586 36352 15934 36408
rect 15990 36352 15995 36408
rect 12525 36350 15995 36352
rect 12525 36347 12591 36350
rect 15929 36347 15995 36350
rect 12157 36274 12223 36277
rect 13261 36274 13327 36277
rect 12157 36272 13327 36274
rect 12157 36216 12162 36272
rect 12218 36216 13266 36272
rect 13322 36216 13327 36272
rect 12157 36214 13327 36216
rect 12157 36211 12223 36214
rect 13261 36211 13327 36214
rect 10685 36138 10751 36141
rect 18689 36138 18755 36141
rect 10685 36136 18755 36138
rect 10685 36080 10690 36136
rect 10746 36080 18694 36136
rect 18750 36080 18755 36136
rect 10685 36078 18755 36080
rect 10685 36075 10751 36078
rect 18689 36075 18755 36078
rect 11329 36004 11395 36005
rect 11278 36002 11284 36004
rect 11238 35942 11284 36002
rect 11348 36000 11395 36004
rect 11390 35944 11395 36000
rect 11278 35940 11284 35942
rect 11348 35940 11395 35944
rect 11329 35939 11395 35940
rect 15837 36004 15903 36005
rect 15837 36000 15884 36004
rect 15948 36002 15954 36004
rect 15837 35944 15842 36000
rect 15837 35940 15884 35944
rect 15948 35942 15994 36002
rect 15948 35940 15954 35942
rect 15837 35939 15903 35940
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 12709 35866 12775 35869
rect 17953 35866 18019 35869
rect 12709 35864 18019 35866
rect 12709 35808 12714 35864
rect 12770 35808 17958 35864
rect 18014 35808 18019 35864
rect 12709 35806 18019 35808
rect 12709 35803 12775 35806
rect 17953 35803 18019 35806
rect 3877 35730 3943 35733
rect 5349 35730 5415 35733
rect 3877 35728 5415 35730
rect 3877 35672 3882 35728
rect 3938 35672 5354 35728
rect 5410 35672 5415 35728
rect 3877 35670 5415 35672
rect 3877 35667 3943 35670
rect 5349 35667 5415 35670
rect 15142 35668 15148 35732
rect 15212 35730 15218 35732
rect 15469 35730 15535 35733
rect 16941 35730 17007 35733
rect 15212 35728 17007 35730
rect 15212 35672 15474 35728
rect 15530 35672 16946 35728
rect 17002 35672 17007 35728
rect 15212 35670 17007 35672
rect 15212 35668 15218 35670
rect 15469 35667 15535 35670
rect 16941 35667 17007 35670
rect 3785 35594 3851 35597
rect 25313 35594 25379 35597
rect 3785 35592 25379 35594
rect 3785 35536 3790 35592
rect 3846 35536 25318 35592
rect 25374 35536 25379 35592
rect 3785 35534 25379 35536
rect 3785 35531 3851 35534
rect 25313 35531 25379 35534
rect 200 35368 800 35488
rect 7465 35458 7531 35461
rect 13997 35458 14063 35461
rect 7465 35456 14063 35458
rect 7465 35400 7470 35456
rect 7526 35400 14002 35456
rect 14058 35400 14063 35456
rect 7465 35398 14063 35400
rect 7465 35395 7531 35398
rect 13997 35395 14063 35398
rect 14181 35458 14247 35461
rect 18505 35458 18571 35461
rect 14181 35456 18571 35458
rect 14181 35400 14186 35456
rect 14242 35400 18510 35456
rect 18566 35400 18571 35456
rect 14181 35398 18571 35400
rect 14181 35395 14247 35398
rect 18505 35395 18571 35398
rect 38193 35458 38259 35461
rect 39200 35458 39800 35488
rect 38193 35456 39800 35458
rect 38193 35400 38198 35456
rect 38254 35400 39800 35456
rect 38193 35398 39800 35400
rect 38193 35395 38259 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 39200 35368 39800 35398
rect 34930 35327 35246 35328
rect 12249 35322 12315 35325
rect 13077 35322 13143 35325
rect 17953 35322 18019 35325
rect 12249 35320 18019 35322
rect 12249 35264 12254 35320
rect 12310 35264 13082 35320
rect 13138 35264 17958 35320
rect 18014 35264 18019 35320
rect 12249 35262 18019 35264
rect 12249 35259 12315 35262
rect 13077 35259 13143 35262
rect 17953 35259 18019 35262
rect 10777 35186 10843 35189
rect 15193 35186 15259 35189
rect 10777 35184 15259 35186
rect 10777 35128 10782 35184
rect 10838 35128 15198 35184
rect 15254 35128 15259 35184
rect 10777 35126 15259 35128
rect 10777 35123 10843 35126
rect 15193 35123 15259 35126
rect 4061 35050 4127 35053
rect 18781 35050 18847 35053
rect 4061 35048 18847 35050
rect 4061 34992 4066 35048
rect 4122 34992 18786 35048
rect 18842 34992 18847 35048
rect 4061 34990 18847 34992
rect 4061 34987 4127 34990
rect 18781 34987 18847 34990
rect 19374 34988 19380 35052
rect 19444 35050 19450 35052
rect 19517 35050 19583 35053
rect 19444 35048 19583 35050
rect 19444 34992 19522 35048
rect 19578 34992 19583 35048
rect 19444 34990 19583 34992
rect 19444 34988 19450 34990
rect 19517 34987 19583 34990
rect 7741 34914 7807 34917
rect 11237 34914 11303 34917
rect 7741 34912 11303 34914
rect 7741 34856 7746 34912
rect 7802 34856 11242 34912
rect 11298 34856 11303 34912
rect 7741 34854 11303 34856
rect 7741 34851 7807 34854
rect 11237 34851 11303 34854
rect 14641 34914 14707 34917
rect 17033 34914 17099 34917
rect 14641 34912 17099 34914
rect 14641 34856 14646 34912
rect 14702 34856 17038 34912
rect 17094 34856 17099 34912
rect 14641 34854 17099 34856
rect 14641 34851 14707 34854
rect 17033 34851 17099 34854
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 12709 34778 12775 34781
rect 16113 34778 16179 34781
rect 12709 34776 16179 34778
rect 12709 34720 12714 34776
rect 12770 34720 16118 34776
rect 16174 34720 16179 34776
rect 12709 34718 16179 34720
rect 12709 34715 12775 34718
rect 16113 34715 16179 34718
rect 9622 34580 9628 34644
rect 9692 34642 9698 34644
rect 9765 34642 9831 34645
rect 9692 34640 9831 34642
rect 9692 34584 9770 34640
rect 9826 34584 9831 34640
rect 9692 34582 9831 34584
rect 9692 34580 9698 34582
rect 9765 34579 9831 34582
rect 10869 34642 10935 34645
rect 12801 34642 12867 34645
rect 10869 34640 12867 34642
rect 10869 34584 10874 34640
rect 10930 34584 12806 34640
rect 12862 34584 12867 34640
rect 10869 34582 12867 34584
rect 10869 34579 10935 34582
rect 12801 34579 12867 34582
rect 13997 34642 14063 34645
rect 17953 34642 18019 34645
rect 13997 34640 18019 34642
rect 13997 34584 14002 34640
rect 14058 34584 17958 34640
rect 18014 34584 18019 34640
rect 13997 34582 18019 34584
rect 13997 34579 14063 34582
rect 17953 34579 18019 34582
rect 12249 34506 12315 34509
rect 13813 34506 13879 34509
rect 12249 34504 13879 34506
rect 12249 34448 12254 34504
rect 12310 34448 13818 34504
rect 13874 34448 13879 34504
rect 12249 34446 13879 34448
rect 12249 34443 12315 34446
rect 13813 34443 13879 34446
rect 6821 34370 6887 34373
rect 12341 34370 12407 34373
rect 6821 34368 12407 34370
rect 6821 34312 6826 34368
rect 6882 34312 12346 34368
rect 12402 34312 12407 34368
rect 6821 34310 12407 34312
rect 6821 34307 6887 34310
rect 12341 34307 12407 34310
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 8201 34234 8267 34237
rect 12341 34234 12407 34237
rect 8201 34232 12407 34234
rect 8201 34176 8206 34232
rect 8262 34176 12346 34232
rect 12402 34176 12407 34232
rect 8201 34174 12407 34176
rect 8201 34171 8267 34174
rect 12341 34171 12407 34174
rect 12525 34234 12591 34237
rect 19517 34234 19583 34237
rect 12525 34232 19583 34234
rect 12525 34176 12530 34232
rect 12586 34176 19522 34232
rect 19578 34176 19583 34232
rect 12525 34174 19583 34176
rect 12525 34171 12591 34174
rect 19517 34171 19583 34174
rect 9305 34098 9371 34101
rect 11789 34098 11855 34101
rect 9305 34096 11855 34098
rect 9305 34040 9310 34096
rect 9366 34040 11794 34096
rect 11850 34040 11855 34096
rect 9305 34038 11855 34040
rect 9305 34035 9371 34038
rect 11789 34035 11855 34038
rect 14365 34098 14431 34101
rect 15653 34098 15719 34101
rect 14365 34096 15719 34098
rect 14365 34040 14370 34096
rect 14426 34040 15658 34096
rect 15714 34040 15719 34096
rect 14365 34038 15719 34040
rect 14365 34035 14431 34038
rect 15653 34035 15719 34038
rect 19885 34098 19951 34101
rect 20621 34098 20687 34101
rect 19885 34096 20687 34098
rect 19885 34040 19890 34096
rect 19946 34040 20626 34096
rect 20682 34040 20687 34096
rect 19885 34038 20687 34040
rect 19885 34035 19951 34038
rect 20621 34035 20687 34038
rect 19425 33962 19491 33965
rect 2730 33960 19491 33962
rect 2730 33904 19430 33960
rect 19486 33904 19491 33960
rect 2730 33902 19491 33904
rect 2730 33557 2790 33902
rect 19425 33899 19491 33902
rect 3550 33764 3556 33828
rect 3620 33826 3626 33828
rect 4245 33826 4311 33829
rect 3620 33824 4311 33826
rect 3620 33768 4250 33824
rect 4306 33768 4311 33824
rect 3620 33766 4311 33768
rect 3620 33764 3626 33766
rect 4245 33763 4311 33766
rect 11329 33826 11395 33829
rect 13905 33826 13971 33829
rect 11329 33824 13971 33826
rect 11329 33768 11334 33824
rect 11390 33768 13910 33824
rect 13966 33768 13971 33824
rect 11329 33766 13971 33768
rect 11329 33763 11395 33766
rect 13905 33763 13971 33766
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 7833 33690 7899 33693
rect 13721 33690 13787 33693
rect 17401 33690 17467 33693
rect 7833 33688 17467 33690
rect 7833 33632 7838 33688
rect 7894 33632 13726 33688
rect 13782 33632 17406 33688
rect 17462 33632 17467 33688
rect 7833 33630 17467 33632
rect 7833 33627 7899 33630
rect 13721 33627 13787 33630
rect 17401 33627 17467 33630
rect 2681 33552 2790 33557
rect 2681 33496 2686 33552
rect 2742 33496 2790 33552
rect 2681 33494 2790 33496
rect 8201 33554 8267 33557
rect 12617 33554 12683 33557
rect 8201 33552 12683 33554
rect 8201 33496 8206 33552
rect 8262 33496 12622 33552
rect 12678 33496 12683 33552
rect 8201 33494 12683 33496
rect 2681 33491 2747 33494
rect 8201 33491 8267 33494
rect 12617 33491 12683 33494
rect 12893 33554 12959 33557
rect 18505 33554 18571 33557
rect 12893 33552 18571 33554
rect 12893 33496 12898 33552
rect 12954 33496 18510 33552
rect 18566 33496 18571 33552
rect 12893 33494 18571 33496
rect 12893 33491 12959 33494
rect 18505 33491 18571 33494
rect 200 33418 800 33448
rect 23657 33418 23723 33421
rect 200 33416 23723 33418
rect 200 33360 23662 33416
rect 23718 33360 23723 33416
rect 200 33358 23723 33360
rect 200 33328 800 33358
rect 3233 33282 3299 33285
rect 3734 33282 3740 33284
rect 3233 33280 3740 33282
rect 3233 33224 3238 33280
rect 3294 33224 3740 33280
rect 3233 33222 3740 33224
rect 3233 33219 3299 33222
rect 3734 33220 3740 33222
rect 3804 33220 3810 33284
rect 3926 33146 3986 33358
rect 23657 33355 23723 33358
rect 38193 33418 38259 33421
rect 39200 33418 39800 33448
rect 38193 33416 39800 33418
rect 38193 33360 38198 33416
rect 38254 33360 39800 33416
rect 38193 33358 39800 33360
rect 38193 33355 38259 33358
rect 39200 33328 39800 33358
rect 9857 33284 9923 33285
rect 9806 33282 9812 33284
rect 9766 33222 9812 33282
rect 9876 33280 9923 33284
rect 9918 33224 9923 33280
rect 9806 33220 9812 33222
rect 9876 33220 9923 33224
rect 9857 33219 9923 33220
rect 16665 33282 16731 33285
rect 19609 33282 19675 33285
rect 16665 33280 19675 33282
rect 16665 33224 16670 33280
rect 16726 33224 19614 33280
rect 19670 33224 19675 33280
rect 16665 33222 19675 33224
rect 16665 33219 16731 33222
rect 19609 33219 19675 33222
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 4061 33146 4127 33149
rect 3926 33144 4127 33146
rect 3926 33088 4066 33144
rect 4122 33088 4127 33144
rect 3926 33086 4127 33088
rect 4061 33083 4127 33086
rect 8109 33146 8175 33149
rect 20161 33146 20227 33149
rect 8109 33144 20227 33146
rect 8109 33088 8114 33144
rect 8170 33088 20166 33144
rect 20222 33088 20227 33144
rect 8109 33086 20227 33088
rect 8109 33083 8175 33086
rect 20161 33083 20227 33086
rect 15193 33010 15259 33013
rect 15694 33010 15700 33012
rect 15193 33008 15700 33010
rect 15193 32952 15198 33008
rect 15254 32952 15700 33008
rect 15193 32950 15700 32952
rect 15193 32947 15259 32950
rect 15694 32948 15700 32950
rect 15764 32948 15770 33012
rect 8017 32874 8083 32877
rect 21081 32874 21147 32877
rect 8017 32872 21147 32874
rect 8017 32816 8022 32872
rect 8078 32816 21086 32872
rect 21142 32816 21147 32872
rect 8017 32814 21147 32816
rect 8017 32811 8083 32814
rect 21081 32811 21147 32814
rect 9949 32738 10015 32741
rect 10542 32738 10548 32740
rect 9949 32736 10548 32738
rect 9949 32680 9954 32736
rect 10010 32680 10548 32736
rect 9949 32678 10548 32680
rect 9949 32675 10015 32678
rect 10542 32676 10548 32678
rect 10612 32676 10618 32740
rect 10961 32738 11027 32741
rect 17309 32738 17375 32741
rect 10961 32736 17375 32738
rect 10961 32680 10966 32736
rect 11022 32680 17314 32736
rect 17370 32680 17375 32736
rect 10961 32678 17375 32680
rect 10961 32675 11027 32678
rect 17309 32675 17375 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 11145 32602 11211 32605
rect 11881 32602 11947 32605
rect 11145 32600 11947 32602
rect 11145 32544 11150 32600
rect 11206 32544 11886 32600
rect 11942 32544 11947 32600
rect 11145 32542 11947 32544
rect 11145 32539 11211 32542
rect 11881 32539 11947 32542
rect 13813 32602 13879 32605
rect 19241 32602 19307 32605
rect 13813 32600 19307 32602
rect 13813 32544 13818 32600
rect 13874 32544 19246 32600
rect 19302 32544 19307 32600
rect 13813 32542 19307 32544
rect 13813 32539 13879 32542
rect 19241 32539 19307 32542
rect 3049 32466 3115 32469
rect 9581 32466 9647 32469
rect 3049 32464 9647 32466
rect 3049 32408 3054 32464
rect 3110 32408 9586 32464
rect 9642 32408 9647 32464
rect 3049 32406 9647 32408
rect 3049 32403 3115 32406
rect 9581 32403 9647 32406
rect 13169 32466 13235 32469
rect 18137 32466 18203 32469
rect 13169 32464 18203 32466
rect 13169 32408 13174 32464
rect 13230 32408 18142 32464
rect 18198 32408 18203 32464
rect 13169 32406 18203 32408
rect 13169 32403 13235 32406
rect 18137 32403 18203 32406
rect 4245 32330 4311 32333
rect 4838 32330 4844 32332
rect 4245 32328 4844 32330
rect 4245 32272 4250 32328
rect 4306 32272 4844 32328
rect 4245 32270 4844 32272
rect 4245 32267 4311 32270
rect 4838 32268 4844 32270
rect 4908 32268 4914 32332
rect 9305 32330 9371 32333
rect 12249 32330 12315 32333
rect 9305 32328 12315 32330
rect 9305 32272 9310 32328
rect 9366 32272 12254 32328
rect 12310 32272 12315 32328
rect 9305 32270 12315 32272
rect 9305 32267 9371 32270
rect 12249 32267 12315 32270
rect 12617 32330 12683 32333
rect 17401 32330 17467 32333
rect 12617 32328 17467 32330
rect 12617 32272 12622 32328
rect 12678 32272 17406 32328
rect 17462 32272 17467 32328
rect 12617 32270 17467 32272
rect 12617 32267 12683 32270
rect 17401 32267 17467 32270
rect 12801 32194 12867 32197
rect 19057 32194 19123 32197
rect 12801 32192 19123 32194
rect 12801 32136 12806 32192
rect 12862 32136 19062 32192
rect 19118 32136 19123 32192
rect 12801 32134 19123 32136
rect 12801 32131 12867 32134
rect 19057 32131 19123 32134
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 11513 32058 11579 32061
rect 14641 32058 14707 32061
rect 11513 32056 14707 32058
rect 11513 32000 11518 32056
rect 11574 32000 14646 32056
rect 14702 32000 14707 32056
rect 11513 31998 14707 32000
rect 11513 31995 11579 31998
rect 14641 31995 14707 31998
rect 15469 32058 15535 32061
rect 15837 32058 15903 32061
rect 15469 32056 15903 32058
rect 15469 32000 15474 32056
rect 15530 32000 15842 32056
rect 15898 32000 15903 32056
rect 15469 31998 15903 32000
rect 15469 31995 15535 31998
rect 15837 31995 15903 31998
rect 38193 32058 38259 32061
rect 39200 32058 39800 32088
rect 38193 32056 39800 32058
rect 38193 32000 38198 32056
rect 38254 32000 39800 32056
rect 38193 31998 39800 32000
rect 38193 31995 38259 31998
rect 39200 31968 39800 31998
rect 9489 31922 9555 31925
rect 10869 31922 10935 31925
rect 9489 31920 10935 31922
rect 9489 31864 9494 31920
rect 9550 31864 10874 31920
rect 10930 31864 10935 31920
rect 9489 31862 10935 31864
rect 9489 31859 9555 31862
rect 10869 31859 10935 31862
rect 12249 31922 12315 31925
rect 12617 31922 12683 31925
rect 12249 31920 12683 31922
rect 12249 31864 12254 31920
rect 12310 31864 12622 31920
rect 12678 31864 12683 31920
rect 12249 31862 12683 31864
rect 12249 31859 12315 31862
rect 12617 31859 12683 31862
rect 3417 31786 3483 31789
rect 3918 31786 3924 31788
rect 3417 31784 3924 31786
rect 3417 31728 3422 31784
rect 3478 31728 3924 31784
rect 3417 31726 3924 31728
rect 3417 31723 3483 31726
rect 3918 31724 3924 31726
rect 3988 31724 3994 31788
rect 10961 31786 11027 31789
rect 12617 31786 12683 31789
rect 10961 31784 12683 31786
rect 10961 31728 10966 31784
rect 11022 31728 12622 31784
rect 12678 31728 12683 31784
rect 10961 31726 12683 31728
rect 10961 31723 11027 31726
rect 12617 31723 12683 31726
rect 15101 31786 15167 31789
rect 17953 31786 18019 31789
rect 15101 31784 18019 31786
rect 15101 31728 15106 31784
rect 15162 31728 17958 31784
rect 18014 31728 18019 31784
rect 15101 31726 18019 31728
rect 15101 31723 15167 31726
rect 17953 31723 18019 31726
rect 19425 31786 19491 31789
rect 20529 31786 20595 31789
rect 19425 31784 20595 31786
rect 19425 31728 19430 31784
rect 19486 31728 20534 31784
rect 20590 31728 20595 31784
rect 19425 31726 20595 31728
rect 19425 31723 19491 31726
rect 20529 31723 20595 31726
rect 6361 31652 6427 31653
rect 6310 31588 6316 31652
rect 6380 31650 6427 31652
rect 14917 31650 14983 31653
rect 16941 31650 17007 31653
rect 6380 31648 6472 31650
rect 6422 31592 6472 31648
rect 6380 31590 6472 31592
rect 14917 31648 17007 31650
rect 14917 31592 14922 31648
rect 14978 31592 16946 31648
rect 17002 31592 17007 31648
rect 14917 31590 17007 31592
rect 6380 31588 6427 31590
rect 6361 31587 6427 31588
rect 14917 31587 14983 31590
rect 16941 31587 17007 31590
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 10225 31514 10291 31517
rect 19425 31514 19491 31517
rect 10225 31512 19491 31514
rect 10225 31456 10230 31512
rect 10286 31456 19430 31512
rect 19486 31456 19491 31512
rect 10225 31454 19491 31456
rect 10225 31451 10291 31454
rect 19425 31451 19491 31454
rect 200 31378 800 31408
rect 1669 31378 1735 31381
rect 200 31376 1735 31378
rect 200 31320 1674 31376
rect 1730 31320 1735 31376
rect 200 31318 1735 31320
rect 200 31288 800 31318
rect 1669 31315 1735 31318
rect 10133 31378 10199 31381
rect 12157 31378 12223 31381
rect 10133 31376 12223 31378
rect 10133 31320 10138 31376
rect 10194 31320 12162 31376
rect 12218 31320 12223 31376
rect 10133 31318 12223 31320
rect 10133 31315 10199 31318
rect 12157 31315 12223 31318
rect 13077 31378 13143 31381
rect 16665 31378 16731 31381
rect 13077 31376 16731 31378
rect 13077 31320 13082 31376
rect 13138 31320 16670 31376
rect 16726 31320 16731 31376
rect 13077 31318 16731 31320
rect 13077 31315 13143 31318
rect 16665 31315 16731 31318
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 10869 30970 10935 30973
rect 12341 30970 12407 30973
rect 13997 30970 14063 30973
rect 10869 30968 14063 30970
rect 10869 30912 10874 30968
rect 10930 30912 12346 30968
rect 12402 30912 14002 30968
rect 14058 30912 14063 30968
rect 10869 30910 14063 30912
rect 10869 30907 10935 30910
rect 12341 30907 12407 30910
rect 13997 30907 14063 30910
rect 17401 30970 17467 30973
rect 21357 30970 21423 30973
rect 17401 30968 21423 30970
rect 17401 30912 17406 30968
rect 17462 30912 21362 30968
rect 21418 30912 21423 30968
rect 17401 30910 21423 30912
rect 17401 30907 17467 30910
rect 21357 30907 21423 30910
rect 1577 30834 1643 30837
rect 18413 30834 18479 30837
rect 1577 30832 18479 30834
rect 1577 30776 1582 30832
rect 1638 30776 18418 30832
rect 18474 30776 18479 30832
rect 1577 30774 18479 30776
rect 1577 30771 1643 30774
rect 18413 30771 18479 30774
rect 4061 30698 4127 30701
rect 6637 30698 6703 30701
rect 4061 30696 6703 30698
rect 4061 30640 4066 30696
rect 4122 30640 6642 30696
rect 6698 30640 6703 30696
rect 4061 30638 6703 30640
rect 4061 30635 4127 30638
rect 6637 30635 6703 30638
rect 11513 30698 11579 30701
rect 16665 30698 16731 30701
rect 18873 30698 18939 30701
rect 11513 30696 18939 30698
rect 11513 30640 11518 30696
rect 11574 30640 16670 30696
rect 16726 30640 18878 30696
rect 18934 30640 18939 30696
rect 11513 30638 18939 30640
rect 11513 30635 11579 30638
rect 16665 30635 16731 30638
rect 18873 30635 18939 30638
rect 20069 30562 20135 30565
rect 20345 30562 20411 30565
rect 20069 30560 20411 30562
rect 20069 30504 20074 30560
rect 20130 30504 20350 30560
rect 20406 30504 20411 30560
rect 20069 30502 20411 30504
rect 20069 30499 20135 30502
rect 20345 30499 20411 30502
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 3417 30426 3483 30429
rect 5717 30426 5783 30429
rect 3417 30424 5783 30426
rect 3417 30368 3422 30424
rect 3478 30368 5722 30424
rect 5778 30368 5783 30424
rect 3417 30366 5783 30368
rect 3417 30363 3483 30366
rect 5717 30363 5783 30366
rect 13997 30426 14063 30429
rect 17309 30426 17375 30429
rect 13997 30424 17375 30426
rect 13997 30368 14002 30424
rect 14058 30368 17314 30424
rect 17370 30368 17375 30424
rect 13997 30366 17375 30368
rect 13997 30363 14063 30366
rect 17309 30363 17375 30366
rect 10961 30292 11027 30293
rect 3918 30228 3924 30292
rect 3988 30290 3994 30292
rect 10910 30290 10916 30292
rect 3988 30230 10916 30290
rect 10980 30290 11027 30292
rect 15142 30290 15148 30292
rect 10980 30288 15148 30290
rect 11022 30232 15148 30288
rect 3988 30228 3994 30230
rect 10910 30228 10916 30230
rect 10980 30230 15148 30232
rect 10980 30228 11027 30230
rect 15142 30228 15148 30230
rect 15212 30228 15218 30292
rect 10961 30227 11027 30228
rect 4613 30156 4679 30157
rect 4613 30152 4660 30156
rect 4724 30154 4730 30156
rect 5901 30154 5967 30157
rect 6637 30154 6703 30157
rect 4613 30096 4618 30152
rect 4613 30092 4660 30096
rect 4724 30094 4770 30154
rect 5901 30152 6703 30154
rect 5901 30096 5906 30152
rect 5962 30096 6642 30152
rect 6698 30096 6703 30152
rect 5901 30094 6703 30096
rect 4724 30092 4730 30094
rect 4613 30091 4679 30092
rect 5901 30091 5967 30094
rect 6637 30091 6703 30094
rect 11145 30154 11211 30157
rect 14273 30154 14339 30157
rect 11145 30152 14339 30154
rect 11145 30096 11150 30152
rect 11206 30096 14278 30152
rect 14334 30096 14339 30152
rect 11145 30094 14339 30096
rect 11145 30091 11211 30094
rect 14273 30091 14339 30094
rect 200 30018 800 30048
rect 1669 30018 1735 30021
rect 200 30016 1735 30018
rect 200 29960 1674 30016
rect 1730 29960 1735 30016
rect 200 29958 1735 29960
rect 200 29928 800 29958
rect 1669 29955 1735 29958
rect 11329 30018 11395 30021
rect 12709 30018 12775 30021
rect 11329 30016 12775 30018
rect 11329 29960 11334 30016
rect 11390 29960 12714 30016
rect 12770 29960 12775 30016
rect 11329 29958 12775 29960
rect 11329 29955 11395 29958
rect 12709 29955 12775 29958
rect 38285 30018 38351 30021
rect 39200 30018 39800 30048
rect 38285 30016 39800 30018
rect 38285 29960 38290 30016
rect 38346 29960 39800 30016
rect 38285 29958 39800 29960
rect 38285 29955 38351 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 39200 29928 39800 29958
rect 34930 29887 35246 29888
rect 6637 29882 6703 29885
rect 8661 29882 8727 29885
rect 6637 29880 8727 29882
rect 6637 29824 6642 29880
rect 6698 29824 8666 29880
rect 8722 29824 8727 29880
rect 6637 29822 8727 29824
rect 6637 29819 6703 29822
rect 8661 29819 8727 29822
rect 10133 29882 10199 29885
rect 12801 29882 12867 29885
rect 16389 29882 16455 29885
rect 10133 29880 16455 29882
rect 10133 29824 10138 29880
rect 10194 29824 12806 29880
rect 12862 29824 16394 29880
rect 16450 29824 16455 29880
rect 10133 29822 16455 29824
rect 10133 29819 10199 29822
rect 12801 29819 12867 29822
rect 16389 29819 16455 29822
rect 3601 29748 3667 29749
rect 3550 29746 3556 29748
rect 3474 29686 3556 29746
rect 3620 29746 3667 29748
rect 9305 29746 9371 29749
rect 3620 29744 9371 29746
rect 3662 29688 9310 29744
rect 9366 29688 9371 29744
rect 3550 29684 3556 29686
rect 3620 29686 9371 29688
rect 3620 29684 3667 29686
rect 3601 29683 3667 29684
rect 9305 29683 9371 29686
rect 10409 29744 10475 29749
rect 10409 29688 10414 29744
rect 10470 29688 10475 29744
rect 10409 29683 10475 29688
rect 10777 29746 10843 29749
rect 14273 29746 14339 29749
rect 10777 29744 14339 29746
rect 10777 29688 10782 29744
rect 10838 29688 14278 29744
rect 14334 29688 14339 29744
rect 10777 29686 14339 29688
rect 10777 29683 10843 29686
rect 14273 29683 14339 29686
rect 15653 29746 15719 29749
rect 18045 29746 18111 29749
rect 15653 29744 18111 29746
rect 15653 29688 15658 29744
rect 15714 29688 18050 29744
rect 18106 29688 18111 29744
rect 15653 29686 18111 29688
rect 15653 29683 15719 29686
rect 18045 29683 18111 29686
rect 2405 29610 2471 29613
rect 8293 29610 8359 29613
rect 2405 29608 8359 29610
rect 2405 29552 2410 29608
rect 2466 29552 8298 29608
rect 8354 29552 8359 29608
rect 2405 29550 8359 29552
rect 10412 29610 10472 29683
rect 11237 29610 11303 29613
rect 10412 29608 11303 29610
rect 10412 29552 11242 29608
rect 11298 29552 11303 29608
rect 10412 29550 11303 29552
rect 2405 29547 2471 29550
rect 8293 29547 8359 29550
rect 11237 29547 11303 29550
rect 6269 29474 6335 29477
rect 6637 29474 6703 29477
rect 9581 29474 9647 29477
rect 6269 29472 6562 29474
rect 6269 29416 6274 29472
rect 6330 29416 6562 29472
rect 6269 29414 6562 29416
rect 6269 29411 6335 29414
rect 5625 29338 5691 29341
rect 6177 29338 6243 29341
rect 5625 29336 6243 29338
rect 5625 29280 5630 29336
rect 5686 29280 6182 29336
rect 6238 29280 6243 29336
rect 5625 29278 6243 29280
rect 6502 29338 6562 29414
rect 6637 29472 9647 29474
rect 6637 29416 6642 29472
rect 6698 29416 9586 29472
rect 9642 29416 9647 29472
rect 6637 29414 9647 29416
rect 6637 29411 6703 29414
rect 9581 29411 9647 29414
rect 9765 29472 9831 29477
rect 9765 29416 9770 29472
rect 9826 29416 9831 29472
rect 9765 29411 9831 29416
rect 7373 29338 7439 29341
rect 8017 29338 8083 29341
rect 6502 29336 8083 29338
rect 6502 29280 7378 29336
rect 7434 29280 8022 29336
rect 8078 29280 8083 29336
rect 6502 29278 8083 29280
rect 5625 29275 5691 29278
rect 6177 29275 6243 29278
rect 7373 29275 7439 29278
rect 8017 29275 8083 29278
rect 8293 29338 8359 29341
rect 9768 29338 9828 29411
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 8293 29336 9828 29338
rect 8293 29280 8298 29336
rect 8354 29280 9828 29336
rect 8293 29278 9828 29280
rect 11513 29338 11579 29341
rect 11973 29338 12039 29341
rect 11513 29336 12039 29338
rect 11513 29280 11518 29336
rect 11574 29280 11978 29336
rect 12034 29280 12039 29336
rect 11513 29278 12039 29280
rect 8293 29275 8359 29278
rect 11513 29275 11579 29278
rect 11973 29275 12039 29278
rect 20253 29338 20319 29341
rect 20437 29338 20503 29341
rect 20253 29336 20503 29338
rect 20253 29280 20258 29336
rect 20314 29280 20442 29336
rect 20498 29280 20503 29336
rect 20253 29278 20503 29280
rect 20253 29275 20319 29278
rect 20437 29275 20503 29278
rect 6177 29202 6243 29205
rect 6310 29202 6316 29204
rect 6177 29200 6316 29202
rect 6177 29144 6182 29200
rect 6238 29144 6316 29200
rect 6177 29142 6316 29144
rect 6177 29139 6243 29142
rect 6310 29140 6316 29142
rect 6380 29140 6386 29204
rect 6545 29202 6611 29205
rect 9765 29202 9831 29205
rect 6545 29200 9831 29202
rect 6545 29144 6550 29200
rect 6606 29144 9770 29200
rect 9826 29144 9831 29200
rect 6545 29142 9831 29144
rect 6545 29139 6611 29142
rect 9765 29139 9831 29142
rect 10409 29202 10475 29205
rect 10409 29200 17970 29202
rect 10409 29144 10414 29200
rect 10470 29144 17970 29200
rect 10409 29142 17970 29144
rect 10409 29139 10475 29142
rect 5257 29066 5323 29069
rect 6269 29066 6335 29069
rect 5257 29064 6335 29066
rect 5257 29008 5262 29064
rect 5318 29008 6274 29064
rect 6330 29008 6335 29064
rect 5257 29006 6335 29008
rect 5257 29003 5323 29006
rect 6269 29003 6335 29006
rect 6729 29066 6795 29069
rect 7925 29066 7991 29069
rect 6729 29064 7991 29066
rect 6729 29008 6734 29064
rect 6790 29008 7930 29064
rect 7986 29008 7991 29064
rect 6729 29006 7991 29008
rect 6729 29003 6795 29006
rect 7925 29003 7991 29006
rect 9029 29066 9095 29069
rect 10409 29066 10475 29069
rect 10542 29066 10548 29068
rect 9029 29064 9644 29066
rect 9029 29008 9034 29064
rect 9090 29008 9644 29064
rect 9029 29006 9644 29008
rect 9029 29003 9095 29006
rect 6269 28930 6335 28933
rect 9397 28930 9463 28933
rect 6269 28928 9463 28930
rect 6269 28872 6274 28928
rect 6330 28872 9402 28928
rect 9458 28872 9463 28928
rect 6269 28870 9463 28872
rect 9584 28930 9644 29006
rect 10409 29064 10548 29066
rect 10409 29008 10414 29064
rect 10470 29008 10548 29064
rect 10409 29006 10548 29008
rect 10409 29003 10475 29006
rect 10542 29004 10548 29006
rect 10612 29004 10618 29068
rect 14273 29066 14339 29069
rect 14273 29064 17050 29066
rect 14273 29008 14278 29064
rect 14334 29008 17050 29064
rect 14273 29006 17050 29008
rect 14273 29003 14339 29006
rect 14089 28930 14155 28933
rect 9584 28928 14155 28930
rect 9584 28872 14094 28928
rect 14150 28872 14155 28928
rect 9584 28870 14155 28872
rect 16990 28930 17050 29006
rect 17125 28930 17191 28933
rect 17401 28930 17467 28933
rect 16990 28928 17467 28930
rect 16990 28872 17130 28928
rect 17186 28872 17406 28928
rect 17462 28872 17467 28928
rect 16990 28870 17467 28872
rect 6269 28867 6335 28870
rect 9397 28867 9463 28870
rect 14089 28867 14155 28870
rect 17125 28867 17191 28870
rect 17401 28867 17467 28870
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 5349 28794 5415 28797
rect 11278 28794 11284 28796
rect 5349 28792 11284 28794
rect 5349 28736 5354 28792
rect 5410 28736 11284 28792
rect 5349 28734 11284 28736
rect 5349 28731 5415 28734
rect 11278 28732 11284 28734
rect 11348 28732 11354 28796
rect 11605 28794 11671 28797
rect 16665 28794 16731 28797
rect 11605 28792 16731 28794
rect 11605 28736 11610 28792
rect 11666 28736 16670 28792
rect 16726 28736 16731 28792
rect 11605 28734 16731 28736
rect 11605 28731 11671 28734
rect 16665 28731 16731 28734
rect 11145 28658 11211 28661
rect 13629 28658 13695 28661
rect 11145 28656 13695 28658
rect 11145 28600 11150 28656
rect 11206 28600 13634 28656
rect 13690 28600 13695 28656
rect 11145 28598 13695 28600
rect 17910 28658 17970 29142
rect 19374 29140 19380 29204
rect 19444 29202 19450 29204
rect 19609 29202 19675 29205
rect 19444 29200 19675 29202
rect 19444 29144 19614 29200
rect 19670 29144 19675 29200
rect 19444 29142 19675 29144
rect 19444 29140 19450 29142
rect 19609 29139 19675 29142
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 18597 28658 18663 28661
rect 17910 28656 18663 28658
rect 17910 28600 18602 28656
rect 18658 28600 18663 28656
rect 17910 28598 18663 28600
rect 11145 28595 11211 28598
rect 13629 28595 13695 28598
rect 18597 28595 18663 28598
rect 38285 28658 38351 28661
rect 39200 28658 39800 28688
rect 38285 28656 39800 28658
rect 38285 28600 38290 28656
rect 38346 28600 39800 28656
rect 38285 28598 39800 28600
rect 38285 28595 38351 28598
rect 39200 28568 39800 28598
rect 4705 28524 4771 28525
rect 4654 28460 4660 28524
rect 4724 28522 4771 28524
rect 6637 28522 6703 28525
rect 8385 28522 8451 28525
rect 11697 28522 11763 28525
rect 4724 28520 4816 28522
rect 4766 28464 4816 28520
rect 4724 28462 4816 28464
rect 6637 28520 11763 28522
rect 6637 28464 6642 28520
rect 6698 28464 8390 28520
rect 8446 28464 11702 28520
rect 11758 28464 11763 28520
rect 6637 28462 11763 28464
rect 4724 28460 4771 28462
rect 4705 28459 4771 28460
rect 6637 28459 6703 28462
rect 8385 28459 8451 28462
rect 11697 28459 11763 28462
rect 9213 28386 9279 28389
rect 10041 28386 10107 28389
rect 9213 28384 10107 28386
rect 9213 28328 9218 28384
rect 9274 28328 10046 28384
rect 10102 28328 10107 28384
rect 9213 28326 10107 28328
rect 9213 28323 9279 28326
rect 10041 28323 10107 28326
rect 11789 28386 11855 28389
rect 12525 28386 12591 28389
rect 11789 28384 12591 28386
rect 11789 28328 11794 28384
rect 11850 28328 12530 28384
rect 12586 28328 12591 28384
rect 11789 28326 12591 28328
rect 11789 28323 11855 28326
rect 12525 28323 12591 28326
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 14181 28250 14247 28253
rect 12206 28248 14247 28250
rect 12206 28192 14186 28248
rect 14242 28192 14247 28248
rect 12206 28190 14247 28192
rect 12206 28114 12266 28190
rect 14181 28187 14247 28190
rect 9492 28054 12266 28114
rect 12341 28114 12407 28117
rect 12525 28114 12591 28117
rect 12341 28112 12591 28114
rect 12341 28056 12346 28112
rect 12402 28056 12530 28112
rect 12586 28056 12591 28112
rect 12341 28054 12591 28056
rect 200 27978 800 28008
rect 1761 27978 1827 27981
rect 200 27976 1827 27978
rect 200 27920 1766 27976
rect 1822 27920 1827 27976
rect 200 27918 1827 27920
rect 200 27888 800 27918
rect 1761 27915 1827 27918
rect 3734 27916 3740 27980
rect 3804 27978 3810 27980
rect 9029 27978 9095 27981
rect 9492 27978 9552 28054
rect 12341 28051 12407 28054
rect 12525 28051 12591 28054
rect 12801 28114 12867 28117
rect 15694 28114 15700 28116
rect 12801 28112 15700 28114
rect 12801 28056 12806 28112
rect 12862 28056 15700 28112
rect 12801 28054 15700 28056
rect 12801 28051 12867 28054
rect 15694 28052 15700 28054
rect 15764 28114 15770 28116
rect 16113 28114 16179 28117
rect 15764 28112 16179 28114
rect 15764 28056 16118 28112
rect 16174 28056 16179 28112
rect 15764 28054 16179 28056
rect 15764 28052 15770 28054
rect 16113 28051 16179 28054
rect 3804 27976 9552 27978
rect 3804 27920 9034 27976
rect 9090 27920 9552 27976
rect 3804 27918 9552 27920
rect 3804 27916 3810 27918
rect 9029 27915 9095 27918
rect 10041 27842 10107 27845
rect 16849 27842 16915 27845
rect 10041 27840 16915 27842
rect 10041 27784 10046 27840
rect 10102 27784 16854 27840
rect 16910 27784 16915 27840
rect 10041 27782 16915 27784
rect 10041 27779 10107 27782
rect 16849 27779 16915 27782
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 10133 27706 10199 27709
rect 12249 27706 12315 27709
rect 10133 27704 12315 27706
rect 10133 27648 10138 27704
rect 10194 27648 12254 27704
rect 12310 27648 12315 27704
rect 10133 27646 12315 27648
rect 10133 27643 10199 27646
rect 12249 27643 12315 27646
rect 4061 27570 4127 27573
rect 9622 27570 9628 27572
rect 4061 27568 9628 27570
rect 4061 27512 4066 27568
rect 4122 27512 9628 27568
rect 4061 27510 9628 27512
rect 4061 27507 4127 27510
rect 9622 27508 9628 27510
rect 9692 27508 9698 27572
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 19701 27026 19767 27029
rect 23381 27026 23447 27029
rect 19701 27024 23447 27026
rect 19701 26968 19706 27024
rect 19762 26968 23386 27024
rect 23442 26968 23447 27024
rect 19701 26966 23447 26968
rect 19701 26963 19767 26966
rect 23381 26963 23447 26966
rect 10133 26890 10199 26893
rect 10685 26890 10751 26893
rect 10133 26888 10751 26890
rect 10133 26832 10138 26888
rect 10194 26832 10690 26888
rect 10746 26832 10751 26888
rect 10133 26830 10751 26832
rect 10133 26827 10199 26830
rect 10685 26827 10751 26830
rect 12525 26890 12591 26893
rect 12525 26888 12634 26890
rect 12525 26832 12530 26888
rect 12586 26832 12634 26888
rect 12525 26827 12634 26832
rect 7465 26754 7531 26757
rect 10225 26754 10291 26757
rect 10358 26754 10364 26756
rect 7465 26752 10364 26754
rect 7465 26696 7470 26752
rect 7526 26696 10230 26752
rect 10286 26696 10364 26752
rect 7465 26694 10364 26696
rect 7465 26691 7531 26694
rect 10225 26691 10291 26694
rect 10358 26692 10364 26694
rect 10428 26692 10434 26756
rect 4210 26688 4526 26689
rect 200 26618 800 26648
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 1669 26618 1735 26621
rect 200 26616 1735 26618
rect 200 26560 1674 26616
rect 1730 26560 1735 26616
rect 200 26558 1735 26560
rect 200 26528 800 26558
rect 1669 26555 1735 26558
rect 12433 26482 12499 26485
rect 12574 26482 12634 26827
rect 14457 26754 14523 26757
rect 18413 26754 18479 26757
rect 14457 26752 18479 26754
rect 14457 26696 14462 26752
rect 14518 26696 18418 26752
rect 18474 26696 18479 26752
rect 14457 26694 18479 26696
rect 14457 26691 14523 26694
rect 18413 26691 18479 26694
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 38193 26618 38259 26621
rect 39200 26618 39800 26648
rect 38193 26616 39800 26618
rect 38193 26560 38198 26616
rect 38254 26560 39800 26616
rect 38193 26558 39800 26560
rect 38193 26555 38259 26558
rect 39200 26528 39800 26558
rect 16205 26482 16271 26485
rect 17677 26482 17743 26485
rect 12433 26480 17743 26482
rect 12433 26424 12438 26480
rect 12494 26424 16210 26480
rect 16266 26424 17682 26480
rect 17738 26424 17743 26480
rect 12433 26422 17743 26424
rect 12433 26419 12499 26422
rect 16205 26419 16271 26422
rect 17677 26419 17743 26422
rect 19333 26346 19399 26349
rect 20897 26346 20963 26349
rect 19333 26344 20963 26346
rect 19333 26288 19338 26344
rect 19394 26288 20902 26344
rect 20958 26288 20963 26344
rect 19333 26286 20963 26288
rect 19333 26283 19399 26286
rect 20897 26283 20963 26286
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 12525 26074 12591 26077
rect 16941 26074 17007 26077
rect 17953 26074 18019 26077
rect 12525 26072 18019 26074
rect 12525 26016 12530 26072
rect 12586 26016 16946 26072
rect 17002 26016 17958 26072
rect 18014 26016 18019 26072
rect 12525 26014 18019 26016
rect 12525 26011 12591 26014
rect 16941 26011 17007 26014
rect 17953 26011 18019 26014
rect 11053 25802 11119 25805
rect 14365 25802 14431 25805
rect 11053 25800 14431 25802
rect 11053 25744 11058 25800
rect 11114 25744 14370 25800
rect 14426 25744 14431 25800
rect 11053 25742 14431 25744
rect 11053 25739 11119 25742
rect 14365 25739 14431 25742
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 10317 25258 10383 25261
rect 14273 25258 14339 25261
rect 10317 25256 14339 25258
rect 10317 25200 10322 25256
rect 10378 25200 14278 25256
rect 14334 25200 14339 25256
rect 10317 25198 14339 25200
rect 10317 25195 10383 25198
rect 14273 25195 14339 25198
rect 10133 25122 10199 25125
rect 12249 25122 12315 25125
rect 10133 25120 12315 25122
rect 10133 25064 10138 25120
rect 10194 25064 12254 25120
rect 12310 25064 12315 25120
rect 10133 25062 12315 25064
rect 10133 25059 10199 25062
rect 12249 25059 12315 25062
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 7281 24850 7347 24853
rect 15653 24850 15719 24853
rect 7281 24848 15719 24850
rect 7281 24792 7286 24848
rect 7342 24792 15658 24848
rect 15714 24792 15719 24848
rect 7281 24790 15719 24792
rect 7281 24787 7347 24790
rect 15653 24787 15719 24790
rect 13353 24714 13419 24717
rect 17677 24714 17743 24717
rect 13353 24712 17743 24714
rect 13353 24656 13358 24712
rect 13414 24656 17682 24712
rect 17738 24656 17743 24712
rect 13353 24654 17743 24656
rect 13353 24651 13419 24654
rect 17677 24651 17743 24654
rect 200 24578 800 24608
rect 1577 24578 1643 24581
rect 200 24576 1643 24578
rect 200 24520 1582 24576
rect 1638 24520 1643 24576
rect 200 24518 1643 24520
rect 200 24488 800 24518
rect 1577 24515 1643 24518
rect 8661 24578 8727 24581
rect 17585 24578 17651 24581
rect 8661 24576 17651 24578
rect 8661 24520 8666 24576
rect 8722 24520 17590 24576
rect 17646 24520 17651 24576
rect 8661 24518 17651 24520
rect 8661 24515 8727 24518
rect 17585 24515 17651 24518
rect 38285 24578 38351 24581
rect 39200 24578 39800 24608
rect 38285 24576 39800 24578
rect 38285 24520 38290 24576
rect 38346 24520 39800 24576
rect 38285 24518 39800 24520
rect 38285 24515 38351 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 39200 24488 39800 24518
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 10961 23898 11027 23901
rect 12709 23898 12775 23901
rect 10961 23896 12775 23898
rect 10961 23840 10966 23896
rect 11022 23840 12714 23896
rect 12770 23840 12775 23896
rect 10961 23838 12775 23840
rect 10961 23835 11027 23838
rect 12709 23835 12775 23838
rect 9673 23762 9739 23765
rect 9806 23762 9812 23764
rect 9673 23760 9812 23762
rect 9673 23704 9678 23760
rect 9734 23704 9812 23760
rect 9673 23702 9812 23704
rect 9673 23699 9739 23702
rect 9806 23700 9812 23702
rect 9876 23700 9882 23764
rect 11973 23762 12039 23765
rect 13997 23762 14063 23765
rect 11973 23760 14063 23762
rect 11973 23704 11978 23760
rect 12034 23704 14002 23760
rect 14058 23704 14063 23760
rect 11973 23702 14063 23704
rect 11973 23699 12039 23702
rect 13997 23699 14063 23702
rect 8385 23626 8451 23629
rect 11053 23626 11119 23629
rect 8385 23624 11119 23626
rect 8385 23568 8390 23624
rect 8446 23568 11058 23624
rect 11114 23568 11119 23624
rect 8385 23566 11119 23568
rect 8385 23563 8451 23566
rect 11053 23563 11119 23566
rect 11881 23626 11947 23629
rect 12617 23626 12683 23629
rect 11881 23624 12683 23626
rect 11881 23568 11886 23624
rect 11942 23568 12622 23624
rect 12678 23568 12683 23624
rect 11881 23566 12683 23568
rect 11881 23563 11947 23566
rect 12617 23563 12683 23566
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 4838 23156 4844 23220
rect 4908 23218 4914 23220
rect 13445 23218 13511 23221
rect 4908 23216 13511 23218
rect 4908 23160 13450 23216
rect 13506 23160 13511 23216
rect 4908 23158 13511 23160
rect 4908 23156 4914 23158
rect 13445 23155 13511 23158
rect 38193 23218 38259 23221
rect 39200 23218 39800 23248
rect 38193 23216 39800 23218
rect 38193 23160 38198 23216
rect 38254 23160 39800 23216
rect 38193 23158 39800 23160
rect 38193 23155 38259 23158
rect 39200 23128 39800 23158
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 15878 22748 15884 22812
rect 15948 22810 15954 22812
rect 18045 22810 18111 22813
rect 15948 22808 18111 22810
rect 15948 22752 18050 22808
rect 18106 22752 18111 22808
rect 15948 22750 18111 22752
rect 15948 22748 15954 22750
rect 18045 22747 18111 22750
rect 200 22538 800 22568
rect 1669 22538 1735 22541
rect 200 22536 1735 22538
rect 200 22480 1674 22536
rect 1730 22480 1735 22536
rect 200 22478 1735 22480
rect 200 22448 800 22478
rect 1669 22475 1735 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 10133 22130 10199 22133
rect 11697 22130 11763 22133
rect 12249 22130 12315 22133
rect 10133 22128 12315 22130
rect 10133 22072 10138 22128
rect 10194 22072 11702 22128
rect 11758 22072 12254 22128
rect 12310 22072 12315 22128
rect 10133 22070 12315 22072
rect 10133 22067 10199 22070
rect 11697 22067 11763 22070
rect 12249 22067 12315 22070
rect 15653 21994 15719 21997
rect 16389 21994 16455 21997
rect 15653 21992 16455 21994
rect 15653 21936 15658 21992
rect 15714 21936 16394 21992
rect 16450 21936 16455 21992
rect 15653 21934 16455 21936
rect 15653 21931 15719 21934
rect 16389 21931 16455 21934
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 200 21178 800 21208
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 1669 21178 1735 21181
rect 200 21176 1735 21178
rect 200 21120 1674 21176
rect 1730 21120 1735 21176
rect 200 21118 1735 21120
rect 200 21088 800 21118
rect 1669 21115 1735 21118
rect 38193 21178 38259 21181
rect 39200 21178 39800 21208
rect 38193 21176 39800 21178
rect 38193 21120 38198 21176
rect 38254 21120 39800 21176
rect 38193 21118 39800 21120
rect 38193 21115 38259 21118
rect 39200 21088 39800 21118
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 38193 19818 38259 19821
rect 39200 19818 39800 19848
rect 38193 19816 39800 19818
rect 38193 19760 38198 19816
rect 38254 19760 39800 19816
rect 38193 19758 39800 19760
rect 38193 19755 38259 19758
rect 39200 19728 39800 19758
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 200 19138 800 19168
rect 1669 19138 1735 19141
rect 200 19136 1735 19138
rect 200 19080 1674 19136
rect 1730 19080 1735 19136
rect 200 19078 1735 19080
rect 200 19048 800 19078
rect 1669 19075 1735 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 200 17778 800 17808
rect 1669 17778 1735 17781
rect 200 17776 1735 17778
rect 200 17720 1674 17776
rect 1730 17720 1735 17776
rect 200 17718 1735 17720
rect 200 17688 800 17718
rect 1669 17715 1735 17718
rect 39200 17688 39800 17808
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 200 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 1669 15738 1735 15741
rect 200 15736 1735 15738
rect 200 15680 1674 15736
rect 1730 15680 1735 15736
rect 200 15678 1735 15680
rect 200 15648 800 15678
rect 1669 15675 1735 15678
rect 38193 15738 38259 15741
rect 39200 15738 39800 15768
rect 38193 15736 39800 15738
rect 38193 15680 38198 15736
rect 38254 15680 39800 15736
rect 38193 15678 39800 15680
rect 38193 15675 38259 15678
rect 39200 15648 39800 15678
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 38285 14378 38351 14381
rect 39200 14378 39800 14408
rect 38285 14376 39800 14378
rect 38285 14320 38290 14376
rect 38346 14320 39800 14376
rect 38285 14318 39800 14320
rect 38285 14315 38351 14318
rect 39200 14288 39800 14318
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 200 13698 800 13728
rect 1669 13698 1735 13701
rect 200 13696 1735 13698
rect 200 13640 1674 13696
rect 1730 13640 1735 13696
rect 200 13638 1735 13640
rect 200 13608 800 13638
rect 1669 13635 1735 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 9806 12684 9812 12748
rect 9876 12746 9882 12748
rect 37457 12746 37523 12749
rect 9876 12744 37523 12746
rect 9876 12688 37462 12744
rect 37518 12688 37523 12744
rect 9876 12686 37523 12688
rect 9876 12684 9882 12686
rect 37457 12683 37523 12686
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 200 12338 800 12368
rect 1669 12338 1735 12341
rect 200 12336 1735 12338
rect 200 12280 1674 12336
rect 1730 12280 1735 12336
rect 200 12278 1735 12280
rect 200 12248 800 12278
rect 1669 12275 1735 12278
rect 38193 12338 38259 12341
rect 39200 12338 39800 12368
rect 38193 12336 39800 12338
rect 38193 12280 38198 12336
rect 38254 12280 39800 12336
rect 38193 12278 39800 12280
rect 38193 12275 38259 12278
rect 39200 12248 39800 12278
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 38193 10978 38259 10981
rect 39200 10978 39800 11008
rect 38193 10976 39800 10978
rect 38193 10920 38198 10976
rect 38254 10920 39800 10976
rect 38193 10918 39800 10920
rect 38193 10915 38259 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 39200 10888 39800 10918
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 200 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 1669 10298 1735 10301
rect 200 10296 1735 10298
rect 200 10240 1674 10296
rect 1730 10240 1735 10296
rect 200 10238 1735 10240
rect 200 10208 800 10238
rect 1669 10235 1735 10238
rect 10358 10236 10364 10300
rect 10428 10298 10434 10300
rect 12709 10298 12775 10301
rect 10428 10296 12775 10298
rect 10428 10240 12714 10296
rect 12770 10240 12775 10296
rect 10428 10238 12775 10240
rect 10428 10236 10434 10238
rect 12709 10235 12775 10238
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 200 8938 800 8968
rect 1669 8938 1735 8941
rect 200 8936 1735 8938
rect 200 8880 1674 8936
rect 1730 8880 1735 8936
rect 200 8878 1735 8880
rect 200 8848 800 8878
rect 1669 8875 1735 8878
rect 38193 8938 38259 8941
rect 39200 8938 39800 8968
rect 38193 8936 39800 8938
rect 38193 8880 38198 8936
rect 38254 8880 39800 8936
rect 38193 8878 39800 8880
rect 38193 8875 38259 8878
rect 39200 8848 39800 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 200 6898 800 6928
rect 1577 6898 1643 6901
rect 200 6896 1643 6898
rect 200 6840 1582 6896
rect 1638 6840 1643 6896
rect 200 6838 1643 6840
rect 200 6808 800 6838
rect 1577 6835 1643 6838
rect 38193 6898 38259 6901
rect 39200 6898 39800 6928
rect 38193 6896 39800 6898
rect 38193 6840 38198 6896
rect 38254 6840 39800 6896
rect 38193 6838 39800 6840
rect 38193 6835 38259 6838
rect 39200 6808 39800 6838
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 38193 5538 38259 5541
rect 39200 5538 39800 5568
rect 38193 5536 39800 5538
rect 38193 5480 38198 5536
rect 38254 5480 39800 5536
rect 38193 5478 39800 5480
rect 38193 5475 38259 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 39200 5448 39800 5478
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 200 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 1577 4858 1643 4861
rect 200 4856 1643 4858
rect 200 4800 1582 4856
rect 1638 4800 1643 4856
rect 200 4798 1643 4800
rect 200 4768 800 4798
rect 1577 4795 1643 4798
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 200 3498 800 3528
rect 1669 3498 1735 3501
rect 200 3496 1735 3498
rect 200 3440 1674 3496
rect 1730 3440 1735 3496
rect 200 3438 1735 3440
rect 200 3408 800 3438
rect 1669 3435 1735 3438
rect 38193 3498 38259 3501
rect 39200 3498 39800 3528
rect 38193 3496 39800 3498
rect 38193 3440 38198 3496
rect 38254 3440 39800 3496
rect 38193 3438 39800 3440
rect 38193 3435 38259 3438
rect 39200 3408 39800 3438
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 10910 2620 10916 2684
rect 10980 2682 10986 2684
rect 11881 2682 11947 2685
rect 10980 2680 11947 2682
rect 10980 2624 11886 2680
rect 11942 2624 11947 2680
rect 10980 2622 11947 2624
rect 10980 2620 10986 2622
rect 11881 2619 11947 2622
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 35801 2138 35867 2141
rect 39200 2138 39800 2168
rect 35801 2136 39800 2138
rect 35801 2080 35806 2136
rect 35862 2080 39800 2136
rect 35801 2078 39800 2080
rect 35801 2075 35867 2078
rect 39200 2048 39800 2078
rect 200 1458 800 1488
rect 1669 1458 1735 1461
rect 200 1456 1735 1458
rect 200 1400 1674 1456
rect 1730 1400 1735 1456
rect 200 1398 1735 1400
rect 200 1368 800 1398
rect 1669 1395 1735 1398
rect 37641 98 37707 101
rect 39200 98 39800 128
rect 37641 96 39800 98
rect 37641 40 37646 96
rect 37702 40 39800 96
rect 37641 38 39800 40
rect 37641 35 37707 38
rect 39200 8 39800 38
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 11284 36000 11348 36004
rect 11284 35944 11334 36000
rect 11334 35944 11348 36000
rect 11284 35940 11348 35944
rect 15884 36000 15948 36004
rect 15884 35944 15898 36000
rect 15898 35944 15948 36000
rect 15884 35940 15948 35944
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 15148 35668 15212 35732
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19380 34988 19444 35052
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 9628 34580 9692 34644
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 3556 33764 3620 33828
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 3740 33220 3804 33284
rect 9812 33280 9876 33284
rect 9812 33224 9862 33280
rect 9862 33224 9876 33280
rect 9812 33220 9876 33224
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 15700 32948 15764 33012
rect 10548 32676 10612 32740
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4844 32268 4908 32332
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 3924 31724 3988 31788
rect 6316 31648 6380 31652
rect 6316 31592 6366 31648
rect 6366 31592 6380 31648
rect 6316 31588 6380 31592
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 3924 30228 3988 30292
rect 10916 30288 10980 30292
rect 10916 30232 10966 30288
rect 10966 30232 10980 30288
rect 10916 30228 10980 30232
rect 15148 30228 15212 30292
rect 4660 30152 4724 30156
rect 4660 30096 4674 30152
rect 4674 30096 4724 30152
rect 4660 30092 4724 30096
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 3556 29744 3620 29748
rect 3556 29688 3606 29744
rect 3606 29688 3620 29744
rect 3556 29684 3620 29688
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 6316 29140 6380 29204
rect 10548 29004 10612 29068
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 11284 28732 11348 28796
rect 19380 29140 19444 29204
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 4660 28520 4724 28524
rect 4660 28464 4710 28520
rect 4710 28464 4724 28520
rect 4660 28460 4724 28464
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 3740 27916 3804 27980
rect 15700 28052 15764 28116
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 9628 27508 9692 27572
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 10364 26692 10428 26756
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 9812 23700 9876 23764
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 4844 23156 4908 23220
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 15884 22748 15948 22812
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 9812 12684 9876 12748
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 10364 10236 10428 10300
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 10916 2620 10980 2684
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 11283 36004 11349 36005
rect 11283 35940 11284 36004
rect 11348 35940 11349 36004
rect 11283 35939 11349 35940
rect 15883 36004 15949 36005
rect 15883 35940 15884 36004
rect 15948 35940 15949 36004
rect 15883 35939 15949 35940
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 9627 34644 9693 34645
rect 9627 34580 9628 34644
rect 9692 34580 9693 34644
rect 9627 34579 9693 34580
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 3555 33828 3621 33829
rect 3555 33764 3556 33828
rect 3620 33764 3621 33828
rect 3555 33763 3621 33764
rect 3558 29749 3618 33763
rect 3739 33284 3805 33285
rect 3739 33220 3740 33284
rect 3804 33220 3805 33284
rect 3739 33219 3805 33220
rect 3555 29748 3621 29749
rect 3555 29684 3556 29748
rect 3620 29684 3621 29748
rect 3555 29683 3621 29684
rect 3742 27981 3802 33219
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4843 32332 4909 32333
rect 4843 32268 4844 32332
rect 4908 32268 4909 32332
rect 4843 32267 4909 32268
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 3923 31788 3989 31789
rect 3923 31724 3924 31788
rect 3988 31724 3989 31788
rect 3923 31723 3989 31724
rect 3926 30293 3986 31723
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 3923 30292 3989 30293
rect 3923 30228 3924 30292
rect 3988 30228 3989 30292
rect 3923 30227 3989 30228
rect 4208 29952 4528 30976
rect 4659 30156 4725 30157
rect 4659 30092 4660 30156
rect 4724 30092 4725 30156
rect 4659 30091 4725 30092
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 3739 27980 3805 27981
rect 3739 27916 3740 27980
rect 3804 27916 3805 27980
rect 3739 27915 3805 27916
rect 4208 27776 4528 28800
rect 4662 28525 4722 30091
rect 4659 28524 4725 28525
rect 4659 28460 4660 28524
rect 4724 28460 4725 28524
rect 4659 28459 4725 28460
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4846 23221 4906 32267
rect 6315 31652 6381 31653
rect 6315 31588 6316 31652
rect 6380 31588 6381 31652
rect 6315 31587 6381 31588
rect 6318 29205 6378 31587
rect 6315 29204 6381 29205
rect 6315 29140 6316 29204
rect 6380 29140 6381 29204
rect 6315 29139 6381 29140
rect 9630 27573 9690 34579
rect 9811 33284 9877 33285
rect 9811 33220 9812 33284
rect 9876 33220 9877 33284
rect 9811 33219 9877 33220
rect 9627 27572 9693 27573
rect 9627 27508 9628 27572
rect 9692 27508 9693 27572
rect 9627 27507 9693 27508
rect 9814 23765 9874 33219
rect 10547 32740 10613 32741
rect 10547 32676 10548 32740
rect 10612 32676 10613 32740
rect 10547 32675 10613 32676
rect 10550 29069 10610 32675
rect 10915 30292 10981 30293
rect 10915 30228 10916 30292
rect 10980 30228 10981 30292
rect 10915 30227 10981 30228
rect 10547 29068 10613 29069
rect 10547 29004 10548 29068
rect 10612 29004 10613 29068
rect 10547 29003 10613 29004
rect 10363 26756 10429 26757
rect 10363 26692 10364 26756
rect 10428 26692 10429 26756
rect 10363 26691 10429 26692
rect 9811 23764 9877 23765
rect 9811 23700 9812 23764
rect 9876 23700 9877 23764
rect 9811 23699 9877 23700
rect 4843 23220 4909 23221
rect 4843 23156 4844 23220
rect 4908 23156 4909 23220
rect 4843 23155 4909 23156
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 9814 12749 9874 23699
rect 9811 12748 9877 12749
rect 9811 12684 9812 12748
rect 9876 12684 9877 12748
rect 9811 12683 9877 12684
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 10366 10301 10426 26691
rect 10363 10300 10429 10301
rect 10363 10236 10364 10300
rect 10428 10236 10429 10300
rect 10363 10235 10429 10236
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 10918 2685 10978 30227
rect 11286 28797 11346 35939
rect 15147 35732 15213 35733
rect 15147 35668 15148 35732
rect 15212 35668 15213 35732
rect 15147 35667 15213 35668
rect 15150 30293 15210 35667
rect 15699 33012 15765 33013
rect 15699 32948 15700 33012
rect 15764 32948 15765 33012
rect 15699 32947 15765 32948
rect 15147 30292 15213 30293
rect 15147 30228 15148 30292
rect 15212 30228 15213 30292
rect 15147 30227 15213 30228
rect 11283 28796 11349 28797
rect 11283 28732 11284 28796
rect 11348 28732 11349 28796
rect 11283 28731 11349 28732
rect 15702 28117 15762 32947
rect 15699 28116 15765 28117
rect 15699 28052 15700 28116
rect 15764 28052 15765 28116
rect 15699 28051 15765 28052
rect 15886 22813 15946 35939
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19379 35052 19445 35053
rect 19379 34988 19380 35052
rect 19444 34988 19445 35052
rect 19379 34987 19445 34988
rect 19382 29205 19442 34987
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19379 29204 19445 29205
rect 19379 29140 19380 29204
rect 19444 29140 19445 29204
rect 19379 29139 19445 29140
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 15883 22812 15949 22813
rect 15883 22748 15884 22812
rect 15948 22748 15949 22812
rect 15883 22747 15949 22748
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 10915 2684 10981 2685
rect 10915 2620 10916 2684
rect 10980 2620 10981 2684
rect 10915 2619 10981 2620
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__213__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 18676 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__223__A
timestamp 1667941163
transform -1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__224__A
timestamp 1667941163
transform -1 0 10580 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__A
timestamp 1667941163
transform -1 0 7452 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__A
timestamp 1667941163
transform -1 0 14076 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__A
timestamp 1667941163
transform 1 0 8004 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__A
timestamp 1667941163
transform 1 0 6532 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__232__A
timestamp 1667941163
transform 1 0 9200 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__A
timestamp 1667941163
transform 1 0 6532 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__A
timestamp 1667941163
transform -1 0 6716 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__A
timestamp 1667941163
transform -1 0 5520 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__A
timestamp 1667941163
transform -1 0 10212 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A
timestamp 1667941163
transform -1 0 12512 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__A
timestamp 1667941163
transform -1 0 10856 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__A
timestamp 1667941163
transform 1 0 12880 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__248__A
timestamp 1667941163
transform -1 0 24012 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__249__A
timestamp 1667941163
transform -1 0 24748 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__A
timestamp 1667941163
transform -1 0 23000 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__A
timestamp 1667941163
transform -1 0 24012 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__A
timestamp 1667941163
transform -1 0 22816 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__A
timestamp 1667941163
transform -1 0 18768 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__A
timestamp 1667941163
transform -1 0 12236 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__A
timestamp 1667941163
transform -1 0 6808 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__A
timestamp 1667941163
transform 1 0 21804 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__A
timestamp 1667941163
transform 1 0 14260 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__A
timestamp 1667941163
transform -1 0 18124 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__266__A
timestamp 1667941163
transform 1 0 22908 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__A
timestamp 1667941163
transform 1 0 21528 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__A
timestamp 1667941163
transform 1 0 19412 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__272__A
timestamp 1667941163
transform 1 0 18860 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__273__A
timestamp 1667941163
transform 1 0 6624 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__A
timestamp 1667941163
transform 1 0 17940 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__A
timestamp 1667941163
transform -1 0 21896 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__277__A
timestamp 1667941163
transform -1 0 17020 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__A
timestamp 1667941163
transform -1 0 9292 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__A
timestamp 1667941163
transform -1 0 17020 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__A
timestamp 1667941163
transform -1 0 17572 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__A
timestamp 1667941163
transform -1 0 23460 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__A
timestamp 1667941163
transform -1 0 20700 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__A
timestamp 1667941163
transform -1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__287__A
timestamp 1667941163
transform -1 0 7084 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__288__A
timestamp 1667941163
transform -1 0 21344 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__A
timestamp 1667941163
transform -1 0 17664 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__A
timestamp 1667941163
transform 1 0 12328 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__A
timestamp 1667941163
transform -1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__293__A
timestamp 1667941163
transform 1 0 21252 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__296__A
timestamp 1667941163
transform -1 0 22908 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__297__A
timestamp 1667941163
transform -1 0 23920 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__300__A
timestamp 1667941163
transform 1 0 21252 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__301__A
timestamp 1667941163
transform 1 0 22172 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__304__A
timestamp 1667941163
transform -1 0 8004 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__305__A
timestamp 1667941163
transform 1 0 19964 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__307__A
timestamp 1667941163
transform 1 0 21344 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__308__A
timestamp 1667941163
transform 1 0 22632 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__309__A
timestamp 1667941163
transform 1 0 6808 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__311__A
timestamp 1667941163
transform 1 0 22356 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__312__A
timestamp 1667941163
transform -1 0 23552 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__313__A
timestamp 1667941163
transform 1 0 8464 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__314__A
timestamp 1667941163
transform 1 0 21160 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__315__A
timestamp 1667941163
transform 1 0 21988 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__316__A
timestamp 1667941163
transform 1 0 7176 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__317__A
timestamp 1667941163
transform -1 0 13156 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__319__A
timestamp 1667941163
transform 1 0 11684 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__320__A
timestamp 1667941163
transform 1 0 6072 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__321__A
timestamp 1667941163
transform 1 0 11776 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__323__A
timestamp 1667941163
transform -1 0 10028 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__324__A
timestamp 1667941163
transform -1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__325__A
timestamp 1667941163
transform -1 0 14076 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__327__A
timestamp 1667941163
transform 1 0 14260 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__328__A
timestamp 1667941163
transform -1 0 23920 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__329__A
timestamp 1667941163
transform -1 0 16008 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__331__A
timestamp 1667941163
transform -1 0 22172 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__333__A
timestamp 1667941163
transform -1 0 11868 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__A
timestamp 1667941163
transform 1 0 19412 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__336__A
timestamp 1667941163
transform 1 0 15272 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__337__A
timestamp 1667941163
transform -1 0 20608 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__338__A
timestamp 1667941163
transform -1 0 15272 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__A
timestamp 1667941163
transform -1 0 16008 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__340__A
timestamp 1667941163
transform 1 0 7912 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__A
timestamp 1667941163
transform 1 0 12420 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__A
timestamp 1667941163
transform 1 0 17388 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__A
timestamp 1667941163
transform 1 0 30544 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__344__A
timestamp 1667941163
transform -1 0 20884 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__345__A
timestamp 1667941163
transform 1 0 17664 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__347__A
timestamp 1667941163
transform 1 0 6808 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__A
timestamp 1667941163
transform 1 0 22632 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__A
timestamp 1667941163
transform 1 0 7268 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__350__A
timestamp 1667941163
transform -1 0 15640 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__352__A
timestamp 1667941163
transform 1 0 7544 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__353__A
timestamp 1667941163
transform -1 0 23184 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__A
timestamp 1667941163
transform -1 0 21896 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__360__A
timestamp 1667941163
transform 1 0 9200 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__361__A
timestamp 1667941163
transform 1 0 11500 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__362__A
timestamp 1667941163
transform 1 0 24932 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__363__A
timestamp 1667941163
transform 1 0 22540 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__364__A
timestamp 1667941163
transform -1 0 8004 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__365__A
timestamp 1667941163
transform -1 0 33304 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__366__A
timestamp 1667941163
transform 1 0 17940 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__368__A
timestamp 1667941163
transform -1 0 22172 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__A
timestamp 1667941163
transform 1 0 22264 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__371__A
timestamp 1667941163
transform -1 0 16560 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__372__A
timestamp 1667941163
transform -1 0 35144 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__373__A
timestamp 1667941163
transform 1 0 11316 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__375__A
timestamp 1667941163
transform 1 0 7360 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__376__A
timestamp 1667941163
transform 1 0 17940 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__377__A
timestamp 1667941163
transform -1 0 33120 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__380__A
timestamp 1667941163
transform 1 0 22264 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__381__A
timestamp 1667941163
transform 1 0 13708 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__383__A
timestamp 1667941163
transform 1 0 23184 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__A
timestamp 1667941163
transform 1 0 7176 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__387__A
timestamp 1667941163
transform 1 0 27140 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__389__A
timestamp 1667941163
transform 1 0 21620 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__390__A
timestamp 1667941163
transform -1 0 3496 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__393__A
timestamp 1667941163
transform 1 0 2668 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__394__A
timestamp 1667941163
transform -1 0 2576 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__395__A
timestamp 1667941163
transform -1 0 1748 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__396__A
timestamp 1667941163
transform 1 0 4600 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__397__A
timestamp 1667941163
transform 1 0 4968 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__398__A
timestamp 1667941163
transform -1 0 21988 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__399__A
timestamp 1667941163
transform -1 0 1748 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__400__A
timestamp 1667941163
transform 1 0 4232 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__401__A
timestamp 1667941163
transform 1 0 2392 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__402__A
timestamp 1667941163
transform 1 0 6072 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__404__A
timestamp 1667941163
transform -1 0 3680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__405__A
timestamp 1667941163
transform 1 0 3864 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__406__A
timestamp 1667941163
transform 1 0 4876 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__407__A
timestamp 1667941163
transform 1 0 2760 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__408__A
timestamp 1667941163
transform 1 0 5152 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__409__A
timestamp 1667941163
transform 1 0 2668 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__410__A
timestamp 1667941163
transform -1 0 22724 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__411__A
timestamp 1667941163
transform 1 0 3220 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__412__A
timestamp 1667941163
transform 1 0 3404 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__413__A
timestamp 1667941163
transform -1 0 1840 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__415__A
timestamp 1667941163
transform 1 0 4416 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__416__A
timestamp 1667941163
transform 1 0 5152 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__417__A
timestamp 1667941163
transform 1 0 4140 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__418__A
timestamp 1667941163
transform 1 0 4232 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__419__A
timestamp 1667941163
transform 1 0 4232 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__420__A
timestamp 1667941163
transform 1 0 4508 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__421__A
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__A
timestamp 1667941163
transform 1 0 3312 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__423__A
timestamp 1667941163
transform -1 0 3128 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__424__A
timestamp 1667941163
transform 1 0 4048 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__426__A
timestamp 1667941163
transform -1 0 3404 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__427__A
timestamp 1667941163
transform 1 0 2392 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__428__A
timestamp 1667941163
transform 1 0 2944 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__429__A
timestamp 1667941163
transform 1 0 5428 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__430__A
timestamp 1667941163
transform 1 0 5888 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__431__A
timestamp 1667941163
transform 1 0 3312 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__432__A
timestamp 1667941163
transform 1 0 2116 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__433__A
timestamp 1667941163
transform 1 0 2760 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__434__A
timestamp 1667941163
transform 1 0 2208 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__435__A
timestamp 1667941163
transform -1 0 1748 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__437__A
timestamp 1667941163
transform -1 0 22172 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__438__A
timestamp 1667941163
transform 1 0 21804 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__439__A
timestamp 1667941163
transform 1 0 18400 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__440__A
timestamp 1667941163
transform -1 0 17572 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__441__A
timestamp 1667941163
transform 1 0 19688 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__442__A
timestamp 1667941163
transform 1 0 21252 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__443__A
timestamp 1667941163
transform 1 0 20608 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__444__A
timestamp 1667941163
transform 1 0 21344 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__445__A
timestamp 1667941163
transform -1 0 5704 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__446__A
timestamp 1667941163
transform -1 0 4968 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__464__CLK
timestamp 1667941163
transform 1 0 4048 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__465__CLK
timestamp 1667941163
transform 1 0 4600 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__466__CLK
timestamp 1667941163
transform 1 0 4600 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__466__D
timestamp 1667941163
transform 1 0 4784 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__467__CLK
timestamp 1667941163
transform 1 0 6440 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__467__D
timestamp 1667941163
transform -1 0 23092 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__468__CLK
timestamp 1667941163
transform 1 0 1564 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__468__D
timestamp 1667941163
transform -1 0 7544 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__469__CLK
timestamp 1667941163
transform 1 0 19964 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__469__D
timestamp 1667941163
transform -1 0 18860 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__470__CLK
timestamp 1667941163
transform 1 0 5428 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__471__CLK
timestamp 1667941163
transform 1 0 23092 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__472__CLK
timestamp 1667941163
transform 1 0 3312 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__472__D
timestamp 1667941163
transform 1 0 5336 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__473__CLK
timestamp 1667941163
transform 1 0 5888 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__473__D
timestamp 1667941163
transform -1 0 3772 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__474__CLK
timestamp 1667941163
transform 1 0 6532 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__474__D
timestamp 1667941163
transform -1 0 23644 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__475__CLK
timestamp 1667941163
transform 1 0 23552 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__476__CLK
timestamp 1667941163
transform 1 0 25116 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__476__D
timestamp 1667941163
transform -1 0 24748 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__477__CLK
timestamp 1667941163
transform 1 0 23828 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__478__CLK
timestamp 1667941163
transform 1 0 24564 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__478__D
timestamp 1667941163
transform -1 0 3680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__479__CLK
timestamp 1667941163
transform 1 0 24196 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__479__D
timestamp 1667941163
transform -1 0 22172 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__480__CLK
timestamp 1667941163
transform 1 0 3956 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__480__D
timestamp 1667941163
transform -1 0 24380 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__481__CLK
timestamp 1667941163
transform 1 0 22172 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__482__CLK
timestamp 1667941163
transform 1 0 23276 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__483__CLK
timestamp 1667941163
transform 1 0 24012 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__484__CLK
timestamp 1667941163
transform 1 0 21068 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__484__D
timestamp 1667941163
transform 1 0 20516 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__485__CLK
timestamp 1667941163
transform 1 0 5244 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__485__D
timestamp 1667941163
transform -1 0 6716 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__486__CLK
timestamp 1667941163
transform 1 0 22540 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__487__CLK
timestamp 1667941163
transform 1 0 20056 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__488__CLK
timestamp 1667941163
transform 1 0 21160 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__489__CLK
timestamp 1667941163
transform 1 0 19412 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__490__CLK
timestamp 1667941163
transform 1 0 20792 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__490__D
timestamp 1667941163
transform -1 0 19688 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__491__CLK
timestamp 1667941163
transform 1 0 4324 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__491__D
timestamp 1667941163
transform -1 0 5060 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__492__CLK
timestamp 1667941163
transform 1 0 23644 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__492__D
timestamp 1667941163
transform 1 0 23000 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__493__CLK
timestamp 1667941163
transform 1 0 19964 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__494__CLK
timestamp 1667941163
transform 1 0 23644 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__495__CLK
timestamp 1667941163
transform 1 0 2116 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__496__CLK
timestamp 1667941163
transform 1 0 4508 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__496__D
timestamp 1667941163
transform 1 0 3312 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__497__CLK
timestamp 1667941163
transform 1 0 6808 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__497__D
timestamp 1667941163
transform -1 0 4876 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__498__CLK
timestamp 1667941163
transform 1 0 23092 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__498__D
timestamp 1667941163
transform -1 0 22724 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__499__CLK
timestamp 1667941163
transform 1 0 21068 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__500__CLK
timestamp 1667941163
transform 1 0 24748 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__500__D
timestamp 1667941163
transform -1 0 24748 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__501__CLK
timestamp 1667941163
transform 1 0 24564 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__501__D
timestamp 1667941163
transform -1 0 25852 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__502__CLK
timestamp 1667941163
transform 1 0 24564 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__502__D
timestamp 1667941163
transform -1 0 23460 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__503__CLK
timestamp 1667941163
transform 1 0 22356 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__504__CLK
timestamp 1667941163
transform 1 0 5704 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__505__CLK
timestamp 1667941163
transform 1 0 23092 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__506__CLK
timestamp 1667941163
transform 1 0 21988 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__507__CLK
timestamp 1667941163
transform 1 0 22540 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__508__CLK
timestamp 1667941163
transform 1 0 23276 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__508__D
timestamp 1667941163
transform 1 0 22724 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__509__CLK
timestamp 1667941163
transform 1 0 20608 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__509__D
timestamp 1667941163
transform -1 0 20700 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__510__CLK
timestamp 1667941163
transform 1 0 21068 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__510__D
timestamp 1667941163
transform 1 0 22356 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__511__CLK
timestamp 1667941163
transform 1 0 22172 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__512__CLK
timestamp 1667941163
transform 1 0 24196 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__513__CLK
timestamp 1667941163
transform 1 0 3772 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__514__CLK
timestamp 1667941163
transform 1 0 4048 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__515__CLK
timestamp 1667941163
transform 1 0 23092 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__515__D
timestamp 1667941163
transform -1 0 21528 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__516__CLK
timestamp 1667941163
transform 1 0 20240 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__516__D
timestamp 1667941163
transform -1 0 20884 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__517__CLK
timestamp 1667941163
transform 1 0 21988 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__518__CLK
timestamp 1667941163
transform 1 0 22540 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__519__CLK
timestamp 1667941163
transform 1 0 22724 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__520__CLK
timestamp 1667941163
transform 1 0 23828 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__520__D
timestamp 1667941163
transform -1 0 22908 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__520__RESET_B
timestamp 1667941163
transform -1 0 21804 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__521__CLK
timestamp 1667941163
transform 1 0 22448 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__522__CLK
timestamp 1667941163
transform 1 0 5888 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__522__D
timestamp 1667941163
transform -1 0 6440 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__523__CLK
timestamp 1667941163
transform 1 0 22908 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__524__CLK
timestamp 1667941163
transform 1 0 23644 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__525__CLK
timestamp 1667941163
transform 1 0 23460 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__525__D
timestamp 1667941163
transform -1 0 24932 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__525__RESET_B
timestamp 1667941163
transform -1 0 23276 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__526__CLK
timestamp 1667941163
transform 1 0 5428 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__527__CLK
timestamp 1667941163
transform 1 0 21896 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__528__CLK
timestamp 1667941163
transform 1 0 21252 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__529__CLK
timestamp 1667941163
transform 1 0 22540 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__541__A
timestamp 1667941163
transform -1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__542__A
timestamp 1667941163
transform -1 0 18308 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__543__A
timestamp 1667941163
transform -1 0 20792 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__546__A
timestamp 1667941163
transform 1 0 20332 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__547__A
timestamp 1667941163
transform 1 0 12696 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__548__A
timestamp 1667941163
transform -1 0 17020 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__549__A
timestamp 1667941163
transform -1 0 30728 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__550__A
timestamp 1667941163
transform -1 0 22172 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__553__A
timestamp 1667941163
transform 1 0 21436 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__554__A
timestamp 1667941163
transform 1 0 18032 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__555__A
timestamp 1667941163
transform -1 0 25208 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__556__A
timestamp 1667941163
transform -1 0 20148 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__557__A
timestamp 1667941163
transform 1 0 23828 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__559__A
timestamp 1667941163
transform 1 0 16836 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__560__A
timestamp 1667941163
transform -1 0 19136 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__562__A
timestamp 1667941163
transform -1 0 7636 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__563__A
timestamp 1667941163
transform -1 0 20792 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__564__A
timestamp 1667941163
transform -1 0 6164 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__565__A
timestamp 1667941163
transform 1 0 5888 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__568__A
timestamp 1667941163
transform -1 0 34684 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__570__A
timestamp 1667941163
transform 1 0 24564 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__571__A
timestamp 1667941163
transform 1 0 4600 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__572__A
timestamp 1667941163
transform 1 0 38088 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__573__A
timestamp 1667941163
transform -1 0 16284 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__574__A
timestamp 1667941163
transform -1 0 26220 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__576__A
timestamp 1667941163
transform 1 0 19412 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__577__A
timestamp 1667941163
transform 1 0 2944 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__578__A
timestamp 1667941163
transform -1 0 6164 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__593__A
timestamp 1667941163
transform 1 0 16376 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__613__A
timestamp 1667941163
transform -1 0 8648 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__615__A
timestamp 1667941163
transform -1 0 19596 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__621__A
timestamp 1667941163
transform -1 0 18584 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__640__TE_B
timestamp 1667941163
transform -1 0 23368 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__653__A
timestamp 1667941163
transform -1 0 18032 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__671__A
timestamp 1667941163
transform 1 0 21988 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__693__A
timestamp 1667941163
transform 1 0 10672 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1667941163
transform -1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1667941163
transform -1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1667941163
transform -1 0 2852 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1667941163
transform -1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1667941163
transform -1 0 14536 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1667941163
transform -1 0 1748 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1667941163
transform -1 0 37628 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1667941163
transform -1 0 20332 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1667941163
transform -1 0 2300 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1667941163
transform -1 0 23828 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1667941163
transform -1 0 37628 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1667941163
transform -1 0 9384 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1667941163
transform -1 0 38364 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1667941163
transform -1 0 17756 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1667941163
transform -1 0 37628 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1667941163
transform -1 0 1748 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1667941163
transform 1 0 23920 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1667941163
transform -1 0 38364 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1667941163
transform -1 0 5336 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1667941163
transform -1 0 3036 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1667941163
transform -1 0 21804 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1667941163
transform -1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1667941163
transform -1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1667941163
transform -1 0 33212 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1667941163
transform -1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1667941163
transform -1 0 37628 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1667941163
transform -1 0 1748 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1667941163
transform -1 0 25484 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1667941163
transform -1 0 37628 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1667941163
transform -1 0 1748 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1667941163
transform -1 0 37628 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1667941163
transform -1 0 2392 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1667941163
transform -1 0 29716 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1667941163
transform -1 0 38364 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1667941163
transform -1 0 20700 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1667941163
transform -1 0 24380 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1667941163
transform -1 0 17756 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1667941163
transform -1 0 2484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1667941163
transform -1 0 22908 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1667941163
transform -1 0 29992 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output49_A
timestamp 1667941163
transform -1 0 37628 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output56_A
timestamp 1667941163
transform -1 0 26680 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output57_A
timestamp 1667941163
transform -1 0 35236 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output58_A
timestamp 1667941163
transform -1 0 2484 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output59_A
timestamp 1667941163
transform 1 0 37444 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output64_A
timestamp 1667941163
transform 1 0 5612 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output74_A
timestamp 1667941163
transform 1 0 2300 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output79_A
timestamp 1667941163
transform -1 0 37628 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output80_A
timestamp 1667941163
transform -1 0 2484 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output82_A
timestamp 1667941163
transform 1 0 7268 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output86_A
timestamp 1667941163
transform 1 0 21344 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output87_A
timestamp 1667941163
transform -1 0 31832 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2668 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1667941163
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41
timestamp 1667941163
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49
timestamp 1667941163
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1667941163
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63
timestamp 1667941163
transform 1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 7452 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77
timestamp 1667941163
transform 1 0 8188 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1667941163
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_85 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90
timestamp 1667941163
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_104
timestamp 1667941163
transform 1 0 10672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1667941163
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119
timestamp 1667941163
transform 1 0 12052 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_127
timestamp 1667941163
transform 1 0 12788 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_133
timestamp 1667941163
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1667941163
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1667941163
transform 1 0 14536 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 15272 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1667941163
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1667941163
transform 1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181
timestamp 1667941163
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_189
timestamp 1667941163
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1667941163
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_205
timestamp 1667941163
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_210
timestamp 1667941163
transform 1 0 20424 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1667941163
transform 1 0 21160 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1667941163
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_231
timestamp 1667941163
transform 1 0 22356 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_237
timestamp 1667941163
transform 1 0 22908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_245
timestamp 1667941163
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1667941163
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_261
timestamp 1667941163
transform 1 0 25116 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_266
timestamp 1667941163
transform 1 0 25576 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1667941163
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_287
timestamp 1667941163
transform 1 0 27508 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_295
timestamp 1667941163
transform 1 0 28244 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1667941163
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1667941163
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_321
timestamp 1667941163
transform 1 0 30636 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_329
timestamp 1667941163
transform 1 0 31372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_334
timestamp 1667941163
transform 1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_343
timestamp 1667941163
transform 1 0 32660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_349
timestamp 1667941163
transform 1 0 33212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_357
timestamp 1667941163
transform 1 0 33948 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1667941163
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_371
timestamp 1667941163
transform 1 0 35236 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_377
timestamp 1667941163
transform 1 0 35788 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_382
timestamp 1667941163
transform 1 0 36248 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1667941163
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_399
timestamp 1667941163
transform 1 0 37812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_405
timestamp 1667941163
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1667941163
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_15
timestamp 1667941163
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_21
timestamp 1667941163
transform 1 0 3036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_33
timestamp 1667941163
transform 1 0 4140 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_45
timestamp 1667941163
transform 1 0 5244 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1667941163
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1667941163
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_69
timestamp 1667941163
transform 1 0 7452 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_77
timestamp 1667941163
transform 1 0 8188 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_82
timestamp 1667941163
transform 1 0 8648 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_94
timestamp 1667941163
transform 1 0 9752 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_106
timestamp 1667941163
transform 1 0 10856 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_125
timestamp 1667941163
transform 1 0 12604 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1667941163
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1667941163
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1667941163
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1667941163
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1667941163
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1667941163
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_208
timestamp 1667941163
transform 1 0 20240 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_214
timestamp 1667941163
transform 1 0 20792 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1667941163
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1667941163
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1667941163
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1667941163
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1667941163
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1667941163
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1667941163
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_305
timestamp 1667941163
transform 1 0 29164 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_311
timestamp 1667941163
transform 1 0 29716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_323
timestamp 1667941163
transform 1 0 30820 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1667941163
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_349
timestamp 1667941163
transform 1 0 33212 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_355
timestamp 1667941163
transform 1 0 33764 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_359
timestamp 1667941163
transform 1 0 34132 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_365
timestamp 1667941163
transform 1 0 34684 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_371
timestamp 1667941163
transform 1 0 35236 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_383
timestamp 1667941163
transform 1 0 36340 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1667941163
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_397
timestamp 1667941163
transform 1 0 37628 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_9
timestamp 1667941163
transform 1 0 1932 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1667941163
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1667941163
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1667941163
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1667941163
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1667941163
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1667941163
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1667941163
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1667941163
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1667941163
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1667941163
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1667941163
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1667941163
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1667941163
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1667941163
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1667941163
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1667941163
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1667941163
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1667941163
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1667941163
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1667941163
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1667941163
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1667941163
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1667941163
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1667941163
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1667941163
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1667941163
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1667941163
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1667941163
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1667941163
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1667941163
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1667941163
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1667941163
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_389
timestamp 1667941163
transform 1 0 36892 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_397
timestamp 1667941163
transform 1 0 37628 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_405
timestamp 1667941163
transform 1 0 38364 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1667941163
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1667941163
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1667941163
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1667941163
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1667941163
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1667941163
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1667941163
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1667941163
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1667941163
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1667941163
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1667941163
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1667941163
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1667941163
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1667941163
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1667941163
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1667941163
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1667941163
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1667941163
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1667941163
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1667941163
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1667941163
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1667941163
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1667941163
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1667941163
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1667941163
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1667941163
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1667941163
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1667941163
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1667941163
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1667941163
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1667941163
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1667941163
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1667941163
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1667941163
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7
timestamp 1667941163
transform 1 0 1748 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_19
timestamp 1667941163
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1667941163
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1667941163
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1667941163
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1667941163
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1667941163
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1667941163
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1667941163
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1667941163
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1667941163
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1667941163
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1667941163
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1667941163
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1667941163
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1667941163
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1667941163
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1667941163
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1667941163
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1667941163
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1667941163
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1667941163
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1667941163
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1667941163
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1667941163
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1667941163
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1667941163
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1667941163
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1667941163
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1667941163
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1667941163
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1667941163
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1667941163
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_401
timestamp 1667941163
transform 1 0 37996 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_9
timestamp 1667941163
transform 1 0 1932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_21
timestamp 1667941163
transform 1 0 3036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_33
timestamp 1667941163
transform 1 0 4140 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_45
timestamp 1667941163
transform 1 0 5244 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1667941163
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1667941163
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1667941163
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1667941163
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1667941163
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1667941163
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1667941163
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1667941163
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1667941163
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1667941163
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1667941163
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1667941163
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1667941163
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1667941163
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1667941163
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1667941163
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1667941163
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1667941163
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1667941163
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1667941163
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1667941163
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1667941163
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1667941163
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1667941163
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1667941163
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1667941163
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1667941163
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1667941163
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1667941163
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1667941163
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1667941163
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1667941163
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1667941163
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1667941163
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1667941163
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1667941163
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1667941163
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1667941163
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1667941163
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1667941163
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1667941163
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1667941163
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1667941163
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1667941163
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1667941163
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1667941163
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1667941163
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1667941163
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1667941163
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1667941163
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1667941163
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1667941163
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1667941163
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1667941163
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1667941163
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1667941163
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1667941163
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1667941163
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1667941163
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1667941163
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1667941163
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1667941163
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1667941163
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1667941163
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1667941163
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_389
timestamp 1667941163
transform 1 0 36892 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_397
timestamp 1667941163
transform 1 0 37628 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_405
timestamp 1667941163
transform 1 0 38364 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1667941163
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1667941163
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1667941163
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1667941163
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1667941163
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1667941163
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1667941163
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1667941163
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1667941163
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1667941163
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1667941163
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1667941163
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1667941163
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1667941163
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1667941163
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1667941163
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1667941163
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1667941163
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1667941163
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1667941163
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1667941163
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1667941163
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1667941163
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1667941163
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1667941163
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1667941163
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1667941163
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1667941163
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1667941163
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1667941163
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_342
timestamp 1667941163
transform 1 0 32568 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_348
timestamp 1667941163
transform 1 0 33120 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_360
timestamp 1667941163
transform 1 0 34224 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_372
timestamp 1667941163
transform 1 0 35328 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_384
timestamp 1667941163
transform 1 0 36432 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7
timestamp 1667941163
transform 1 0 1748 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_19
timestamp 1667941163
transform 1 0 2852 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1667941163
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1667941163
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_53
timestamp 1667941163
transform 1 0 5980 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_62
timestamp 1667941163
transform 1 0 6808 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_68
timestamp 1667941163
transform 1 0 7360 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1667941163
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1667941163
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1667941163
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1667941163
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1667941163
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1667941163
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1667941163
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1667941163
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1667941163
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1667941163
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1667941163
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1667941163
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1667941163
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1667941163
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_248
timestamp 1667941163
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_257
timestamp 1667941163
transform 1 0 24748 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_269
timestamp 1667941163
transform 1 0 25852 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_281
timestamp 1667941163
transform 1 0 26956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_293
timestamp 1667941163
transform 1 0 28060 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_305
timestamp 1667941163
transform 1 0 29164 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1667941163
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1667941163
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1667941163
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1667941163
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1667941163
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1667941163
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_401
timestamp 1667941163
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_9
timestamp 1667941163
transform 1 0 1932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_21
timestamp 1667941163
transform 1 0 3036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_33
timestamp 1667941163
transform 1 0 4140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_45
timestamp 1667941163
transform 1 0 5244 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1667941163
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1667941163
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1667941163
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1667941163
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1667941163
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1667941163
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1667941163
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1667941163
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1667941163
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1667941163
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1667941163
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1667941163
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1667941163
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1667941163
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1667941163
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1667941163
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1667941163
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1667941163
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1667941163
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1667941163
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1667941163
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1667941163
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1667941163
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1667941163
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1667941163
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1667941163
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1667941163
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1667941163
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1667941163
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1667941163
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_397
timestamp 1667941163
transform 1 0 37628 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1667941163
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1667941163
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1667941163
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1667941163
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1667941163
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1667941163
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1667941163
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1667941163
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1667941163
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1667941163
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1667941163
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1667941163
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1667941163
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1667941163
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1667941163
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1667941163
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1667941163
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1667941163
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1667941163
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1667941163
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1667941163
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1667941163
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1667941163
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1667941163
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1667941163
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1667941163
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1667941163
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1667941163
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1667941163
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1667941163
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1667941163
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1667941163
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1667941163
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_401
timestamp 1667941163
transform 1 0 37996 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_7
timestamp 1667941163
transform 1 0 1748 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_19
timestamp 1667941163
transform 1 0 2852 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_31
timestamp 1667941163
transform 1 0 3956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_43
timestamp 1667941163
transform 1 0 5060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1667941163
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1667941163
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1667941163
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1667941163
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1667941163
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1667941163
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1667941163
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1667941163
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1667941163
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1667941163
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1667941163
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1667941163
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1667941163
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1667941163
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1667941163
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1667941163
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1667941163
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1667941163
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1667941163
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1667941163
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1667941163
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1667941163
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1667941163
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1667941163
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1667941163
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1667941163
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1667941163
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1667941163
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1667941163
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_9
timestamp 1667941163
transform 1 0 1932 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_21
timestamp 1667941163
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1667941163
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1667941163
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1667941163
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1667941163
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1667941163
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1667941163
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1667941163
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1667941163
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1667941163
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1667941163
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1667941163
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1667941163
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1667941163
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1667941163
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1667941163
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1667941163
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1667941163
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1667941163
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1667941163
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1667941163
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1667941163
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1667941163
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1667941163
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1667941163
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1667941163
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1667941163
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1667941163
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1667941163
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1667941163
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1667941163
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1667941163
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1667941163
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_405
timestamp 1667941163
transform 1 0 38364 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1667941163
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1667941163
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1667941163
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1667941163
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1667941163
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1667941163
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1667941163
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1667941163
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1667941163
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1667941163
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1667941163
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1667941163
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1667941163
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1667941163
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1667941163
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1667941163
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1667941163
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_205
timestamp 1667941163
transform 1 0 19964 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_215
timestamp 1667941163
transform 1 0 20884 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1667941163
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1667941163
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1667941163
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1667941163
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1667941163
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1667941163
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1667941163
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1667941163
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1667941163
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1667941163
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1667941163
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1667941163
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1667941163
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1667941163
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1667941163
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1667941163
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1667941163
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1667941163
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1667941163
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1667941163
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1667941163
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1667941163
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_93
timestamp 1667941163
transform 1 0 9660 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1667941163
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1667941163
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_121
timestamp 1667941163
transform 1 0 12236 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_125
timestamp 1667941163
transform 1 0 12604 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_128
timestamp 1667941163
transform 1 0 12880 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_135
timestamp 1667941163
transform 1 0 13524 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1667941163
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1667941163
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1667941163
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1667941163
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1667941163
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1667941163
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1667941163
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1667941163
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1667941163
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1667941163
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1667941163
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1667941163
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1667941163
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1667941163
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1667941163
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1667941163
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1667941163
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1667941163
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1667941163
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1667941163
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1667941163
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1667941163
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_401
timestamp 1667941163
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_9
timestamp 1667941163
transform 1 0 1932 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1667941163
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1667941163
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1667941163
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1667941163
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1667941163
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1667941163
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1667941163
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1667941163
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1667941163
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1667941163
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_125
timestamp 1667941163
transform 1 0 12604 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_129
timestamp 1667941163
transform 1 0 12972 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_133
timestamp 1667941163
transform 1 0 13340 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_139
timestamp 1667941163
transform 1 0 13892 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_151
timestamp 1667941163
transform 1 0 14996 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_163
timestamp 1667941163
transform 1 0 16100 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1667941163
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1667941163
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1667941163
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1667941163
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1667941163
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1667941163
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1667941163
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1667941163
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1667941163
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1667941163
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1667941163
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1667941163
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1667941163
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1667941163
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1667941163
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1667941163
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1667941163
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1667941163
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1667941163
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1667941163
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1667941163
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1667941163
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1667941163
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1667941163
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1667941163
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1667941163
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1667941163
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1667941163
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1667941163
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1667941163
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1667941163
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1667941163
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1667941163
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1667941163
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1667941163
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1667941163
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1667941163
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1667941163
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1667941163
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1667941163
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1667941163
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1667941163
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1667941163
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1667941163
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1667941163
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1667941163
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1667941163
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1667941163
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1667941163
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1667941163
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1667941163
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_389
timestamp 1667941163
transform 1 0 36892 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_397
timestamp 1667941163
transform 1 0 37628 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_405
timestamp 1667941163
transform 1 0 38364 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1667941163
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1667941163
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1667941163
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1667941163
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1667941163
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1667941163
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1667941163
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1667941163
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1667941163
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1667941163
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1667941163
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1667941163
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1667941163
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1667941163
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1667941163
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1667941163
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1667941163
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1667941163
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1667941163
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1667941163
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1667941163
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_249
timestamp 1667941163
transform 1 0 24012 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_255
timestamp 1667941163
transform 1 0 24564 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1667941163
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1667941163
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1667941163
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1667941163
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1667941163
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1667941163
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1667941163
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1667941163
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1667941163
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1667941163
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1667941163
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1667941163
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1667941163
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1667941163
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1667941163
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1667941163
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1667941163
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1667941163
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1667941163
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1667941163
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1667941163
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1667941163
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1667941163
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1667941163
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1667941163
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_153
timestamp 1667941163
transform 1 0 15180 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_159
timestamp 1667941163
transform 1 0 15732 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1667941163
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1667941163
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1667941163
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1667941163
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1667941163
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1667941163
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1667941163
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1667941163
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1667941163
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1667941163
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1667941163
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1667941163
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1667941163
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1667941163
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1667941163
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1667941163
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1667941163
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1667941163
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1667941163
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_389
timestamp 1667941163
transform 1 0 36892 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_397
timestamp 1667941163
transform 1 0 37628 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_402
timestamp 1667941163
transform 1 0 38088 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_406
timestamp 1667941163
transform 1 0 38456 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_9
timestamp 1667941163
transform 1 0 1932 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_21
timestamp 1667941163
transform 1 0 3036 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_33
timestamp 1667941163
transform 1 0 4140 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_45
timestamp 1667941163
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1667941163
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1667941163
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1667941163
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1667941163
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1667941163
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1667941163
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1667941163
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1667941163
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1667941163
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_161
timestamp 1667941163
transform 1 0 15916 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1667941163
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_173
timestamp 1667941163
transform 1 0 17020 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_185
timestamp 1667941163
transform 1 0 18124 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_197
timestamp 1667941163
transform 1 0 19228 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_209
timestamp 1667941163
transform 1 0 20332 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_221
timestamp 1667941163
transform 1 0 21436 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1667941163
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1667941163
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1667941163
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1667941163
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1667941163
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1667941163
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1667941163
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1667941163
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1667941163
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1667941163
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1667941163
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1667941163
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1667941163
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1667941163
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_397
timestamp 1667941163
transform 1 0 37628 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1667941163
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1667941163
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1667941163
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1667941163
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1667941163
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1667941163
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1667941163
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1667941163
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1667941163
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1667941163
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_121
timestamp 1667941163
transform 1 0 12236 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_129
timestamp 1667941163
transform 1 0 12972 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_134
timestamp 1667941163
transform 1 0 13432 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1667941163
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1667941163
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1667941163
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1667941163
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1667941163
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_201
timestamp 1667941163
transform 1 0 19596 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_205
timestamp 1667941163
transform 1 0 19964 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_211
timestamp 1667941163
transform 1 0 20516 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_223
timestamp 1667941163
transform 1 0 21620 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_235
timestamp 1667941163
transform 1 0 22724 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_247
timestamp 1667941163
transform 1 0 23828 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1667941163
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1667941163
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1667941163
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1667941163
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1667941163
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1667941163
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1667941163
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1667941163
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1667941163
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1667941163
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1667941163
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_401
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_9
timestamp 1667941163
transform 1 0 1932 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_21
timestamp 1667941163
transform 1 0 3036 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_33
timestamp 1667941163
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_45
timestamp 1667941163
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1667941163
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1667941163
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1667941163
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1667941163
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1667941163
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1667941163
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1667941163
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1667941163
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1667941163
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1667941163
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1667941163
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1667941163
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1667941163
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1667941163
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1667941163
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1667941163
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1667941163
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1667941163
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1667941163
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1667941163
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1667941163
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1667941163
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1667941163
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1667941163
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1667941163
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1667941163
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1667941163
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1667941163
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_401
timestamp 1667941163
transform 1 0 37996 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1667941163
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1667941163
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1667941163
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1667941163
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1667941163
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1667941163
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1667941163
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1667941163
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1667941163
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1667941163
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1667941163
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1667941163
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1667941163
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1667941163
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1667941163
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1667941163
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1667941163
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1667941163
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1667941163
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1667941163
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1667941163
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1667941163
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1667941163
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1667941163
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1667941163
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1667941163
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1667941163
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1667941163
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1667941163
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1667941163
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1667941163
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1667941163
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1667941163
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_389
timestamp 1667941163
transform 1 0 36892 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_405
timestamp 1667941163
transform 1 0 38364 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1667941163
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1667941163
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1667941163
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1667941163
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1667941163
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1667941163
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1667941163
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1667941163
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1667941163
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1667941163
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1667941163
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1667941163
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1667941163
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1667941163
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1667941163
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1667941163
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1667941163
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1667941163
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1667941163
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1667941163
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1667941163
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1667941163
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1667941163
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1667941163
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1667941163
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1667941163
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1667941163
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1667941163
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1667941163
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1667941163
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1667941163
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1667941163
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1667941163
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1667941163
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1667941163
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1667941163
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1667941163
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1667941163
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1667941163
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1667941163
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1667941163
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1667941163
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1667941163
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1667941163
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1667941163
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1667941163
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1667941163
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1667941163
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1667941163
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1667941163
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1667941163
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1667941163
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1667941163
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1667941163
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1667941163
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1667941163
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1667941163
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1667941163
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1667941163
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1667941163
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1667941163
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1667941163
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1667941163
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1667941163
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1667941163
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1667941163
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1667941163
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1667941163
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_401
timestamp 1667941163
transform 1 0 37996 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_9
timestamp 1667941163
transform 1 0 1932 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_21
timestamp 1667941163
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_33
timestamp 1667941163
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1667941163
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1667941163
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1667941163
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1667941163
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1667941163
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1667941163
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1667941163
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1667941163
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1667941163
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1667941163
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1667941163
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1667941163
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1667941163
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1667941163
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1667941163
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1667941163
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1667941163
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1667941163
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1667941163
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1667941163
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1667941163
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1667941163
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1667941163
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1667941163
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1667941163
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1667941163
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1667941163
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1667941163
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1667941163
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1667941163
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1667941163
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1667941163
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1667941163
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1667941163
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1667941163
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1667941163
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1667941163
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1667941163
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1667941163
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1667941163
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1667941163
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1667941163
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1667941163
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1667941163
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1667941163
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1667941163
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1667941163
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1667941163
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1667941163
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_209
timestamp 1667941163
transform 1 0 20332 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_220
timestamp 1667941163
transform 1 0 21344 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_226
timestamp 1667941163
transform 1 0 21896 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_238
timestamp 1667941163
transform 1 0 23000 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1667941163
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1667941163
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1667941163
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1667941163
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1667941163
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1667941163
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1667941163
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1667941163
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1667941163
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1667941163
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1667941163
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1667941163
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_401
timestamp 1667941163
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1667941163
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1667941163
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1667941163
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1667941163
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1667941163
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1667941163
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1667941163
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1667941163
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1667941163
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1667941163
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1667941163
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_137
timestamp 1667941163
transform 1 0 13708 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_141
timestamp 1667941163
transform 1 0 14076 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_148
timestamp 1667941163
transform 1 0 14720 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_154
timestamp 1667941163
transform 1 0 15272 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1667941163
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1667941163
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1667941163
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1667941163
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1667941163
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1667941163
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1667941163
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_249
timestamp 1667941163
transform 1 0 24012 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_257
timestamp 1667941163
transform 1 0 24748 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_262
timestamp 1667941163
transform 1 0 25208 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_270
timestamp 1667941163
transform 1 0 25944 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1667941163
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1667941163
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1667941163
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1667941163
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1667941163
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1667941163
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1667941163
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1667941163
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1667941163
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1667941163
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1667941163
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1667941163
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1667941163
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1667941163
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1667941163
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1667941163
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1667941163
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1667941163
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1667941163
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1667941163
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1667941163
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_121
timestamp 1667941163
transform 1 0 12236 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_131
timestamp 1667941163
transform 1 0 13156 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1667941163
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_152
timestamp 1667941163
transform 1 0 15088 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_158
timestamp 1667941163
transform 1 0 15640 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_170
timestamp 1667941163
transform 1 0 16744 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_182
timestamp 1667941163
transform 1 0 17848 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1667941163
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1667941163
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1667941163
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1667941163
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1667941163
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1667941163
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1667941163
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1667941163
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1667941163
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1667941163
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1667941163
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_318
timestamp 1667941163
transform 1 0 30360 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_330
timestamp 1667941163
transform 1 0 31464 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_342
timestamp 1667941163
transform 1 0 32568 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_354
timestamp 1667941163
transform 1 0 33672 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_362
timestamp 1667941163
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1667941163
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1667941163
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_9
timestamp 1667941163
transform 1 0 1932 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1667941163
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_27
timestamp 1667941163
transform 1 0 3588 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_35
timestamp 1667941163
transform 1 0 4324 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_40
timestamp 1667941163
transform 1 0 4784 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_52
timestamp 1667941163
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1667941163
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1667941163
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1667941163
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1667941163
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1667941163
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_118
timestamp 1667941163
transform 1 0 11960 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_124
timestamp 1667941163
transform 1 0 12512 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_131
timestamp 1667941163
transform 1 0 13156 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_138
timestamp 1667941163
transform 1 0 13800 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_144
timestamp 1667941163
transform 1 0 14352 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_148
timestamp 1667941163
transform 1 0 14720 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_156
timestamp 1667941163
transform 1 0 15456 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_162
timestamp 1667941163
transform 1 0 16008 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1667941163
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1667941163
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1667941163
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1667941163
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1667941163
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1667941163
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1667941163
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1667941163
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1667941163
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1667941163
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1667941163
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1667941163
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1667941163
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1667941163
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1667941163
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1667941163
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1667941163
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1667941163
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1667941163
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1667941163
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1667941163
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1667941163
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_34
timestamp 1667941163
transform 1 0 4232 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_40
timestamp 1667941163
transform 1 0 4784 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_52
timestamp 1667941163
transform 1 0 5888 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_64
timestamp 1667941163
transform 1 0 6992 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_76
timestamp 1667941163
transform 1 0 8096 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_99
timestamp 1667941163
transform 1 0 10212 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_103
timestamp 1667941163
transform 1 0 10580 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_106
timestamp 1667941163
transform 1 0 10856 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_112
timestamp 1667941163
transform 1 0 11408 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_115
timestamp 1667941163
transform 1 0 11684 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_121
timestamp 1667941163
transform 1 0 12236 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_128
timestamp 1667941163
transform 1 0 12880 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_132
timestamp 1667941163
transform 1 0 13248 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1667941163
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_148
timestamp 1667941163
transform 1 0 14720 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_155
timestamp 1667941163
transform 1 0 15364 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_159
timestamp 1667941163
transform 1 0 15732 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_162
timestamp 1667941163
transform 1 0 16008 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_168
timestamp 1667941163
transform 1 0 16560 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_180
timestamp 1667941163
transform 1 0 17664 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_192
timestamp 1667941163
transform 1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1667941163
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1667941163
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1667941163
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1667941163
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1667941163
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1667941163
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1667941163
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1667941163
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1667941163
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1667941163
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1667941163
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1667941163
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1667941163
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1667941163
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1667941163
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1667941163
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1667941163
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_401
timestamp 1667941163
transform 1 0 37996 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_9
timestamp 1667941163
transform 1 0 1932 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_21
timestamp 1667941163
transform 1 0 3036 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_33
timestamp 1667941163
transform 1 0 4140 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_45
timestamp 1667941163
transform 1 0 5244 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1667941163
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1667941163
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_93
timestamp 1667941163
transform 1 0 9660 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_97
timestamp 1667941163
transform 1 0 10028 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_103
timestamp 1667941163
transform 1 0 10580 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1667941163
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_117
timestamp 1667941163
transform 1 0 11868 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_126
timestamp 1667941163
transform 1 0 12696 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_137
timestamp 1667941163
transform 1 0 13708 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_150
timestamp 1667941163
transform 1 0 14904 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_159
timestamp 1667941163
transform 1 0 15732 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1667941163
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_173
timestamp 1667941163
transform 1 0 17020 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_179
timestamp 1667941163
transform 1 0 17572 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_191
timestamp 1667941163
transform 1 0 18676 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_203
timestamp 1667941163
transform 1 0 19780 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_215
timestamp 1667941163
transform 1 0 20884 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1667941163
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1667941163
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1667941163
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1667941163
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1667941163
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1667941163
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1667941163
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1667941163
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1667941163
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1667941163
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1667941163
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1667941163
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1667941163
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1667941163
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1667941163
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1667941163
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1667941163
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1667941163
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1667941163
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1667941163
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1667941163
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_68
timestamp 1667941163
transform 1 0 7360 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_80
timestamp 1667941163
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_90
timestamp 1667941163
transform 1 0 9384 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_97
timestamp 1667941163
transform 1 0 10028 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_104
timestamp 1667941163
transform 1 0 10672 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_111
timestamp 1667941163
transform 1 0 11316 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_124
timestamp 1667941163
transform 1 0 12512 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_128
timestamp 1667941163
transform 1 0 12880 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1667941163
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_145
timestamp 1667941163
transform 1 0 14444 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_158
timestamp 1667941163
transform 1 0 15640 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_165
timestamp 1667941163
transform 1 0 16284 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_173
timestamp 1667941163
transform 1 0 17020 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_179
timestamp 1667941163
transform 1 0 17572 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_185
timestamp 1667941163
transform 1 0 18124 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_193
timestamp 1667941163
transform 1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1667941163
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_223
timestamp 1667941163
transform 1 0 21620 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_231
timestamp 1667941163
transform 1 0 22356 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_243
timestamp 1667941163
transform 1 0 23460 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1667941163
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1667941163
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1667941163
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1667941163
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1667941163
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1667941163
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1667941163
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1667941163
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1667941163
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1667941163
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1667941163
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1667941163
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_405
timestamp 1667941163
transform 1 0 38364 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_15
timestamp 1667941163
transform 1 0 2484 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_23
timestamp 1667941163
transform 1 0 3220 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_28
timestamp 1667941163
transform 1 0 3680 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_40
timestamp 1667941163
transform 1 0 4784 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_52
timestamp 1667941163
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1667941163
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_81
timestamp 1667941163
transform 1 0 8556 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_87
timestamp 1667941163
transform 1 0 9108 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_90
timestamp 1667941163
transform 1 0 9384 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_97
timestamp 1667941163
transform 1 0 10028 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1667941163
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_117
timestamp 1667941163
transform 1 0 11868 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_130
timestamp 1667941163
transform 1 0 13064 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_137
timestamp 1667941163
transform 1 0 13708 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_150
timestamp 1667941163
transform 1 0 14904 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_157
timestamp 1667941163
transform 1 0 15548 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1667941163
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_174
timestamp 1667941163
transform 1 0 17112 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_180
timestamp 1667941163
transform 1 0 17664 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_186
timestamp 1667941163
transform 1 0 18216 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_192
timestamp 1667941163
transform 1 0 18768 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_204
timestamp 1667941163
transform 1 0 19872 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_216
timestamp 1667941163
transform 1 0 20976 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1667941163
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1667941163
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1667941163
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1667941163
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1667941163
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1667941163
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1667941163
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1667941163
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1667941163
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1667941163
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1667941163
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1667941163
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1667941163
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1667941163
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_402
timestamp 1667941163
transform 1 0 38088 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_406
timestamp 1667941163
transform 1 0 38456 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_13
timestamp 1667941163
transform 1 0 2300 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_19
timestamp 1667941163
transform 1 0 2852 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_23
timestamp 1667941163
transform 1 0 3220 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1667941163
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_33
timestamp 1667941163
transform 1 0 4140 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_39
timestamp 1667941163
transform 1 0 4692 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_51
timestamp 1667941163
transform 1 0 5796 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_63
timestamp 1667941163
transform 1 0 6900 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_75
timestamp 1667941163
transform 1 0 8004 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_79
timestamp 1667941163
transform 1 0 8372 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1667941163
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_94
timestamp 1667941163
transform 1 0 9752 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_107
timestamp 1667941163
transform 1 0 10948 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_113
timestamp 1667941163
transform 1 0 11500 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_125
timestamp 1667941163
transform 1 0 12604 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1667941163
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_147
timestamp 1667941163
transform 1 0 14628 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_157
timestamp 1667941163
transform 1 0 15548 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_161
timestamp 1667941163
transform 1 0 15916 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_165
timestamp 1667941163
transform 1 0 16284 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_172
timestamp 1667941163
transform 1 0 16928 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_179
timestamp 1667941163
transform 1 0 17572 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_185
timestamp 1667941163
transform 1 0 18124 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_189
timestamp 1667941163
transform 1 0 18492 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1667941163
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_201
timestamp 1667941163
transform 1 0 19596 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_213
timestamp 1667941163
transform 1 0 20700 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_225
timestamp 1667941163
transform 1 0 21804 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_237
timestamp 1667941163
transform 1 0 22908 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_249
timestamp 1667941163
transform 1 0 24012 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1667941163
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1667941163
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1667941163
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1667941163
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1667941163
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1667941163
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1667941163
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1667941163
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1667941163
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1667941163
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1667941163
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_401
timestamp 1667941163
transform 1 0 37996 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_9
timestamp 1667941163
transform 1 0 1932 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_13
timestamp 1667941163
transform 1 0 2300 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_16
timestamp 1667941163
transform 1 0 2576 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_22
timestamp 1667941163
transform 1 0 3128 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_28
timestamp 1667941163
transform 1 0 3680 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_34
timestamp 1667941163
transform 1 0 4232 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_40
timestamp 1667941163
transform 1 0 4784 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_46
timestamp 1667941163
transform 1 0 5336 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1667941163
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_61
timestamp 1667941163
transform 1 0 6716 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_69
timestamp 1667941163
transform 1 0 7452 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_72
timestamp 1667941163
transform 1 0 7728 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_79
timestamp 1667941163
transform 1 0 8372 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_86
timestamp 1667941163
transform 1 0 9016 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_93
timestamp 1667941163
transform 1 0 9660 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1667941163
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_119
timestamp 1667941163
transform 1 0 12052 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_129
timestamp 1667941163
transform 1 0 12972 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_146
timestamp 1667941163
transform 1 0 14536 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_150
timestamp 1667941163
transform 1 0 14904 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_160
timestamp 1667941163
transform 1 0 15824 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1667941163
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_176
timestamp 1667941163
transform 1 0 17296 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_182
timestamp 1667941163
transform 1 0 17848 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_189
timestamp 1667941163
transform 1 0 18492 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_195
timestamp 1667941163
transform 1 0 19044 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_206
timestamp 1667941163
transform 1 0 20056 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_212
timestamp 1667941163
transform 1 0 20608 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1667941163
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1667941163
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1667941163
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1667941163
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1667941163
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1667941163
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1667941163
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1667941163
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1667941163
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1667941163
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1667941163
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1667941163
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1667941163
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1667941163
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1667941163
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_7
timestamp 1667941163
transform 1 0 1748 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_13
timestamp 1667941163
transform 1 0 2300 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_16
timestamp 1667941163
transform 1 0 2576 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1667941163
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_34
timestamp 1667941163
transform 1 0 4232 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_40
timestamp 1667941163
transform 1 0 4784 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_44
timestamp 1667941163
transform 1 0 5152 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_48
timestamp 1667941163
transform 1 0 5520 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_54
timestamp 1667941163
transform 1 0 6072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_60
timestamp 1667941163
transform 1 0 6624 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_66
timestamp 1667941163
transform 1 0 7176 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_69
timestamp 1667941163
transform 1 0 7452 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_75
timestamp 1667941163
transform 1 0 8004 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1667941163
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_89
timestamp 1667941163
transform 1 0 9292 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_96
timestamp 1667941163
transform 1 0 9936 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_103
timestamp 1667941163
transform 1 0 10580 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_116
timestamp 1667941163
transform 1 0 11776 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_120
timestamp 1667941163
transform 1 0 12144 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_124
timestamp 1667941163
transform 1 0 12512 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_137
timestamp 1667941163
transform 1 0 13708 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_145
timestamp 1667941163
transform 1 0 14444 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_155
timestamp 1667941163
transform 1 0 15364 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_159
timestamp 1667941163
transform 1 0 15732 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_164
timestamp 1667941163
transform 1 0 16192 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_36_175
timestamp 1667941163
transform 1 0 17204 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_36_190
timestamp 1667941163
transform 1 0 18584 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_201
timestamp 1667941163
transform 1 0 19596 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_207
timestamp 1667941163
transform 1 0 20148 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_213
timestamp 1667941163
transform 1 0 20700 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_220
timestamp 1667941163
transform 1 0 21344 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_226
timestamp 1667941163
transform 1 0 21896 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_238
timestamp 1667941163
transform 1 0 23000 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1667941163
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1667941163
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1667941163
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1667941163
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1667941163
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1667941163
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1667941163
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1667941163
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1667941163
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1667941163
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1667941163
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1667941163
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_389
timestamp 1667941163
transform 1 0 36892 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_397
timestamp 1667941163
transform 1 0 37628 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_402
timestamp 1667941163
transform 1 0 38088 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_406
timestamp 1667941163
transform 1 0 38456 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_9
timestamp 1667941163
transform 1 0 1932 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_16
timestamp 1667941163
transform 1 0 2576 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_22
timestamp 1667941163
transform 1 0 3128 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_28
timestamp 1667941163
transform 1 0 3680 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_31
timestamp 1667941163
transform 1 0 3956 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_39
timestamp 1667941163
transform 1 0 4692 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_42
timestamp 1667941163
transform 1 0 4968 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_48
timestamp 1667941163
transform 1 0 5520 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1667941163
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_61
timestamp 1667941163
transform 1 0 6716 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_64
timestamp 1667941163
transform 1 0 6992 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_68
timestamp 1667941163
transform 1 0 7360 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_71
timestamp 1667941163
transform 1 0 7636 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_77
timestamp 1667941163
transform 1 0 8188 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_84
timestamp 1667941163
transform 1 0 8832 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_91
timestamp 1667941163
transform 1 0 9476 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_98
timestamp 1667941163
transform 1 0 10120 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1667941163
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_124
timestamp 1667941163
transform 1 0 12512 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_128
timestamp 1667941163
transform 1 0 12880 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_132
timestamp 1667941163
transform 1 0 13248 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_145
timestamp 1667941163
transform 1 0 14444 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_158
timestamp 1667941163
transform 1 0 15640 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_165
timestamp 1667941163
transform 1 0 16284 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_173
timestamp 1667941163
transform 1 0 17020 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_180
timestamp 1667941163
transform 1 0 17664 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_187
timestamp 1667941163
transform 1 0 18308 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_191
timestamp 1667941163
transform 1 0 18676 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_201
timestamp 1667941163
transform 1 0 19596 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_214
timestamp 1667941163
transform 1 0 20792 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1667941163
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1667941163
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1667941163
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1667941163
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1667941163
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1667941163
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1667941163
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1667941163
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1667941163
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1667941163
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1667941163
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1667941163
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1667941163
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1667941163
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1667941163
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_401
timestamp 1667941163
transform 1 0 37996 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_404
timestamp 1667941163
transform 1 0 38272 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_7
timestamp 1667941163
transform 1 0 1748 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_13
timestamp 1667941163
transform 1 0 2300 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_19
timestamp 1667941163
transform 1 0 2852 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_25
timestamp 1667941163
transform 1 0 3404 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_33
timestamp 1667941163
transform 1 0 4140 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_36
timestamp 1667941163
transform 1 0 4416 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_40
timestamp 1667941163
transform 1 0 4784 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_43
timestamp 1667941163
transform 1 0 5060 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_49
timestamp 1667941163
transform 1 0 5612 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_53
timestamp 1667941163
transform 1 0 5980 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_56
timestamp 1667941163
transform 1 0 6256 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_62
timestamp 1667941163
transform 1 0 6808 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_65
timestamp 1667941163
transform 1 0 7084 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_73
timestamp 1667941163
transform 1 0 7820 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1667941163
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_98
timestamp 1667941163
transform 1 0 10120 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_111
timestamp 1667941163
transform 1 0 11316 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_124
timestamp 1667941163
transform 1 0 12512 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_130
timestamp 1667941163
transform 1 0 13064 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1667941163
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_152
timestamp 1667941163
transform 1 0 15088 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_159
timestamp 1667941163
transform 1 0 15732 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_166
timestamp 1667941163
transform 1 0 16376 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_179
timestamp 1667941163
transform 1 0 17572 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_186
timestamp 1667941163
transform 1 0 18216 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_193
timestamp 1667941163
transform 1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_202
timestamp 1667941163
transform 1 0 19688 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_209
timestamp 1667941163
transform 1 0 20332 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_213
timestamp 1667941163
transform 1 0 20700 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_218
timestamp 1667941163
transform 1 0 21160 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_224
timestamp 1667941163
transform 1 0 21712 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_236
timestamp 1667941163
transform 1 0 22816 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1667941163
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1667941163
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1667941163
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1667941163
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1667941163
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1667941163
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_316
timestamp 1667941163
transform 1 0 30176 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_322
timestamp 1667941163
transform 1 0 30728 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_334
timestamp 1667941163
transform 1 0 31832 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_346
timestamp 1667941163
transform 1 0 32936 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_358
timestamp 1667941163
transform 1 0 34040 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1667941163
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1667941163
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 1667941163
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_10
timestamp 1667941163
transform 1 0 2024 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_16
timestamp 1667941163
transform 1 0 2576 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_22
timestamp 1667941163
transform 1 0 3128 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_32
timestamp 1667941163
transform 1 0 4048 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_36
timestamp 1667941163
transform 1 0 4416 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_39
timestamp 1667941163
transform 1 0 4692 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_43
timestamp 1667941163
transform 1 0 5060 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_46
timestamp 1667941163
transform 1 0 5336 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1667941163
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_62
timestamp 1667941163
transform 1 0 6808 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_68
timestamp 1667941163
transform 1 0 7360 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_75
timestamp 1667941163
transform 1 0 8004 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_82
timestamp 1667941163
transform 1 0 8648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_89
timestamp 1667941163
transform 1 0 9292 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_96
timestamp 1667941163
transform 1 0 9936 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_103
timestamp 1667941163
transform 1 0 10580 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1667941163
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_120
timestamp 1667941163
transform 1 0 12144 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_133
timestamp 1667941163
transform 1 0 13340 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_146
timestamp 1667941163
transform 1 0 14536 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_152
timestamp 1667941163
transform 1 0 15088 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1667941163
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_184
timestamp 1667941163
transform 1 0 18032 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_197
timestamp 1667941163
transform 1 0 19228 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_204
timestamp 1667941163
transform 1 0 19872 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_214
timestamp 1667941163
transform 1 0 20792 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1667941163
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_229
timestamp 1667941163
transform 1 0 22172 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_241
timestamp 1667941163
transform 1 0 23276 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_253
timestamp 1667941163
transform 1 0 24380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_265
timestamp 1667941163
transform 1 0 25484 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_271
timestamp 1667941163
transform 1 0 26036 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_275
timestamp 1667941163
transform 1 0 26404 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1667941163
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_285
timestamp 1667941163
transform 1 0 27324 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_297
timestamp 1667941163
transform 1 0 28428 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_309
timestamp 1667941163
transform 1 0 29532 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_316
timestamp 1667941163
transform 1 0 30176 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_322
timestamp 1667941163
transform 1 0 30728 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_334
timestamp 1667941163
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1667941163
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1667941163
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1667941163
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1667941163
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1667941163
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_7
timestamp 1667941163
transform 1 0 1748 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_13
timestamp 1667941163
transform 1 0 2300 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_19
timestamp 1667941163
transform 1 0 2852 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_25
timestamp 1667941163
transform 1 0 3404 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_33
timestamp 1667941163
transform 1 0 4140 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_36
timestamp 1667941163
transform 1 0 4416 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_40
timestamp 1667941163
transform 1 0 4784 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_43
timestamp 1667941163
transform 1 0 5060 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_49
timestamp 1667941163
transform 1 0 5612 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_55
timestamp 1667941163
transform 1 0 6164 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_61
timestamp 1667941163
transform 1 0 6716 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_68
timestamp 1667941163
transform 1 0 7360 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_75
timestamp 1667941163
transform 1 0 8004 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1667941163
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_91
timestamp 1667941163
transform 1 0 9476 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_104
timestamp 1667941163
transform 1 0 10672 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_111
timestamp 1667941163
transform 1 0 11316 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_124
timestamp 1667941163
transform 1 0 12512 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_128
timestamp 1667941163
transform 1 0 12880 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1667941163
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_156
timestamp 1667941163
transform 1 0 15456 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_164
timestamp 1667941163
transform 1 0 16192 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_178
timestamp 1667941163
transform 1 0 17480 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_184
timestamp 1667941163
transform 1 0 18032 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1667941163
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_201
timestamp 1667941163
transform 1 0 19596 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_208
timestamp 1667941163
transform 1 0 20240 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_215
timestamp 1667941163
transform 1 0 20884 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_221
timestamp 1667941163
transform 1 0 21436 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_234
timestamp 1667941163
transform 1 0 22632 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_240
timestamp 1667941163
transform 1 0 23184 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1667941163
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1667941163
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1667941163
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1667941163
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1667941163
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1667941163
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1667941163
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_345
timestamp 1667941163
transform 1 0 32844 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_356
timestamp 1667941163
transform 1 0 33856 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_362
timestamp 1667941163
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1667941163
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_389
timestamp 1667941163
transform 1 0 36892 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_397
timestamp 1667941163
transform 1 0 37628 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_402
timestamp 1667941163
transform 1 0 38088 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_406
timestamp 1667941163
transform 1 0 38456 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_8
timestamp 1667941163
transform 1 0 1840 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_14
timestamp 1667941163
transform 1 0 2392 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_20
timestamp 1667941163
transform 1 0 2944 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_24
timestamp 1667941163
transform 1 0 3312 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_27
timestamp 1667941163
transform 1 0 3588 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_31
timestamp 1667941163
transform 1 0 3956 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_34
timestamp 1667941163
transform 1 0 4232 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_40
timestamp 1667941163
transform 1 0 4784 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_46
timestamp 1667941163
transform 1 0 5336 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_53
timestamp 1667941163
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_62
timestamp 1667941163
transform 1 0 6808 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_66
timestamp 1667941163
transform 1 0 7176 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_69
timestamp 1667941163
transform 1 0 7452 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_76
timestamp 1667941163
transform 1 0 8096 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_83
timestamp 1667941163
transform 1 0 8740 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_90
timestamp 1667941163
transform 1 0 9384 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_97
timestamp 1667941163
transform 1 0 10028 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1667941163
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_124
timestamp 1667941163
transform 1 0 12512 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_137
timestamp 1667941163
transform 1 0 13708 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_41_156
timestamp 1667941163
transform 1 0 15456 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_162
timestamp 1667941163
transform 1 0 16008 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1667941163
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_175
timestamp 1667941163
transform 1 0 17204 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_182
timestamp 1667941163
transform 1 0 17848 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_189
timestamp 1667941163
transform 1 0 18492 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_202
timestamp 1667941163
transform 1 0 19688 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_215
timestamp 1667941163
transform 1 0 20884 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1667941163
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_230
timestamp 1667941163
transform 1 0 22264 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_236
timestamp 1667941163
transform 1 0 22816 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_242
timestamp 1667941163
transform 1 0 23368 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_248
timestamp 1667941163
transform 1 0 23920 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_260
timestamp 1667941163
transform 1 0 25024 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_272
timestamp 1667941163
transform 1 0 26128 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1667941163
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_305
timestamp 1667941163
transform 1 0 29164 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_312
timestamp 1667941163
transform 1 0 29808 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_324
timestamp 1667941163
transform 1 0 30912 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1667941163
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1667941163
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1667941163
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1667941163
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1667941163
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_8
timestamp 1667941163
transform 1 0 1840 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_14
timestamp 1667941163
transform 1 0 2392 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_20
timestamp 1667941163
transform 1 0 2944 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_26
timestamp 1667941163
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_35
timestamp 1667941163
transform 1 0 4324 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_38
timestamp 1667941163
transform 1 0 4600 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_44
timestamp 1667941163
transform 1 0 5152 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_50
timestamp 1667941163
transform 1 0 5704 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_56
timestamp 1667941163
transform 1 0 6256 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_62
timestamp 1667941163
transform 1 0 6808 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_69
timestamp 1667941163
transform 1 0 7452 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_75
timestamp 1667941163
transform 1 0 8004 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1667941163
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_91
timestamp 1667941163
transform 1 0 9476 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_104
timestamp 1667941163
transform 1 0 10672 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_121
timestamp 1667941163
transform 1 0 12236 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1667941163
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_147
timestamp 1667941163
transform 1 0 14628 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_162
timestamp 1667941163
transform 1 0 16008 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_175
timestamp 1667941163
transform 1 0 17204 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1667941163
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_202
timestamp 1667941163
transform 1 0 19688 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_206
timestamp 1667941163
transform 1 0 20056 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_216
timestamp 1667941163
transform 1 0 20976 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_223
timestamp 1667941163
transform 1 0 21620 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_229
timestamp 1667941163
transform 1 0 22172 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1667941163
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1667941163
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1667941163
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1667941163
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1667941163
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1667941163
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_314
timestamp 1667941163
transform 1 0 29992 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_326
timestamp 1667941163
transform 1 0 31096 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_338
timestamp 1667941163
transform 1 0 32200 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_350
timestamp 1667941163
transform 1 0 33304 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_362
timestamp 1667941163
transform 1 0 34408 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1667941163
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_401
timestamp 1667941163
transform 1 0 37996 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_405
timestamp 1667941163
transform 1 0 38364 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_7
timestamp 1667941163
transform 1 0 1748 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_11
timestamp 1667941163
transform 1 0 2116 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_18
timestamp 1667941163
transform 1 0 2760 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_26
timestamp 1667941163
transform 1 0 3496 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_29
timestamp 1667941163
transform 1 0 3772 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_35
timestamp 1667941163
transform 1 0 4324 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_41
timestamp 1667941163
transform 1 0 4876 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_47
timestamp 1667941163
transform 1 0 5428 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_54
timestamp 1667941163
transform 1 0 6072 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_61
timestamp 1667941163
transform 1 0 6716 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_68
timestamp 1667941163
transform 1 0 7360 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_75
timestamp 1667941163
transform 1 0 8004 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_82
timestamp 1667941163
transform 1 0 8648 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_95
timestamp 1667941163
transform 1 0 9844 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1667941163
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_118
timestamp 1667941163
transform 1 0 11960 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_131
timestamp 1667941163
transform 1 0 13156 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_144
timestamp 1667941163
transform 1 0 14352 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_157
timestamp 1667941163
transform 1 0 15548 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_43_166
timestamp 1667941163
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_173
timestamp 1667941163
transform 1 0 17020 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_177
timestamp 1667941163
transform 1 0 17388 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_184
timestamp 1667941163
transform 1 0 18032 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_191
timestamp 1667941163
transform 1 0 18676 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_208
timestamp 1667941163
transform 1 0 20240 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_215
timestamp 1667941163
transform 1 0 20884 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1667941163
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_236
timestamp 1667941163
transform 1 0 22816 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_243
timestamp 1667941163
transform 1 0 23460 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1667941163
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1667941163
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1667941163
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1667941163
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1667941163
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1667941163
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1667941163
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1667941163
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1667941163
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1667941163
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1667941163
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1667941163
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1667941163
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1667941163
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_7
timestamp 1667941163
transform 1 0 1748 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_11
timestamp 1667941163
transform 1 0 2116 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_18
timestamp 1667941163
transform 1 0 2760 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_25
timestamp 1667941163
transform 1 0 3404 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_37
timestamp 1667941163
transform 1 0 4508 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_43
timestamp 1667941163
transform 1 0 5060 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_49
timestamp 1667941163
transform 1 0 5612 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_55
timestamp 1667941163
transform 1 0 6164 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_61
timestamp 1667941163
transform 1 0 6716 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_68
timestamp 1667941163
transform 1 0 7360 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_75
timestamp 1667941163
transform 1 0 8004 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_82
timestamp 1667941163
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_100
timestamp 1667941163
transform 1 0 10304 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_106
timestamp 1667941163
transform 1 0 10856 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_119
timestamp 1667941163
transform 1 0 12052 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_125
timestamp 1667941163
transform 1 0 12604 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1667941163
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_146
timestamp 1667941163
transform 1 0 14536 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_159
timestamp 1667941163
transform 1 0 15732 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_166
timestamp 1667941163
transform 1 0 16376 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_179
timestamp 1667941163
transform 1 0 17572 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_185
timestamp 1667941163
transform 1 0 18124 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_193
timestamp 1667941163
transform 1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_208
timestamp 1667941163
transform 1 0 20240 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_214
timestamp 1667941163
transform 1 0 20792 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_224
timestamp 1667941163
transform 1 0 21712 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_232
timestamp 1667941163
transform 1 0 22448 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_236
timestamp 1667941163
transform 1 0 22816 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_243
timestamp 1667941163
transform 1 0 23460 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_249
timestamp 1667941163
transform 1 0 24012 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_257
timestamp 1667941163
transform 1 0 24748 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_269
timestamp 1667941163
transform 1 0 25852 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_281
timestamp 1667941163
transform 1 0 26956 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_293
timestamp 1667941163
transform 1 0 28060 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_305
timestamp 1667941163
transform 1 0 29164 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_314
timestamp 1667941163
transform 1 0 29992 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_326
timestamp 1667941163
transform 1 0 31096 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_338
timestamp 1667941163
transform 1 0 32200 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_350
timestamp 1667941163
transform 1 0 33304 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_362
timestamp 1667941163
transform 1 0 34408 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1667941163
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1667941163
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_401
timestamp 1667941163
transform 1 0 37996 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_9
timestamp 1667941163
transform 1 0 1932 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_16
timestamp 1667941163
transform 1 0 2576 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_23
timestamp 1667941163
transform 1 0 3220 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_30
timestamp 1667941163
transform 1 0 3864 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_36
timestamp 1667941163
transform 1 0 4416 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_42
timestamp 1667941163
transform 1 0 4968 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_48
timestamp 1667941163
transform 1 0 5520 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1667941163
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_61
timestamp 1667941163
transform 1 0 6716 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_64
timestamp 1667941163
transform 1 0 6992 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_70
timestamp 1667941163
transform 1 0 7544 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_77
timestamp 1667941163
transform 1 0 8188 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_94
timestamp 1667941163
transform 1 0 9752 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_103
timestamp 1667941163
transform 1 0 10580 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1667941163
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_126
timestamp 1667941163
transform 1 0 12696 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_130
timestamp 1667941163
transform 1 0 13064 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_140
timestamp 1667941163
transform 1 0 13984 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_153
timestamp 1667941163
transform 1 0 15180 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1667941163
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_182
timestamp 1667941163
transform 1 0 17848 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_197
timestamp 1667941163
transform 1 0 19228 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_210
timestamp 1667941163
transform 1 0 20424 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_221
timestamp 1667941163
transform 1 0 21436 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_236
timestamp 1667941163
transform 1 0 22816 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1667941163
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1667941163
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1667941163
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1667941163
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1667941163
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1667941163
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1667941163
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1667941163
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1667941163
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1667941163
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1667941163
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1667941163
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1667941163
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1667941163
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1667941163
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_9
timestamp 1667941163
transform 1 0 1932 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_13
timestamp 1667941163
transform 1 0 2300 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_20
timestamp 1667941163
transform 1 0 2944 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_26
timestamp 1667941163
transform 1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_34
timestamp 1667941163
transform 1 0 4232 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_49
timestamp 1667941163
transform 1 0 5612 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_52
timestamp 1667941163
transform 1 0 5888 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_58
timestamp 1667941163
transform 1 0 6440 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_64
timestamp 1667941163
transform 1 0 6992 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_70
timestamp 1667941163
transform 1 0 7544 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_76
timestamp 1667941163
transform 1 0 8096 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_82
timestamp 1667941163
transform 1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_92
timestamp 1667941163
transform 1 0 9568 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_105
timestamp 1667941163
transform 1 0 10764 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_118
timestamp 1667941163
transform 1 0 11960 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_124
timestamp 1667941163
transform 1 0 12512 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_131
timestamp 1667941163
transform 1 0 13156 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1667941163
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_156
timestamp 1667941163
transform 1 0 15456 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_164
timestamp 1667941163
transform 1 0 16192 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_168
timestamp 1667941163
transform 1 0 16560 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_181
timestamp 1667941163
transform 1 0 17756 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1667941163
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_202
timestamp 1667941163
transform 1 0 19688 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_219
timestamp 1667941163
transform 1 0 21252 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_226
timestamp 1667941163
transform 1 0 21896 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_232
timestamp 1667941163
transform 1 0 22448 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_238
timestamp 1667941163
transform 1 0 23000 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_244
timestamp 1667941163
transform 1 0 23552 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_250
timestamp 1667941163
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1667941163
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1667941163
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1667941163
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1667941163
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1667941163
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1667941163
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1667941163
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1667941163
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1667941163
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1667941163
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1667941163
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_401
timestamp 1667941163
transform 1 0 37996 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_9
timestamp 1667941163
transform 1 0 1932 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_16
timestamp 1667941163
transform 1 0 2576 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_23
timestamp 1667941163
transform 1 0 3220 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_30
timestamp 1667941163
transform 1 0 3864 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_37
timestamp 1667941163
transform 1 0 4508 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_44
timestamp 1667941163
transform 1 0 5152 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_50
timestamp 1667941163
transform 1 0 5704 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_54
timestamp 1667941163
transform 1 0 6072 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_61
timestamp 1667941163
transform 1 0 6716 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_65
timestamp 1667941163
transform 1 0 7084 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_72
timestamp 1667941163
transform 1 0 7728 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_82
timestamp 1667941163
transform 1 0 8648 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_106
timestamp 1667941163
transform 1 0 10856 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_124
timestamp 1667941163
transform 1 0 12512 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_137
timestamp 1667941163
transform 1 0 13708 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_47_154
timestamp 1667941163
transform 1 0 15272 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_162
timestamp 1667941163
transform 1 0 16008 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_166
timestamp 1667941163
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_180
timestamp 1667941163
transform 1 0 17664 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_195
timestamp 1667941163
transform 1 0 19044 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_202
timestamp 1667941163
transform 1 0 19688 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_209
timestamp 1667941163
transform 1 0 20332 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_216
timestamp 1667941163
transform 1 0 20976 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1667941163
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_230
timestamp 1667941163
transform 1 0 22264 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_236
timestamp 1667941163
transform 1 0 22816 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_242
timestamp 1667941163
transform 1 0 23368 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_248
timestamp 1667941163
transform 1 0 23920 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_260
timestamp 1667941163
transform 1 0 25024 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_272
timestamp 1667941163
transform 1 0 26128 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1667941163
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1667941163
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1667941163
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1667941163
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1667941163
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1667941163
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1667941163
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1667941163
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1667941163
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1667941163
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1667941163
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_7
timestamp 1667941163
transform 1 0 1748 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_14
timestamp 1667941163
transform 1 0 2392 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_21
timestamp 1667941163
transform 1 0 3036 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_34
timestamp 1667941163
transform 1 0 4232 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_41
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_48
timestamp 1667941163
transform 1 0 5520 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_55
timestamp 1667941163
transform 1 0 6164 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_48_66
timestamp 1667941163
transform 1 0 7176 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_75
timestamp 1667941163
transform 1 0 8004 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_82
timestamp 1667941163
transform 1 0 8648 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_91
timestamp 1667941163
transform 1 0 9476 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_95
timestamp 1667941163
transform 1 0 9844 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_120
timestamp 1667941163
transform 1 0 12144 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_131
timestamp 1667941163
transform 1 0 13156 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_138
timestamp 1667941163
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_145
timestamp 1667941163
transform 1 0 14444 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_158
timestamp 1667941163
transform 1 0 15640 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_171
timestamp 1667941163
transform 1 0 16836 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_184
timestamp 1667941163
transform 1 0 18032 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_191
timestamp 1667941163
transform 1 0 18676 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1667941163
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_202
timestamp 1667941163
transform 1 0 19688 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_208
timestamp 1667941163
transform 1 0 20240 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_212
timestamp 1667941163
transform 1 0 20608 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_219
timestamp 1667941163
transform 1 0 21252 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_225
timestamp 1667941163
transform 1 0 21804 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_231
timestamp 1667941163
transform 1 0 22356 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_237
timestamp 1667941163
transform 1 0 22908 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_243
timestamp 1667941163
transform 1 0 23460 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1667941163
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1667941163
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1667941163
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1667941163
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1667941163
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1667941163
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1667941163
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1667941163
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1667941163
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1667941163
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1667941163
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1667941163
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_401
timestamp 1667941163
transform 1 0 37996 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_405
timestamp 1667941163
transform 1 0 38364 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_7
timestamp 1667941163
transform 1 0 1748 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_14
timestamp 1667941163
transform 1 0 2392 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_22
timestamp 1667941163
transform 1 0 3128 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_43
timestamp 1667941163
transform 1 0 5060 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_54
timestamp 1667941163
transform 1 0 6072 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_62
timestamp 1667941163
transform 1 0 6808 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_69
timestamp 1667941163
transform 1 0 7452 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_76
timestamp 1667941163
transform 1 0 8096 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_101
timestamp 1667941163
transform 1 0 10396 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_110
timestamp 1667941163
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_120
timestamp 1667941163
transform 1 0 12144 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_127
timestamp 1667941163
transform 1 0 12788 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_140
timestamp 1667941163
transform 1 0 13984 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_153
timestamp 1667941163
transform 1 0 15180 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_166
timestamp 1667941163
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_174
timestamp 1667941163
transform 1 0 17112 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_187
timestamp 1667941163
transform 1 0 18308 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_200
timestamp 1667941163
transform 1 0 19504 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_213
timestamp 1667941163
transform 1 0 20700 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_220
timestamp 1667941163
transform 1 0 21344 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_230
timestamp 1667941163
transform 1 0 22264 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_236
timestamp 1667941163
transform 1 0 22816 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_243
timestamp 1667941163
transform 1 0 23460 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1667941163
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1667941163
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1667941163
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1667941163
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1667941163
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_305
timestamp 1667941163
transform 1 0 29164 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_313
timestamp 1667941163
transform 1 0 29900 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_318
timestamp 1667941163
transform 1 0 30360 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_330
timestamp 1667941163
transform 1 0 31464 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1667941163
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1667941163
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1667941163
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_26
timestamp 1667941163
transform 1 0 3496 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_51
timestamp 1667941163
transform 1 0 5796 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_59
timestamp 1667941163
transform 1 0 6532 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_63
timestamp 1667941163
transform 1 0 6900 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_70
timestamp 1667941163
transform 1 0 7544 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1667941163
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1667941163
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_92
timestamp 1667941163
transform 1 0 9568 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_119
timestamp 1667941163
transform 1 0 12052 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_50_134
timestamp 1667941163
transform 1 0 13432 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_152
timestamp 1667941163
transform 1 0 15088 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_156
timestamp 1667941163
transform 1 0 15456 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_166
timestamp 1667941163
transform 1 0 16376 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_181
timestamp 1667941163
transform 1 0 17756 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1667941163
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_212
timestamp 1667941163
transform 1 0 20608 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_219
timestamp 1667941163
transform 1 0 21252 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_226
timestamp 1667941163
transform 1 0 21896 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_232
timestamp 1667941163
transform 1 0 22448 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_244
timestamp 1667941163
transform 1 0 23552 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1667941163
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1667941163
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1667941163
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1667941163
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1667941163
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1667941163
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1667941163
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1667941163
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1667941163
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1667941163
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1667941163
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1667941163
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_401
timestamp 1667941163
transform 1 0 37996 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_405
timestamp 1667941163
transform 1 0 38364 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_9
timestamp 1667941163
transform 1 0 1932 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_30
timestamp 1667941163
transform 1 0 3864 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_54
timestamp 1667941163
transform 1 0 6072 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_63
timestamp 1667941163
transform 1 0 6900 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_87
timestamp 1667941163
transform 1 0 9108 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_96
timestamp 1667941163
transform 1 0 9936 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_103
timestamp 1667941163
transform 1 0 10580 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1667941163
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_136
timestamp 1667941163
transform 1 0 13616 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_142
timestamp 1667941163
transform 1 0 14168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_146
timestamp 1667941163
transform 1 0 14536 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_159
timestamp 1667941163
transform 1 0 15732 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1667941163
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_184
timestamp 1667941163
transform 1 0 18032 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_190
timestamp 1667941163
transform 1 0 18584 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_203
timestamp 1667941163
transform 1 0 19780 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_216
timestamp 1667941163
transform 1 0 20976 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1667941163
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_229
timestamp 1667941163
transform 1 0 22172 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_235
timestamp 1667941163
transform 1 0 22724 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_247
timestamp 1667941163
transform 1 0 23828 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_259
timestamp 1667941163
transform 1 0 24932 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_271
timestamp 1667941163
transform 1 0 26036 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1667941163
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1667941163
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1667941163
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1667941163
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1667941163
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1667941163
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1667941163
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1667941163
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1667941163
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1667941163
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1667941163
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_9
timestamp 1667941163
transform 1 0 1932 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_16
timestamp 1667941163
transform 1 0 2576 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_22
timestamp 1667941163
transform 1 0 3128 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_26
timestamp 1667941163
transform 1 0 3496 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_51
timestamp 1667941163
transform 1 0 5796 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_82
timestamp 1667941163
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_91
timestamp 1667941163
transform 1 0 9476 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_95
timestamp 1667941163
transform 1 0 9844 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_122
timestamp 1667941163
transform 1 0 12328 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_131
timestamp 1667941163
transform 1 0 13156 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1667941163
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_150
timestamp 1667941163
transform 1 0 14904 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_163
timestamp 1667941163
transform 1 0 16100 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_170
timestamp 1667941163
transform 1 0 16744 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_183
timestamp 1667941163
transform 1 0 17940 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_190
timestamp 1667941163
transform 1 0 18584 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_208
timestamp 1667941163
transform 1 0 20240 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_215
timestamp 1667941163
transform 1 0 20884 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_221
timestamp 1667941163
transform 1 0 21436 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_227
timestamp 1667941163
transform 1 0 21988 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_233
timestamp 1667941163
transform 1 0 22540 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_239
timestamp 1667941163
transform 1 0 23092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1667941163
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1667941163
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1667941163
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1667941163
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1667941163
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1667941163
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1667941163
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1667941163
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1667941163
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1667941163
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1667941163
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1667941163
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1667941163
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_401
timestamp 1667941163
transform 1 0 37996 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_9
timestamp 1667941163
transform 1 0 1932 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_17
timestamp 1667941163
transform 1 0 2668 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_23
timestamp 1667941163
transform 1 0 3220 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_27
timestamp 1667941163
transform 1 0 3588 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1667941163
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1667941163
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_83
timestamp 1667941163
transform 1 0 8740 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 1667941163
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_138
timestamp 1667941163
transform 1 0 13800 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_53_153
timestamp 1667941163
transform 1 0 15180 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_53_162
timestamp 1667941163
transform 1 0 16008 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_184
timestamp 1667941163
transform 1 0 18032 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_191
timestamp 1667941163
transform 1 0 18676 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_204
timestamp 1667941163
transform 1 0 19872 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_211
timestamp 1667941163
transform 1 0 20516 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_218
timestamp 1667941163
transform 1 0 21160 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_229
timestamp 1667941163
transform 1 0 22172 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_235
timestamp 1667941163
transform 1 0 22724 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_241
timestamp 1667941163
transform 1 0 23276 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_253
timestamp 1667941163
transform 1 0 24380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_265
timestamp 1667941163
transform 1 0 25484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_277
timestamp 1667941163
transform 1 0 26588 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1667941163
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1667941163
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1667941163
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1667941163
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1667941163
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1667941163
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1667941163
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1667941163
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1667941163
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1667941163
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1667941163
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_9
timestamp 1667941163
transform 1 0 1932 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_20
timestamp 1667941163
transform 1 0 2944 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_26
timestamp 1667941163
transform 1 0 3496 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_51
timestamp 1667941163
transform 1 0 5796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_57
timestamp 1667941163
transform 1 0 6348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_81
timestamp 1667941163
transform 1 0 8556 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_89
timestamp 1667941163
transform 1 0 9292 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_111
timestamp 1667941163
transform 1 0 11316 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_117
timestamp 1667941163
transform 1 0 11868 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_124
timestamp 1667941163
transform 1 0 12512 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_131
timestamp 1667941163
transform 1 0 13156 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_138
timestamp 1667941163
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_145
timestamp 1667941163
transform 1 0 14444 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_149
timestamp 1667941163
transform 1 0 14812 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_162
timestamp 1667941163
transform 1 0 16008 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_173
timestamp 1667941163
transform 1 0 17020 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_190
timestamp 1667941163
transform 1 0 18584 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_208
timestamp 1667941163
transform 1 0 20240 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_215
timestamp 1667941163
transform 1 0 20884 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_221
timestamp 1667941163
transform 1 0 21436 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_227
timestamp 1667941163
transform 1 0 21988 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_233
timestamp 1667941163
transform 1 0 22540 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_239
timestamp 1667941163
transform 1 0 23092 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1667941163
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1667941163
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1667941163
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1667941163
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1667941163
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1667941163
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1667941163
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1667941163
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1667941163
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1667941163
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1667941163
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1667941163
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_401
timestamp 1667941163
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_27
timestamp 1667941163
transform 1 0 3588 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_54
timestamp 1667941163
transform 1 0 6072 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_82
timestamp 1667941163
transform 1 0 8648 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_88
timestamp 1667941163
transform 1 0 9200 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_110
timestamp 1667941163
transform 1 0 11224 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_135
timestamp 1667941163
transform 1 0 13524 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_148
timestamp 1667941163
transform 1 0 14720 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_163
timestamp 1667941163
transform 1 0 16100 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1667941163
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_176
timestamp 1667941163
transform 1 0 17296 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_189
timestamp 1667941163
transform 1 0 18492 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_198
timestamp 1667941163
transform 1 0 19320 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_205
timestamp 1667941163
transform 1 0 19964 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_212
timestamp 1667941163
transform 1 0 20608 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_219
timestamp 1667941163
transform 1 0 21252 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1667941163
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_229
timestamp 1667941163
transform 1 0 22172 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_235
timestamp 1667941163
transform 1 0 22724 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_241
timestamp 1667941163
transform 1 0 23276 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_247
timestamp 1667941163
transform 1 0 23828 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_253
timestamp 1667941163
transform 1 0 24380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_265
timestamp 1667941163
transform 1 0 25484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_277
timestamp 1667941163
transform 1 0 26588 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1667941163
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1667941163
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1667941163
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1667941163
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1667941163
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1667941163
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1667941163
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1667941163
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1667941163
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_397
timestamp 1667941163
transform 1 0 37628 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1667941163
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_26
timestamp 1667941163
transform 1 0 3496 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_35
timestamp 1667941163
transform 1 0 4324 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_43
timestamp 1667941163
transform 1 0 5060 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_74
timestamp 1667941163
transform 1 0 7912 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_56_81
timestamp 1667941163
transform 1 0 8556 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_91
timestamp 1667941163
transform 1 0 9476 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_95
timestamp 1667941163
transform 1 0 9844 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_102
timestamp 1667941163
transform 1 0 10488 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_129
timestamp 1667941163
transform 1 0 12972 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_138
timestamp 1667941163
transform 1 0 13800 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_148
timestamp 1667941163
transform 1 0 14720 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_155
timestamp 1667941163
transform 1 0 15364 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_159
timestamp 1667941163
transform 1 0 15732 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_169
timestamp 1667941163
transform 1 0 16652 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_179
timestamp 1667941163
transform 1 0 17572 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_186
timestamp 1667941163
transform 1 0 18216 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_56_193
timestamp 1667941163
transform 1 0 18860 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_202
timestamp 1667941163
transform 1 0 19688 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_209
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_216
timestamp 1667941163
transform 1 0 20976 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_222
timestamp 1667941163
transform 1 0 21528 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_228
timestamp 1667941163
transform 1 0 22080 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_234
timestamp 1667941163
transform 1 0 22632 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_240
timestamp 1667941163
transform 1 0 23184 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_246
timestamp 1667941163
transform 1 0 23736 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_257
timestamp 1667941163
transform 1 0 24748 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_269
timestamp 1667941163
transform 1 0 25852 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_281
timestamp 1667941163
transform 1 0 26956 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_293
timestamp 1667941163
transform 1 0 28060 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_305
timestamp 1667941163
transform 1 0 29164 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1667941163
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1667941163
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1667941163
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1667941163
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1667941163
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_401
timestamp 1667941163
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_27
timestamp 1667941163
transform 1 0 3588 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_54
timestamp 1667941163
transform 1 0 6072 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_61
timestamp 1667941163
transform 1 0 6716 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_83
timestamp 1667941163
transform 1 0 8740 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_110
timestamp 1667941163
transform 1 0 11224 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_138
timestamp 1667941163
transform 1 0 13800 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_146
timestamp 1667941163
transform 1 0 14536 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_150
timestamp 1667941163
transform 1 0 14904 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_156
timestamp 1667941163
transform 1 0 15456 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_166
timestamp 1667941163
transform 1 0 16376 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_177
timestamp 1667941163
transform 1 0 17388 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_181
timestamp 1667941163
transform 1 0 17756 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_195
timestamp 1667941163
transform 1 0 19044 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_208
timestamp 1667941163
transform 1 0 20240 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_214
timestamp 1667941163
transform 1 0 20792 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_220
timestamp 1667941163
transform 1 0 21344 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_229
timestamp 1667941163
transform 1 0 22172 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_235
timestamp 1667941163
transform 1 0 22724 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_241
timestamp 1667941163
transform 1 0 23276 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_247
timestamp 1667941163
transform 1 0 23828 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_253
timestamp 1667941163
transform 1 0 24380 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_259
timestamp 1667941163
transform 1 0 24932 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_271
timestamp 1667941163
transform 1 0 26036 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1667941163
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1667941163
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1667941163
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1667941163
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1667941163
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1667941163
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1667941163
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1667941163
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_397
timestamp 1667941163
transform 1 0 37628 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_26
timestamp 1667941163
transform 1 0 3496 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_51
timestamp 1667941163
transform 1 0 5796 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_55
timestamp 1667941163
transform 1 0 6164 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_79
timestamp 1667941163
transform 1 0 8372 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1667941163
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_110
timestamp 1667941163
transform 1 0 11224 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_135
timestamp 1667941163
transform 1 0 13524 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1667941163
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_158
timestamp 1667941163
transform 1 0 15640 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_164
timestamp 1667941163
transform 1 0 16192 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_171
timestamp 1667941163
transform 1 0 16836 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_181
timestamp 1667941163
transform 1 0 17756 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_191
timestamp 1667941163
transform 1 0 18676 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1667941163
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_202
timestamp 1667941163
transform 1 0 19688 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_215
timestamp 1667941163
transform 1 0 20884 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_227
timestamp 1667941163
transform 1 0 21988 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_233
timestamp 1667941163
transform 1 0 22540 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_239
timestamp 1667941163
transform 1 0 23092 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1667941163
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1667941163
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_257
timestamp 1667941163
transform 1 0 24748 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_269
timestamp 1667941163
transform 1 0 25852 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_281
timestamp 1667941163
transform 1 0 26956 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_293
timestamp 1667941163
transform 1 0 28060 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_305
timestamp 1667941163
transform 1 0 29164 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1667941163
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1667941163
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1667941163
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1667941163
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1667941163
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1667941163
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1667941163
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 1667941163
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_27
timestamp 1667941163
transform 1 0 3588 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1667941163
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1667941163
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_81
timestamp 1667941163
transform 1 0 8556 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_108
timestamp 1667941163
transform 1 0 11040 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_135
timestamp 1667941163
transform 1 0 13524 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_152
timestamp 1667941163
transform 1 0 15088 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_159
timestamp 1667941163
transform 1 0 15732 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_166
timestamp 1667941163
transform 1 0 16376 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_177
timestamp 1667941163
transform 1 0 17388 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_184
timestamp 1667941163
transform 1 0 18032 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_191
timestamp 1667941163
transform 1 0 18676 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_198
timestamp 1667941163
transform 1 0 19320 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_204
timestamp 1667941163
transform 1 0 19872 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_210
timestamp 1667941163
transform 1 0 20424 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_216
timestamp 1667941163
transform 1 0 20976 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_222
timestamp 1667941163
transform 1 0 21528 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_229
timestamp 1667941163
transform 1 0 22172 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_235
timestamp 1667941163
transform 1 0 22724 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_241
timestamp 1667941163
transform 1 0 23276 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_247
timestamp 1667941163
transform 1 0 23828 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_253
timestamp 1667941163
transform 1 0 24380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_265
timestamp 1667941163
transform 1 0 25484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_277
timestamp 1667941163
transform 1 0 26588 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1667941163
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1667941163
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1667941163
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1667941163
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1667941163
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1667941163
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1667941163
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1667941163
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1667941163
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1667941163
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_26
timestamp 1667941163
transform 1 0 3496 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_51
timestamp 1667941163
transform 1 0 5796 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_55
timestamp 1667941163
transform 1 0 6164 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_79
timestamp 1667941163
transform 1 0 8372 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1667941163
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_105
timestamp 1667941163
transform 1 0 10764 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_129
timestamp 1667941163
transform 1 0 12972 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_60_138
timestamp 1667941163
transform 1 0 13800 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_146
timestamp 1667941163
transform 1 0 14536 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_154
timestamp 1667941163
transform 1 0 15272 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_158
timestamp 1667941163
transform 1 0 15640 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_165
timestamp 1667941163
transform 1 0 16284 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_60_174
timestamp 1667941163
transform 1 0 17112 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_186
timestamp 1667941163
transform 1 0 18216 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_193
timestamp 1667941163
transform 1 0 18860 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_201
timestamp 1667941163
transform 1 0 19596 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_207
timestamp 1667941163
transform 1 0 20148 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_213
timestamp 1667941163
transform 1 0 20700 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_219
timestamp 1667941163
transform 1 0 21252 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_225
timestamp 1667941163
transform 1 0 21804 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_231
timestamp 1667941163
transform 1 0 22356 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_237
timestamp 1667941163
transform 1 0 22908 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_243
timestamp 1667941163
transform 1 0 23460 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_249
timestamp 1667941163
transform 1 0 24012 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_257
timestamp 1667941163
transform 1 0 24748 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_269
timestamp 1667941163
transform 1 0 25852 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_281
timestamp 1667941163
transform 1 0 26956 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_293
timestamp 1667941163
transform 1 0 28060 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_305
timestamp 1667941163
transform 1 0 29164 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1667941163
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1667941163
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1667941163
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1667941163
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1667941163
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1667941163
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1667941163
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_401
timestamp 1667941163
transform 1 0 37996 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_9
timestamp 1667941163
transform 1 0 1932 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_23
timestamp 1667941163
transform 1 0 3220 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_47
timestamp 1667941163
transform 1 0 5428 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1667941163
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_61
timestamp 1667941163
transform 1 0 6716 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_86
timestamp 1667941163
transform 1 0 9016 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_110
timestamp 1667941163
transform 1 0 11224 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_135
timestamp 1667941163
transform 1 0 13524 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_141
timestamp 1667941163
transform 1 0 14076 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_148
timestamp 1667941163
transform 1 0 14720 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_159
timestamp 1667941163
transform 1 0 15732 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_166
timestamp 1667941163
transform 1 0 16376 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_174
timestamp 1667941163
transform 1 0 17112 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_178
timestamp 1667941163
transform 1 0 17480 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_182
timestamp 1667941163
transform 1 0 17848 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_190
timestamp 1667941163
transform 1 0 18584 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_196
timestamp 1667941163
transform 1 0 19136 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_202
timestamp 1667941163
transform 1 0 19688 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_208
timestamp 1667941163
transform 1 0 20240 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_214
timestamp 1667941163
transform 1 0 20792 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_220
timestamp 1667941163
transform 1 0 21344 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_229
timestamp 1667941163
transform 1 0 22172 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_235
timestamp 1667941163
transform 1 0 22724 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_241
timestamp 1667941163
transform 1 0 23276 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_247
timestamp 1667941163
transform 1 0 23828 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_253
timestamp 1667941163
transform 1 0 24380 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_259
timestamp 1667941163
transform 1 0 24932 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_265
timestamp 1667941163
transform 1 0 25484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_277
timestamp 1667941163
transform 1 0 26588 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_285
timestamp 1667941163
transform 1 0 27324 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_289
timestamp 1667941163
transform 1 0 27692 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_301
timestamp 1667941163
transform 1 0 28796 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_313
timestamp 1667941163
transform 1 0 29900 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_325
timestamp 1667941163
transform 1 0 31004 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_333
timestamp 1667941163
transform 1 0 31740 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1667941163
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1667941163
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1667941163
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1667941163
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1667941163
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_397
timestamp 1667941163
transform 1 0 37628 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_26
timestamp 1667941163
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_53
timestamp 1667941163
transform 1 0 5980 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_80
timestamp 1667941163
transform 1 0 8464 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_99
timestamp 1667941163
transform 1 0 10212 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_126
timestamp 1667941163
transform 1 0 12696 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_134
timestamp 1667941163
transform 1 0 13432 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_148
timestamp 1667941163
transform 1 0 14720 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_155
timestamp 1667941163
transform 1 0 15364 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_162
timestamp 1667941163
transform 1 0 16008 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_168
timestamp 1667941163
transform 1 0 16560 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_176
timestamp 1667941163
transform 1 0 17296 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_179
timestamp 1667941163
transform 1 0 17572 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_185
timestamp 1667941163
transform 1 0 18124 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_191
timestamp 1667941163
transform 1 0 18676 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1667941163
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_201
timestamp 1667941163
transform 1 0 19596 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_207
timestamp 1667941163
transform 1 0 20148 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_213
timestamp 1667941163
transform 1 0 20700 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_219
timestamp 1667941163
transform 1 0 21252 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_225
timestamp 1667941163
transform 1 0 21804 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_231
timestamp 1667941163
transform 1 0 22356 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_237
timestamp 1667941163
transform 1 0 22908 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_243
timestamp 1667941163
transform 1 0 23460 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_249
timestamp 1667941163
transform 1 0 24012 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_257
timestamp 1667941163
transform 1 0 24748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_263
timestamp 1667941163
transform 1 0 25300 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_269
timestamp 1667941163
transform 1 0 25852 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_281
timestamp 1667941163
transform 1 0 26956 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_293
timestamp 1667941163
transform 1 0 28060 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_305
timestamp 1667941163
transform 1 0 29164 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1667941163
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1667941163
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1667941163
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1667941163
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1667941163
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1667941163
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_405
timestamp 1667941163
transform 1 0 38364 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_9
timestamp 1667941163
transform 1 0 1932 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_30
timestamp 1667941163
transform 1 0 3864 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_54
timestamp 1667941163
transform 1 0 6072 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_83
timestamp 1667941163
transform 1 0 8740 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_110
timestamp 1667941163
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_138
timestamp 1667941163
transform 1 0 13800 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_146
timestamp 1667941163
transform 1 0 14536 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_153
timestamp 1667941163
transform 1 0 15180 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_159
timestamp 1667941163
transform 1 0 15732 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_163
timestamp 1667941163
transform 1 0 16100 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1667941163
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_174
timestamp 1667941163
transform 1 0 17112 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_178
timestamp 1667941163
transform 1 0 17480 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_182
timestamp 1667941163
transform 1 0 17848 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_190
timestamp 1667941163
transform 1 0 18584 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_194
timestamp 1667941163
transform 1 0 18952 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_201
timestamp 1667941163
transform 1 0 19596 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_207
timestamp 1667941163
transform 1 0 20148 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_213
timestamp 1667941163
transform 1 0 20700 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_219
timestamp 1667941163
transform 1 0 21252 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1667941163
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_229
timestamp 1667941163
transform 1 0 22172 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_235
timestamp 1667941163
transform 1 0 22724 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_241
timestamp 1667941163
transform 1 0 23276 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_245
timestamp 1667941163
transform 1 0 23644 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_251
timestamp 1667941163
transform 1 0 24196 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_257
timestamp 1667941163
transform 1 0 24748 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_263
timestamp 1667941163
transform 1 0 25300 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_267
timestamp 1667941163
transform 1 0 25668 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1667941163
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1667941163
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1667941163
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1667941163
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1667941163
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1667941163
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1667941163
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_344
timestamp 1667941163
transform 1 0 32752 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_350
timestamp 1667941163
transform 1 0 33304 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_358
timestamp 1667941163
transform 1 0 34040 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_364
timestamp 1667941163
transform 1 0 34592 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_370
timestamp 1667941163
transform 1 0 35144 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_382
timestamp 1667941163
transform 1 0 36248 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_390
timestamp 1667941163
transform 1 0 36984 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1667941163
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_26
timestamp 1667941163
transform 1 0 3496 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_53
timestamp 1667941163
transform 1 0 5980 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_61
timestamp 1667941163
transform 1 0 6716 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_82
timestamp 1667941163
transform 1 0 8648 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_107
timestamp 1667941163
transform 1 0 10948 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_111
timestamp 1667941163
transform 1 0 11316 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_135
timestamp 1667941163
transform 1 0 13524 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1667941163
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_153
timestamp 1667941163
transform 1 0 15180 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_161
timestamp 1667941163
transform 1 0 15916 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_167
timestamp 1667941163
transform 1 0 16468 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_175
timestamp 1667941163
transform 1 0 17204 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_181
timestamp 1667941163
transform 1 0 17756 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_187
timestamp 1667941163
transform 1 0 18308 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_193
timestamp 1667941163
transform 1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_203
timestamp 1667941163
transform 1 0 19780 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_209
timestamp 1667941163
transform 1 0 20332 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_216
timestamp 1667941163
transform 1 0 20976 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_222
timestamp 1667941163
transform 1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_231
timestamp 1667941163
transform 1 0 22356 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_237
timestamp 1667941163
transform 1 0 22908 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_243
timestamp 1667941163
transform 1 0 23460 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_247
timestamp 1667941163
transform 1 0 23828 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_250
timestamp 1667941163
transform 1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_259
timestamp 1667941163
transform 1 0 24932 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_267
timestamp 1667941163
transform 1 0 25668 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_275
timestamp 1667941163
transform 1 0 26404 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_278
timestamp 1667941163
transform 1 0 26680 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_287
timestamp 1667941163
transform 1 0 27508 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_299
timestamp 1667941163
transform 1 0 28612 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_306
timestamp 1667941163
transform 1 0 29256 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_314
timestamp 1667941163
transform 1 0 29992 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_328
timestamp 1667941163
transform 1 0 31280 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_334
timestamp 1667941163
transform 1 0 31832 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_343
timestamp 1667941163
transform 1 0 32660 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_351
timestamp 1667941163
transform 1 0 33396 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1667941163
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1667941163
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_373
timestamp 1667941163
transform 1 0 35420 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_378
timestamp 1667941163
transform 1 0 35880 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_390
timestamp 1667941163
transform 1 0 36984 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_393
timestamp 1667941163
transform 1 0 37260 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_399
timestamp 1667941163
transform 1 0 37812 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _213_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14444 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _214_
timestamp 1667941163
transform 1 0 9200 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _215_
timestamp 1667941163
transform 1 0 15732 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _216_
timestamp 1667941163
transform -1 0 18492 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _217_
timestamp 1667941163
transform 1 0 18400 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _218_
timestamp 1667941163
transform 1 0 14260 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _219_
timestamp 1667941163
transform -1 0 8004 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 1667941163
transform -1 0 14536 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _221_
timestamp 1667941163
transform 1 0 18400 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1667941163
transform 1 0 8372 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _223_
timestamp 1667941163
transform 1 0 16284 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _224_
timestamp 1667941163
transform 1 0 11040 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _225_
timestamp 1667941163
transform 1 0 11040 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _226_
timestamp 1667941163
transform 1 0 9660 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _227_
timestamp 1667941163
transform -1 0 15364 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1667941163
transform 1 0 9844 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _229_
timestamp 1667941163
transform 1 0 10948 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _230_
timestamp 1667941163
transform 1 0 7912 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _231_
timestamp 1667941163
transform 1 0 9016 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _232_
timestamp 1667941163
transform 1 0 9752 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _233_
timestamp 1667941163
transform -1 0 9936 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _234_
timestamp 1667941163
transform 1 0 5704 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1667941163
transform 1 0 8372 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _236_
timestamp 1667941163
transform 1 0 7728 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _237_
timestamp 1667941163
transform 1 0 7820 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _238_
timestamp 1667941163
transform 1 0 6532 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 1667941163
transform 1 0 9568 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 1667941163
transform 1 0 8556 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _241_
timestamp 1667941163
transform 1 0 9752 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _242_
timestamp 1667941163
transform 1 0 5796 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1667941163
transform -1 0 13616 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _244_
timestamp 1667941163
transform 1 0 8740 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _245_
timestamp 1667941163
transform 1 0 10396 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _246_
timestamp 1667941163
transform 1 0 13524 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _247_
timestamp 1667941163
transform -1 0 16284 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1667941163
transform -1 0 23460 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 1667941163
transform 1 0 23184 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _250_
timestamp 1667941163
transform 1 0 10212 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1667941163
transform 1 0 19412 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1667941163
transform -1 0 22816 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1667941163
transform -1 0 21528 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1667941163
transform 1 0 16836 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1667941163
transform -1 0 15548 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp 1667941163
transform -1 0 13708 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 1667941163
transform 1 0 9200 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 1667941163
transform -1 0 18584 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1667941163
transform 1 0 11868 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp 1667941163
transform 1 0 17112 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _261_
timestamp 1667941163
transform 1 0 11684 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp 1667941163
transform 1 0 14444 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _263_
timestamp 1667941163
transform -1 0 9936 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1667941163
transform -1 0 18216 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1667941163
transform -1 0 19872 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 1667941163
transform 1 0 14628 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _267_
timestamp 1667941163
transform 1 0 12972 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _268_
timestamp 1667941163
transform -1 0 16376 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _269_
timestamp 1667941163
transform 1 0 20608 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1667941163
transform 1 0 12512 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1667941163
transform -1 0 19688 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _272_
timestamp 1667941163
transform -1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1667941163
transform 1 0 10948 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _274_
timestamp 1667941163
transform 1 0 9568 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _275_
timestamp 1667941163
transform 1 0 19412 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _276_
timestamp 1667941163
transform 1 0 21068 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _277_
timestamp 1667941163
transform 1 0 16008 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _278_
timestamp 1667941163
transform 1 0 9292 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _279_
timestamp 1667941163
transform 1 0 12236 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1667941163
transform -1 0 17296 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _281_
timestamp 1667941163
transform -1 0 16376 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _282_
timestamp 1667941163
transform 1 0 15364 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _283_
timestamp 1667941163
transform 1 0 18400 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _284_
timestamp 1667941163
transform -1 0 15732 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _285_
timestamp 1667941163
transform -1 0 21436 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _286_
timestamp 1667941163
transform 1 0 15456 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _287_
timestamp 1667941163
transform 1 0 10304 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _288_
timestamp 1667941163
transform -1 0 20884 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _289_
timestamp 1667941163
transform -1 0 17204 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _290_
timestamp 1667941163
transform 1 0 16100 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _291_
timestamp 1667941163
transform -1 0 16376 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _292_
timestamp 1667941163
transform 1 0 13524 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _293_
timestamp 1667941163
transform 1 0 21252 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _294_
timestamp 1667941163
transform 1 0 16836 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1667941163
transform -1 0 20608 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1667941163
transform 1 0 19412 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1667941163
transform 1 0 16100 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1667941163
transform 1 0 15732 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1667941163
transform -1 0 18032 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _300_
timestamp 1667941163
transform -1 0 20516 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _301_
timestamp 1667941163
transform -1 0 21252 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _302_
timestamp 1667941163
transform 1 0 14904 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _303_
timestamp 1667941163
transform 1 0 21068 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _304_
timestamp 1667941163
transform 1 0 8372 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _305_
timestamp 1667941163
transform 1 0 13524 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _306_
timestamp 1667941163
transform 1 0 13524 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _307_
timestamp 1667941163
transform -1 0 21252 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _308_
timestamp 1667941163
transform -1 0 22264 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _309_
timestamp 1667941163
transform 1 0 9292 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1667941163
transform 1 0 12236 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _311_
timestamp 1667941163
transform -1 0 16744 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _312_
timestamp 1667941163
transform 1 0 16100 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _313_
timestamp 1667941163
transform 1 0 9476 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _314_
timestamp 1667941163
transform 1 0 17020 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _315_
timestamp 1667941163
transform -1 0 21620 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _316_
timestamp 1667941163
transform 1 0 11868 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _317_
timestamp 1667941163
transform -1 0 13800 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _318_
timestamp 1667941163
transform 1 0 8372 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _319_
timestamp 1667941163
transform 1 0 13524 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _320_
timestamp 1667941163
transform 1 0 8464 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _321_
timestamp 1667941163
transform -1 0 13156 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _322_
timestamp 1667941163
transform 1 0 7728 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _323_
timestamp 1667941163
transform -1 0 11224 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _324_
timestamp 1667941163
transform -1 0 17664 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _325_
timestamp 1667941163
transform -1 0 14720 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _326_
timestamp 1667941163
transform 1 0 7728 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _327_
timestamp 1667941163
transform 1 0 15916 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _328_
timestamp 1667941163
transform 1 0 17572 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _329_
timestamp 1667941163
transform -1 0 15364 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _330_
timestamp 1667941163
transform 1 0 12880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _331_
timestamp 1667941163
transform -1 0 17112 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _332_
timestamp 1667941163
transform 1 0 10948 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _333_
timestamp 1667941163
transform 1 0 13432 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _334_
timestamp 1667941163
transform 1 0 10304 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _335_
timestamp 1667941163
transform 1 0 19964 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _336_
timestamp 1667941163
transform 1 0 15456 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _337_
timestamp 1667941163
transform 1 0 19780 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _338_
timestamp 1667941163
transform -1 0 14720 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp 1667941163
transform -1 0 16284 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _340_
timestamp 1667941163
transform 1 0 12880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _341_
timestamp 1667941163
transform -1 0 18032 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _342_
timestamp 1667941163
transform -1 0 16928 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _343_
timestamp 1667941163
transform -1 0 30176 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _344_
timestamp 1667941163
transform 1 0 21252 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1667941163
transform -1 0 18492 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp 1667941163
transform -1 0 15364 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1667941163
transform 1 0 7084 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _348_
timestamp 1667941163
transform -1 0 20332 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _349_
timestamp 1667941163
transform 1 0 8372 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _350_
timestamp 1667941163
transform -1 0 14720 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _351_
timestamp 1667941163
transform -1 0 4784 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _352_
timestamp 1667941163
transform 1 0 8096 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _353_
timestamp 1667941163
transform -1 0 16376 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _354_
timestamp 1667941163
transform -1 0 29992 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _355_
timestamp 1667941163
transform -1 0 21344 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _356_
timestamp 1667941163
transform -1 0 13432 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _357_
timestamp 1667941163
transform -1 0 30360 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _358_
timestamp 1667941163
transform 1 0 30084 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _359_
timestamp 1667941163
transform -1 0 14720 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _360_
timestamp 1667941163
transform 1 0 9384 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _361_
timestamp 1667941163
transform -1 0 12880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _362_
timestamp 1667941163
transform -1 0 24564 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _363_
timestamp 1667941163
transform -1 0 16376 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _364_
timestamp 1667941163
transform 1 0 10304 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp 1667941163
transform 1 0 32476 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _366_
timestamp 1667941163
transform -1 0 16376 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _367_
timestamp 1667941163
transform 1 0 9752 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _368_
timestamp 1667941163
transform 1 0 9568 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _369_
timestamp 1667941163
transform -1 0 29992 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _370_
timestamp 1667941163
transform -1 0 21896 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _371_
timestamp 1667941163
transform 1 0 14628 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _372_
timestamp 1667941163
transform 1 0 34316 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _373_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 13432 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _374_
timestamp 1667941163
transform 1 0 9108 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _375_
timestamp 1667941163
transform 1 0 10304 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _376_
timestamp 1667941163
transform -1 0 17112 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _377_
timestamp 1667941163
transform 1 0 32292 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _378_
timestamp 1667941163
transform 1 0 29532 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _379_
timestamp 1667941163
transform 1 0 27416 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _380_
timestamp 1667941163
transform -1 0 18860 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _381_
timestamp 1667941163
transform -1 0 13340 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _382_
timestamp 1667941163
transform 1 0 9752 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _383_
timestamp 1667941163
transform -1 0 19688 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _384_
timestamp 1667941163
transform -1 0 6808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _385_
timestamp 1667941163
transform -1 0 7360 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _386_
timestamp 1667941163
transform -1 0 17848 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _387_
timestamp 1667941163
transform -1 0 26404 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _388_
timestamp 1667941163
transform 1 0 7176 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _389_
timestamp 1667941163
transform -1 0 20976 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _390_
timestamp 1667941163
transform 1 0 10948 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _391_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17664 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _392_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17020 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _393_
timestamp 1667941163
transform 1 0 2760 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _394_
timestamp 1667941163
transform 1 0 2300 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _395_
timestamp 1667941163
transform 1 0 2300 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _396_
timestamp 1667941163
transform 1 0 5888 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _397_
timestamp 1667941163
transform 1 0 6900 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _398_
timestamp 1667941163
transform 1 0 8280 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _399_
timestamp 1667941163
transform 1 0 2116 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _400_
timestamp 1667941163
transform 1 0 3956 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _401_
timestamp 1667941163
transform 1 0 2116 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _402_
timestamp 1667941163
transform 1 0 5796 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _403_
timestamp 1667941163
transform 1 0 18124 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _404_
timestamp 1667941163
transform 1 0 3220 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _405_
timestamp 1667941163
transform 1 0 3588 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _406_
timestamp 1667941163
transform 1 0 4600 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _407_
timestamp 1667941163
transform 1 0 2484 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _408_
timestamp 1667941163
transform -1 0 5152 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _409_
timestamp 1667941163
transform 1 0 2300 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _410_
timestamp 1667941163
transform -1 0 6072 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _411_
timestamp 1667941163
transform 1 0 2944 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _412_
timestamp 1667941163
transform 1 0 3128 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _413_
timestamp 1667941163
transform 1 0 1840 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _414_
timestamp 1667941163
transform -1 0 17388 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _415_
timestamp 1667941163
transform 1 0 5796 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _416_
timestamp 1667941163
transform 1 0 7176 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _417_
timestamp 1667941163
transform 1 0 7912 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _418_
timestamp 1667941163
transform 1 0 7452 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _419_
timestamp 1667941163
transform 1 0 3956 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _420_
timestamp 1667941163
transform 1 0 4232 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _421_
timestamp 1667941163
transform 1 0 4600 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _422_
timestamp 1667941163
transform 1 0 6624 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _423_
timestamp 1667941163
transform 1 0 3312 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _424_
timestamp 1667941163
transform 1 0 5244 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _425_
timestamp 1667941163
transform -1 0 16836 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _426_
timestamp 1667941163
transform 1 0 2944 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _427_
timestamp 1667941163
transform 1 0 2024 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _428_
timestamp 1667941163
transform -1 0 2944 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _429_
timestamp 1667941163
transform 1 0 7268 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _430_
timestamp 1667941163
transform 1 0 6532 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _431_
timestamp 1667941163
transform 1 0 6808 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _432_
timestamp 1667941163
transform 1 0 1840 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _433_
timestamp 1667941163
transform -1 0 3864 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _434_
timestamp 1667941163
transform -1 0 2760 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _435_
timestamp 1667941163
transform 1 0 7728 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _436_
timestamp 1667941163
transform 1 0 17204 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _437_
timestamp 1667941163
transform -1 0 18676 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _438_
timestamp 1667941163
transform -1 0 14812 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _439_
timestamp 1667941163
transform -1 0 18860 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _440_
timestamp 1667941163
transform -1 0 17848 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _441_
timestamp 1667941163
transform -1 0 19320 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _442_
timestamp 1667941163
transform -1 0 20884 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _443_
timestamp 1667941163
transform -1 0 18860 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _444_
timestamp 1667941163
transform -1 0 20976 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _445_
timestamp 1667941163
transform -1 0 8096 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _446_
timestamp 1667941163
transform -1 0 8648 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _447_
timestamp 1667941163
transform -1 0 17388 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _448_
timestamp 1667941163
transform -1 0 13156 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _449_
timestamp 1667941163
transform -1 0 13800 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _450_
timestamp 1667941163
transform 1 0 20884 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _451_
timestamp 1667941163
transform -1 0 20332 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _452_
timestamp 1667941163
transform -1 0 18216 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _453_
timestamp 1667941163
transform -1 0 16284 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _454_
timestamp 1667941163
transform 1 0 20976 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _455_
timestamp 1667941163
transform -1 0 20884 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _456_
timestamp 1667941163
transform -1 0 17020 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _457_
timestamp 1667941163
transform -1 0 13156 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _458_
timestamp 1667941163
transform -1 0 18952 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _459_
timestamp 1667941163
transform -1 0 19596 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _460_
timestamp 1667941163
transform 1 0 20332 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _461_
timestamp 1667941163
transform -1 0 19964 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _462_
timestamp 1667941163
transform -1 0 19688 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _463_
timestamp 1667941163
transform -1 0 20332 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _464_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3956 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _465_
timestamp 1667941163
transform -1 0 3864 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _466_
timestamp 1667941163
transform -1 0 5796 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _467_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 8740 0 -1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _468_
timestamp 1667941163
transform -1 0 12052 0 1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _469_
timestamp 1667941163
transform -1 0 13800 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _470_
timestamp 1667941163
transform 1 0 3220 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _471_
timestamp 1667941163
transform -1 0 5428 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _472_
timestamp 1667941163
transform -1 0 5796 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _473_
timestamp 1667941163
transform -1 0 8648 0 1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _474_
timestamp 1667941163
transform -1 0 8556 0 1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _475_
timestamp 1667941163
transform 1 0 5796 0 1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _476_
timestamp 1667941163
transform 1 0 4140 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _477_
timestamp 1667941163
transform 1 0 1656 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _478_
timestamp 1667941163
transform -1 0 3496 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _479_
timestamp 1667941163
transform -1 0 6072 0 -1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _480_
timestamp 1667941163
transform 1 0 3956 0 -1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _481_
timestamp 1667941163
transform -1 0 8464 0 1 35904
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _482_
timestamp 1667941163
transform 1 0 4140 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _483_
timestamp 1667941163
transform -1 0 6072 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _484_
timestamp 1667941163
transform -1 0 13524 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _485_
timestamp 1667941163
transform -1 0 12328 0 1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _486_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 11316 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _487_
timestamp 1667941163
transform 1 0 10856 0 1 34816
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _488_
timestamp 1667941163
transform -1 0 11224 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _489_
timestamp 1667941163
transform -1 0 13524 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _490_
timestamp 1667941163
transform 1 0 11684 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _491_
timestamp 1667941163
transform -1 0 10396 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _492_
timestamp 1667941163
transform -1 0 8648 0 -1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _493_
timestamp 1667941163
transform -1 0 12696 0 1 35904
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _494_
timestamp 1667941163
transform 1 0 3956 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _495_
timestamp 1667941163
transform 1 0 1656 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _496_
timestamp 1667941163
transform -1 0 3588 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _497_
timestamp 1667941163
transform -1 0 9108 0 -1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _498_
timestamp 1667941163
transform -1 0 13800 0 -1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _499_
timestamp 1667941163
transform -1 0 11224 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _500_
timestamp 1667941163
transform -1 0 3496 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _501_
timestamp 1667941163
transform 1 0 2024 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _502_
timestamp 1667941163
transform -1 0 3496 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _503_
timestamp 1667941163
transform -1 0 11224 0 -1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _504_
timestamp 1667941163
transform 1 0 11684 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _505_
timestamp 1667941163
transform 1 0 9292 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _506_
timestamp 1667941163
transform -1 0 10948 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _507_
timestamp 1667941163
transform 1 0 6900 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _508_
timestamp 1667941163
transform -1 0 8648 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _509_
timestamp 1667941163
transform 1 0 8924 0 -1 34816
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _510_
timestamp 1667941163
transform 1 0 9108 0 1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _511_
timestamp 1667941163
transform 1 0 6256 0 1 34816
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _512_
timestamp 1667941163
transform 1 0 3956 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _513_
timestamp 1667941163
transform 1 0 3956 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _514_
timestamp 1667941163
transform -1 0 6072 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _515_
timestamp 1667941163
transform 1 0 6808 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _516_
timestamp 1667941163
transform 1 0 11684 0 -1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _517_
timestamp 1667941163
transform -1 0 9016 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _518_
timestamp 1667941163
transform 1 0 9108 0 -1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _519_
timestamp 1667941163
transform 1 0 1748 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _520_
timestamp 1667941163
transform -1 0 5796 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _521_
timestamp 1667941163
transform 1 0 10856 0 1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _522_
timestamp 1667941163
transform -1 0 12144 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _523_
timestamp 1667941163
transform 1 0 6256 0 1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _524_
timestamp 1667941163
transform 1 0 1656 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _525_
timestamp 1667941163
transform -1 0 3588 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _526_
timestamp 1667941163
transform -1 0 10856 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _527_
timestamp 1667941163
transform -1 0 13524 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _528_
timestamp 1667941163
transform 1 0 11592 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _529_
timestamp 1667941163
transform 1 0 6716 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _541_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 33580 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _542_
timestamp 1667941163
transform -1 0 16100 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _543_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 20792 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _544_
timestamp 1667941163
transform 1 0 14260 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _545_
timestamp 1667941163
transform -1 0 38088 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _546_
timestamp 1667941163
transform -1 0 19964 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _547_
timestamp 1667941163
transform 1 0 13248 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _548_
timestamp 1667941163
transform 1 0 16100 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _549_
timestamp 1667941163
transform -1 0 30176 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _550_
timestamp 1667941163
transform -1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _551_
timestamp 1667941163
transform 1 0 13340 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _552_
timestamp 1667941163
transform 1 0 16836 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _553_
timestamp 1667941163
transform 1 0 21988 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _554_
timestamp 1667941163
transform 1 0 17296 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _555_
timestamp 1667941163
transform 1 0 25576 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _556_
timestamp 1667941163
transform 1 0 15824 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _557_
timestamp 1667941163
transform -1 0 23460 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _558_
timestamp 1667941163
transform -1 0 38088 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _559_
timestamp 1667941163
transform 1 0 18032 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _560_
timestamp 1667941163
transform -1 0 15732 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _561_
timestamp 1667941163
transform 1 0 8372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _562_
timestamp 1667941163
transform 1 0 9200 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _563_
timestamp 1667941163
transform -1 0 20240 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _564_
timestamp 1667941163
transform 1 0 7084 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _565_
timestamp 1667941163
transform 1 0 5244 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _566_
timestamp 1667941163
transform -1 0 7820 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _567_
timestamp 1667941163
transform -1 0 38088 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _568_
timestamp 1667941163
transform -1 0 34132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _569_
timestamp 1667941163
transform 1 0 1748 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _570_
timestamp 1667941163
transform -1 0 23920 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _571_
timestamp 1667941163
transform 1 0 3956 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _572_
timestamp 1667941163
transform 1 0 37812 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _573_
timestamp 1667941163
transform -1 0 15732 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _574_
timestamp 1667941163
transform -1 0 25668 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _575_
timestamp 1667941163
transform -1 0 23644 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _576_
timestamp 1667941163
transform -1 0 18952 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _577_
timestamp 1667941163
transform 1 0 2300 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _578_
timestamp 1667941163
transform 1 0 7084 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _579_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 17756 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _580_
timestamp 1667941163
transform 1 0 13524 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _581_
timestamp 1667941163
transform -1 0 15548 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _582_
timestamp 1667941163
transform 1 0 14076 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _583__91 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 20056 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _583_
timestamp 1667941163
transform 1 0 19964 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _584_
timestamp 1667941163
transform 1 0 17756 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _585_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19044 0 -1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _586_
timestamp 1667941163
transform 1 0 14260 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _587_
timestamp 1667941163
transform 1 0 15548 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _588_
timestamp 1667941163
transform 1 0 13708 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _589_
timestamp 1667941163
transform 1 0 20056 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _590_
timestamp 1667941163
transform 1 0 14260 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _591_
timestamp 1667941163
transform -1 0 10672 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _592__92
timestamp 1667941163
transform -1 0 13800 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _592_
timestamp 1667941163
transform 1 0 14260 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _593_
timestamp 1667941163
transform -1 0 15640 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _594_
timestamp 1667941163
transform -1 0 10948 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _595_
timestamp 1667941163
transform -1 0 13064 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _596_
timestamp 1667941163
transform 1 0 11408 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _597_
timestamp 1667941163
transform -1 0 14444 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _598_
timestamp 1667941163
transform -1 0 19688 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _599_
timestamp 1667941163
transform -1 0 10672 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _600_
timestamp 1667941163
transform -1 0 11224 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _601_
timestamp 1667941163
transform -1 0 17572 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _602_
timestamp 1667941163
transform -1 0 13984 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _603_
timestamp 1667941163
transform 1 0 17112 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _604_
timestamp 1667941163
transform 1 0 14352 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _605_
timestamp 1667941163
transform 1 0 11684 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _606__93
timestamp 1667941163
transform 1 0 21988 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _606_
timestamp 1667941163
transform -1 0 17664 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _607_
timestamp 1667941163
transform 1 0 12972 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _608_
timestamp 1667941163
transform 1 0 12880 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _609_
timestamp 1667941163
transform 1 0 11684 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _610_
timestamp 1667941163
transform -1 0 18952 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _611_
timestamp 1667941163
transform 1 0 15272 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _612_
timestamp 1667941163
transform 1 0 15548 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _613_
timestamp 1667941163
transform -1 0 15272 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _614_
timestamp 1667941163
transform -1 0 19780 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _615_
timestamp 1667941163
transform 1 0 13892 0 -1 34816
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _616_
timestamp 1667941163
transform -1 0 15640 0 1 33728
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _617_
timestamp 1667941163
transform 1 0 17204 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _618__94
timestamp 1667941163
transform -1 0 19320 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _618_
timestamp 1667941163
transform -1 0 20240 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _619_
timestamp 1667941163
transform 1 0 13892 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _620_
timestamp 1667941163
transform 1 0 10396 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _621_
timestamp 1667941163
transform 1 0 18216 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _622_
timestamp 1667941163
transform -1 0 20700 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _623_
timestamp 1667941163
transform -1 0 19044 0 -1 33728
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _624_
timestamp 1667941163
transform -1 0 16652 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _625_
timestamp 1667941163
transform -1 0 20608 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _626_
timestamp 1667941163
transform 1 0 19412 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _627_
timestamp 1667941163
transform 1 0 17388 0 1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _628_
timestamp 1667941163
transform 1 0 16836 0 -1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _629_
timestamp 1667941163
transform -1 0 14536 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _630__95
timestamp 1667941163
transform -1 0 14536 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _630_
timestamp 1667941163
transform 1 0 16376 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _631_
timestamp 1667941163
transform -1 0 21712 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _632_
timestamp 1667941163
transform 1 0 14352 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _633_
timestamp 1667941163
transform -1 0 20424 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _634_
timestamp 1667941163
transform 1 0 14352 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _635_
timestamp 1667941163
transform 1 0 16836 0 -1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _636_
timestamp 1667941163
transform 1 0 14628 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _637_
timestamp 1667941163
transform 1 0 15180 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _638_
timestamp 1667941163
transform -1 0 19504 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _639_
timestamp 1667941163
transform 1 0 15180 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _640_
timestamp 1667941163
transform 1 0 22908 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _641_
timestamp 1667941163
transform 1 0 18768 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _642__96
timestamp 1667941163
transform 1 0 21988 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _642_
timestamp 1667941163
transform 1 0 21804 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _643_
timestamp 1667941163
transform 1 0 14076 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _644_
timestamp 1667941163
transform -1 0 15824 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _645_
timestamp 1667941163
transform 1 0 12972 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _646_
timestamp 1667941163
transform -1 0 17848 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _647_
timestamp 1667941163
transform 1 0 16284 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _648_
timestamp 1667941163
transform 1 0 20148 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _649_
timestamp 1667941163
transform 1 0 14260 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _650_
timestamp 1667941163
transform 1 0 12972 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _651_
timestamp 1667941163
transform 1 0 20148 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _652_
timestamp 1667941163
transform 1 0 16928 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _653_
timestamp 1667941163
transform -1 0 19228 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _654__97
timestamp 1667941163
transform -1 0 17204 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _654_
timestamp 1667941163
transform 1 0 17204 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _655_
timestamp 1667941163
transform -1 0 19228 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _656_
timestamp 1667941163
transform -1 0 15548 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _657_
timestamp 1667941163
transform 1 0 14904 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _658_
timestamp 1667941163
transform -1 0 17572 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _659_
timestamp 1667941163
transform 1 0 17480 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _660_
timestamp 1667941163
transform 1 0 12144 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _661_
timestamp 1667941163
transform 1 0 12512 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _662_
timestamp 1667941163
transform 1 0 14812 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _663_
timestamp 1667941163
transform 1 0 15548 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _664_
timestamp 1667941163
transform -1 0 19872 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _665_
timestamp 1667941163
transform 1 0 20424 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _666__98
timestamp 1667941163
transform -1 0 21896 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _666_
timestamp 1667941163
transform -1 0 22816 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _667_
timestamp 1667941163
transform 1 0 12328 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _668_
timestamp 1667941163
transform 1 0 12972 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _669_
timestamp 1667941163
transform 1 0 23184 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _670_
timestamp 1667941163
transform -1 0 22816 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _671_
timestamp 1667941163
transform 1 0 17664 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _672_
timestamp 1667941163
transform 1 0 19412 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _673_
timestamp 1667941163
transform -1 0 15364 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _674_
timestamp 1667941163
transform 1 0 14812 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _675_
timestamp 1667941163
transform -1 0 11224 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _676_
timestamp 1667941163
transform -1 0 9752 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _677_
timestamp 1667941163
transform 1 0 10948 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _678__99
timestamp 1667941163
transform -1 0 8648 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _678_
timestamp 1667941163
transform 1 0 9292 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _679_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 12696 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _680_
timestamp 1667941163
transform 1 0 10488 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _681_
timestamp 1667941163
transform 1 0 9016 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _682_
timestamp 1667941163
transform 1 0 10396 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _683_
timestamp 1667941163
transform 1 0 9108 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _684_
timestamp 1667941163
transform -1 0 13708 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _685_
timestamp 1667941163
transform -1 0 12604 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _686_
timestamp 1667941163
transform -1 0 12696 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _687_
timestamp 1667941163
transform -1 0 10764 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _688_
timestamp 1667941163
transform -1 0 12512 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _689_
timestamp 1667941163
transform -1 0 15732 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _690__100
timestamp 1667941163
transform -1 0 8648 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _690_
timestamp 1667941163
transform 1 0 12880 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _691_
timestamp 1667941163
transform -1 0 13432 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _692_
timestamp 1667941163
transform 1 0 10488 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _693_
timestamp 1667941163
transform 1 0 12972 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _694_
timestamp 1667941163
transform 1 0 11684 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _695_
timestamp 1667941163
transform -1 0 11960 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _696_
timestamp 1667941163
transform -1 0 15088 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _697_
timestamp 1667941163
transform 1 0 11684 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _698_
timestamp 1667941163
transform -1 0 16836 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _699_
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _700__101
timestamp 1667941163
transform 1 0 19412 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _700_
timestamp 1667941163
transform 1 0 19412 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _701_
timestamp 1667941163
transform -1 0 18952 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _702_
timestamp 1667941163
transform -1 0 13984 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _703_
timestamp 1667941163
transform -1 0 18768 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _704_
timestamp 1667941163
transform 1 0 15548 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _705_
timestamp 1667941163
transform 1 0 15272 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _706_
timestamp 1667941163
transform 1 0 11224 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _707_
timestamp 1667941163
transform 1 0 11684 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1667941163
transform -1 0 32660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1667941163
transform 1 0 20700 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 2944 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1667941163
transform -1 0 37812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1667941163
transform 1 0 14904 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1667941163
transform 1 0 1564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1667941163
transform -1 0 38364 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1667941163
transform -1 0 15180 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1667941163
transform 1 0 2300 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1667941163
transform 1 0 3956 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1667941163
transform -1 0 38364 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1667941163
transform 1 0 9752 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp 1667941163
transform -1 0 38364 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1667941163
transform -1 0 17204 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1667941163
transform -1 0 38364 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1667941163
transform 1 0 1564 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1667941163
transform -1 0 24932 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1667941163
transform -1 0 38364 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1667941163
transform 1 0 4692 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1667941163
transform 1 0 1564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1667941163
transform 1 0 9108 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1667941163
transform 1 0 3956 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1667941163
transform 1 0 11684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1667941163
transform -1 0 33948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1667941163
transform -1 0 38364 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1667941163
transform -1 0 38364 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1667941163
transform 1 0 1564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1667941163
transform 1 0 1564 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1667941163
transform -1 0 36984 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1667941163
transform 1 0 1564 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1667941163
transform -1 0 38364 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1667941163
transform -1 0 1840 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1667941163
transform 1 0 29716 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input34
timestamp 1667941163
transform -1 0 38364 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input35
timestamp 1667941163
transform -1 0 10212 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input36
timestamp 1667941163
transform -1 0 3220 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1667941163
transform 1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1667941163
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1667941163
transform -1 0 23644 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1667941163
transform 1 0 30360 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  output41 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37996 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1667941163
transform 1 0 37996 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1667941163
transform 1 0 37996 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1667941163
transform 1 0 37996 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1667941163
transform 1 0 37996 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1667941163
transform 1 0 35512 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1667941163
transform -1 0 1932 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1667941163
transform -1 0 1932 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1667941163
transform 1 0 37996 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1667941163
transform -1 0 1932 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1667941163
transform 1 0 8280 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1667941163
transform 1 0 19412 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1667941163
transform -1 0 15916 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1667941163
transform 1 0 37996 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1667941163
transform 1 0 25300 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1667941163
transform 1 0 27140 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1667941163
transform -1 0 35236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1667941163
transform -1 0 1932 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1667941163
transform 1 0 37996 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1667941163
transform 1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1667941163
transform -1 0 1932 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1667941163
transform 1 0 35880 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1667941163
transform 1 0 37996 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1667941163
transform -1 0 5612 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1667941163
transform -1 0 1932 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1667941163
transform -1 0 1932 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1667941163
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1667941163
transform -1 0 1932 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1667941163
transform -1 0 13432 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1667941163
transform 1 0 21988 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1667941163
transform 1 0 33580 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1667941163
transform -1 0 1932 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1667941163
transform -1 0 1932 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1667941163
transform -1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1667941163
transform 1 0 37444 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1667941163
transform 1 0 28888 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1667941163
transform 1 0 16836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1667941163
transform -1 0 36984 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1667941163
transform 1 0 37996 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1667941163
transform -1 0 1932 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1667941163
transform 1 0 37996 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1667941163
transform -1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1667941163
transform -1 0 13340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1667941163
transform 1 0 20056 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1667941163
transform 1 0 37996 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1667941163
transform 1 0 21988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1667941163
transform 1 0 32292 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1667941163
transform -1 0 14536 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1667941163
transform 1 0 27140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1667941163
transform -1 0 1932 0 -1 13056
box -38 -48 406 592
<< labels >>
flabel metal3 s 39200 26528 39800 26648 0 FreeSans 480 0 0 0 bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
port 0 nsew signal tristate
flabel metal3 s 39200 37408 39800 37528 0 FreeSans 480 0 0 0 bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
port 1 nsew signal tristate
flabel metal2 s 38658 39200 38714 39800 0 FreeSans 224 90 0 0 bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_
port 2 nsew signal tristate
flabel metal2 s 38014 200 38070 800 0 FreeSans 224 90 0 0 bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
port 3 nsew signal tristate
flabel metal3 s 39200 19728 39800 19848 0 FreeSans 480 0 0 0 bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_
port 4 nsew signal tristate
flabel metal2 s 35438 39200 35494 39800 0 FreeSans 224 90 0 0 bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_
port 5 nsew signal tristate
flabel metal3 s 200 3408 800 3528 0 FreeSans 480 0 0 0 bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_
port 6 nsew signal tristate
flabel metal3 s 200 19048 800 19168 0 FreeSans 480 0 0 0 bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_
port 7 nsew signal tristate
flabel metal2 s 31574 200 31630 800 0 FreeSans 224 90 0 0 ccff_head
port 8 nsew signal input
flabel metal3 s 39200 12248 39800 12368 0 FreeSans 480 0 0 0 ccff_tail
port 9 nsew signal tristate
flabel metal2 s 20626 39200 20682 39800 0 FreeSans 224 90 0 0 chanx_left_in[0]
port 10 nsew signal input
flabel metal2 s 1950 39200 2006 39800 0 FreeSans 224 90 0 0 chanx_left_in[10]
port 11 nsew signal input
flabel metal2 s 36726 200 36782 800 0 FreeSans 224 90 0 0 chanx_left_in[11]
port 12 nsew signal input
flabel metal2 s 14830 200 14886 800 0 FreeSans 224 90 0 0 chanx_left_in[12]
port 13 nsew signal input
flabel metal3 s 200 4768 800 4888 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 14 nsew signal input
flabel metal3 s 39200 33328 39800 33448 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 15 nsew signal input
flabel metal2 s 13542 39200 13598 39800 0 FreeSans 224 90 0 0 chanx_left_in[15]
port 16 nsew signal input
flabel metal3 s 200 38768 800 38888 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 17 nsew signal input
flabel metal3 s 200 33328 800 33448 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 18 nsew signal input
flabel metal3 s 39200 5448 39800 5568 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 19 nsew signal input
flabel metal2 s 9678 200 9734 800 0 FreeSans 224 90 0 0 chanx_left_in[1]
port 20 nsew signal input
flabel metal3 s 39200 28568 39800 28688 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 21 nsew signal input
flabel metal2 s 16762 39200 16818 39800 0 FreeSans 224 90 0 0 chanx_left_in[3]
port 22 nsew signal input
flabel metal3 s 39200 31968 39800 32088 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 23 nsew signal input
flabel metal3 s 200 27888 800 28008 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 24 nsew signal input
flabel metal2 s 23846 39200 23902 39800 0 FreeSans 224 90 0 0 chanx_left_in[6]
port 25 nsew signal input
flabel metal3 s 39200 29928 39800 30048 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 26 nsew signal input
flabel metal2 s 18 39200 74 39800 0 FreeSans 224 90 0 0 chanx_left_in[8]
port 27 nsew signal input
flabel metal3 s 200 1368 800 1488 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 28 nsew signal input
flabel metal3 s 200 15648 800 15768 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 29 nsew signal tristate
flabel metal2 s 8390 200 8446 800 0 FreeSans 224 90 0 0 chanx_left_out[10]
port 30 nsew signal tristate
flabel metal2 s 18694 39200 18750 39800 0 FreeSans 224 90 0 0 chanx_left_out[11]
port 31 nsew signal tristate
flabel metal2 s 15474 39200 15530 39800 0 FreeSans 224 90 0 0 chanx_left_out[12]
port 32 nsew signal tristate
flabel metal3 s 39200 8848 39800 8968 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 33 nsew signal tristate
flabel metal2 s 25134 39200 25190 39800 0 FreeSans 224 90 0 0 chanx_left_out[14]
port 34 nsew signal tristate
flabel metal2 s 27066 39200 27122 39800 0 FreeSans 224 90 0 0 chanx_left_out[15]
port 35 nsew signal tristate
flabel metal2 s 34794 200 34850 800 0 FreeSans 224 90 0 0 chanx_left_out[16]
port 36 nsew signal tristate
flabel metal3 s 200 17688 800 17808 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 37 nsew signal tristate
flabel metal3 s 39200 35368 39800 35488 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 38 nsew signal tristate
flabel metal2 s 25134 200 25190 800 0 FreeSans 224 90 0 0 chanx_left_out[1]
port 39 nsew signal tristate
flabel metal3 s 200 21088 800 21208 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 40 nsew signal tristate
flabel metal3 s 39200 2048 39800 2168 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 41 nsew signal tristate
flabel metal3 s 39200 15648 39800 15768 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 42 nsew signal tristate
flabel metal2 s 4526 200 4582 800 0 FreeSans 224 90 0 0 chanx_left_out[5]
port 43 nsew signal tristate
flabel metal3 s 200 13608 800 13728 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 44 nsew signal tristate
flabel metal3 s 200 31288 800 31408 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 45 nsew signal tristate
flabel metal2 s 28354 200 28410 800 0 FreeSans 224 90 0 0 chanx_left_out[8]
port 46 nsew signal tristate
flabel metal3 s 200 29928 800 30048 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 47 nsew signal tristate
flabel metal2 s 7102 39200 7158 39800 0 FreeSans 224 90 0 0 chanx_right_in[0]
port 48 nsew signal input
flabel metal2 s 3238 200 3294 800 0 FreeSans 224 90 0 0 chanx_right_in[10]
port 49 nsew signal input
flabel metal2 s 11610 200 11666 800 0 FreeSans 224 90 0 0 chanx_right_in[11]
port 50 nsew signal input
flabel metal2 s 33506 200 33562 800 0 FreeSans 224 90 0 0 chanx_right_in[12]
port 51 nsew signal input
flabel metal3 s 39200 14288 39800 14408 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 52 nsew signal input
flabel metal3 s 39200 6808 39800 6928 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 53 nsew signal input
flabel metal3 s 200 6808 800 6928 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 54 nsew signal input
flabel metal3 s 200 36728 800 36848 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 55 nsew signal input
flabel metal3 s 39200 8 39800 128 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 56 nsew signal input
flabel metal3 s 200 8848 800 8968 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 57 nsew signal input
flabel metal3 s 39200 10888 39800 11008 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 58 nsew signal input
flabel metal3 s 200 24488 800 24608 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 59 nsew signal input
flabel metal2 s 29642 200 29698 800 0 FreeSans 224 90 0 0 chanx_right_in[3]
port 60 nsew signal input
flabel metal3 s 39200 24488 39800 24608 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 61 nsew signal input
flabel metal2 s 10322 39200 10378 39800 0 FreeSans 224 90 0 0 chanx_right_in[5]
port 62 nsew signal input
flabel metal2 s 5170 39200 5226 39800 0 FreeSans 224 90 0 0 chanx_right_in[6]
port 63 nsew signal input
flabel metal2 s 18050 200 18106 800 0 FreeSans 224 90 0 0 chanx_right_in[7]
port 64 nsew signal input
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 chanx_right_in[8]
port 65 nsew signal input
flabel metal2 s 23202 200 23258 800 0 FreeSans 224 90 0 0 chanx_right_in[9]
port 66 nsew signal input
flabel metal2 s 12254 39200 12310 39800 0 FreeSans 224 90 0 0 chanx_right_out[0]
port 67 nsew signal tristate
flabel metal2 s 21914 39200 21970 39800 0 FreeSans 224 90 0 0 chanx_right_out[10]
port 68 nsew signal tristate
flabel metal2 s 33506 39200 33562 39800 0 FreeSans 224 90 0 0 chanx_right_out[11]
port 69 nsew signal tristate
flabel metal3 s 200 26528 800 26648 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 70 nsew signal tristate
flabel metal3 s 200 22448 800 22568 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 71 nsew signal tristate
flabel metal2 s 1306 200 1362 800 0 FreeSans 224 90 0 0 chanx_right_out[14]
port 72 nsew signal tristate
flabel metal2 s 37370 39200 37426 39800 0 FreeSans 224 90 0 0 chanx_right_out[15]
port 73 nsew signal tristate
flabel metal2 s 28998 39200 29054 39800 0 FreeSans 224 90 0 0 chanx_right_out[16]
port 74 nsew signal tristate
flabel metal2 s 16762 200 16818 800 0 FreeSans 224 90 0 0 chanx_right_out[17]
port 75 nsew signal tristate
flabel metal3 s 39200 38768 39800 38888 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 76 nsew signal tristate
flabel metal3 s 39200 3408 39800 3528 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 77 nsew signal tristate
flabel metal3 s 200 10208 800 10328 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 78 nsew signal tristate
flabel metal3 s 39200 21088 39800 21208 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 79 nsew signal tristate
flabel metal2 s 6458 200 6514 800 0 FreeSans 224 90 0 0 chanx_right_out[4]
port 80 nsew signal tristate
flabel metal2 s 12898 200 12954 800 0 FreeSans 224 90 0 0 chanx_right_out[5]
port 81 nsew signal tristate
flabel metal2 s 19982 200 20038 800 0 FreeSans 224 90 0 0 chanx_right_out[6]
port 82 nsew signal tristate
flabel metal3 s 39200 23128 39800 23248 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 83 nsew signal tristate
flabel metal2 s 21270 200 21326 800 0 FreeSans 224 90 0 0 chanx_right_out[8]
port 84 nsew signal tristate
flabel metal2 s 32218 39200 32274 39800 0 FreeSans 224 90 0 0 chanx_right_out[9]
port 85 nsew signal tristate
flabel metal2 s 30286 39200 30342 39800 0 FreeSans 224 90 0 0 pReset
port 86 nsew signal input
flabel metal2 s 3882 39200 3938 39800 0 FreeSans 224 90 0 0 prog_clk
port 87 nsew signal input
flabel metal2 s 8390 39200 8446 39800 0 FreeSans 224 90 0 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_
port 88 nsew signal tristate
flabel metal2 s 26422 200 26478 800 0 FreeSans 224 90 0 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_
port 89 nsew signal tristate
flabel metal3 s 200 12248 800 12368 0 FreeSans 480 0 0 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_
port 90 nsew signal tristate
flabel metal3 s 200 35368 800 35488 0 FreeSans 480 0 0 0 vccd1
port 91 nsew signal bidirectional
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 91 nsew signal bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 91 nsew signal bidirectional
flabel metal3 s 39200 17688 39800 17808 0 FreeSans 480 0 0 0 vssd1
port 92 nsew signal bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 92 nsew signal bidirectional
rlabel metal1 19964 37536 19964 37536 0 vccd1
rlabel metal1 19964 36992 19964 36992 0 vssd1
rlabel metal1 3818 28594 3818 28594 0 _000_
rlabel metal2 2438 30396 2438 30396 0 _001_
rlabel via1 4094 28101 4094 28101 0 _002_
rlabel metal1 6532 28662 6532 28662 0 _003_
rlabel metal2 9246 28407 9246 28407 0 _004_
rlabel metal1 9614 33014 9614 33014 0 _005_
rlabel metal2 4646 28934 4646 28934 0 _006_
rlabel metal1 4048 28662 4048 28662 0 _007_
rlabel metal2 4830 29954 4830 29954 0 _008_
rlabel metal1 5980 29274 5980 29274 0 _009_
rlabel metal1 5152 30906 5152 30906 0 _010_
rlabel metal1 5474 27982 5474 27982 0 _011_
rlabel metal1 5244 27574 5244 27574 0 _012_
rlabel metal1 2576 26010 2576 26010 0 _013_
rlabel metal2 2622 30600 2622 30600 0 _014_
rlabel metal1 2346 27098 2346 27098 0 _015_
rlabel metal2 5934 33966 5934 33966 0 _016_
rlabel metal1 8241 36074 8241 36074 0 _017_
rlabel metal2 3404 33014 3404 33014 0 _018_
rlabel metal1 1656 26010 1656 26010 0 _019_
rlabel metal1 6624 27846 6624 27846 0 _020_
rlabel metal1 7966 29036 7966 29036 0 _021_
rlabel metal1 8970 29750 8970 29750 0 _022_
rlabel metal3 9522 34884 9522 34884 0 _023_
rlabel metal3 9729 34612 9729 34612 0 _024_
rlabel metal1 9982 35598 9982 35598 0 _025_
rlabel metal2 12512 33116 12512 33116 0 _026_
rlabel metal1 6716 29818 6716 29818 0 _027_
rlabel metal1 7077 32470 7077 32470 0 _028_
rlabel via3 11339 35972 11339 35972 0 _029_
rlabel metal1 4094 27914 4094 27914 0 _030_
rlabel metal2 3082 28594 3082 28594 0 _031_
rlabel metal2 2714 29988 2714 29988 0 _032_
rlabel metal1 7360 29750 7360 29750 0 _033_
rlabel metal2 6670 29325 6670 29325 0 _034_
rlabel metal2 8326 28713 8326 28713 0 _035_
rlabel metal1 2024 26554 2024 26554 0 _036_
rlabel metal1 3641 36822 3641 36822 0 _037_
rlabel metal1 2392 26554 2392 26554 0 _038_
rlabel metal2 10258 28900 10258 28900 0 _039_
rlabel metal2 18538 30464 18538 30464 0 _040_
rlabel metal2 14674 31875 14674 31875 0 _041_
rlabel metal2 18722 35683 18722 35683 0 _042_
rlabel metal1 16100 35802 16100 35802 0 _043_
rlabel metal2 19182 35496 19182 35496 0 _044_
rlabel metal2 20746 32198 20746 32198 0 _045_
rlabel metal1 18630 33082 18630 33082 0 _046_
rlabel via2 21114 32827 21114 32827 0 _047_
rlabel metal1 7222 29274 7222 29274 0 _048_
rlabel metal1 7728 28390 7728 28390 0 _049_
rlabel metal2 6854 30056 6854 30056 0 _050_
rlabel metal1 13202 30906 13202 30906 0 _051_
rlabel metal1 15502 33626 15502 33626 0 _052_
rlabel metal1 19642 34170 19642 34170 0 _053_
rlabel metal1 16606 33082 16606 33082 0 _054_
rlabel metal1 4646 34680 4646 34680 0 _055_
rlabel metal2 21666 35870 21666 35870 0 _056_
rlabel metal2 20746 30464 20746 30464 0 _057_
rlabel metal1 15272 31994 15272 31994 0 _058_
rlabel metal1 7682 34041 7682 34041 0 _059_
rlabel metal2 18814 35785 18814 35785 0 _060_
rlabel via2 2714 33541 2714 33541 0 _061_
rlabel metal3 20240 30532 20240 30532 0 _062_
rlabel metal2 17434 32249 17434 32249 0 _063_
rlabel metal2 19550 33184 19550 33184 0 _064_
rlabel via2 20194 33099 20194 33099 0 _065_
rlabel metal1 19228 36754 19228 36754 0 _066_
rlabel metal2 21850 33388 21850 33388 0 _067_
rlabel metal1 17572 33898 17572 33898 0 _068_
rlabel metal1 16836 34510 16836 34510 0 _069_
rlabel metal2 12650 33779 12650 33779 0 _070_
rlabel metal1 18538 32878 18538 32878 0 _071_
rlabel metal1 20378 34034 20378 34034 0 _072_
rlabel metal1 17710 26010 17710 26010 0 _073_
rlabel metal1 13616 25942 13616 25942 0 _074_
rlabel metal1 15318 20808 15318 20808 0 _075_
rlabel metal1 14444 18394 14444 18394 0 _076_
rlabel metal1 20056 21658 20056 21658 0 _077_
rlabel metal2 17250 20638 17250 20638 0 _078_
rlabel metal1 15870 25976 15870 25976 0 _079_
rlabel metal3 12742 25772 12742 25772 0 _080_
rlabel metal1 16376 27030 16376 27030 0 _081_
rlabel metal1 13754 23766 13754 23766 0 _082_
rlabel metal1 20010 24106 20010 24106 0 _083_
rlabel metal1 14490 27336 14490 27336 0 _084_
rlabel metal1 9016 23834 9016 23834 0 _085_
rlabel metal2 14582 17442 14582 17442 0 _086_
rlabel metal1 15364 19754 15364 19754 0 _087_
rlabel metal1 10350 20774 10350 20774 0 _088_
rlabel metal1 12926 18394 12926 18394 0 _089_
rlabel metal1 9131 24650 9131 24650 0 _090_
rlabel metal1 14720 22746 14720 22746 0 _091_
rlabel metal1 19182 24854 19182 24854 0 _092_
rlabel metal2 8510 24242 8510 24242 0 _093_
rlabel metal2 11086 19992 11086 19992 0 _094_
rlabel metal1 16100 20502 16100 20502 0 _095_
rlabel metal2 13754 27710 13754 27710 0 _096_
rlabel metal1 17250 32198 17250 32198 0 _097_
rlabel metal1 14076 31382 14076 31382 0 _098_
rlabel metal1 10212 21114 10212 21114 0 _099_
rlabel metal1 16836 26554 16836 26554 0 _100_
rlabel metal1 13432 18394 13432 18394 0 _101_
rlabel metal1 13110 21896 13110 21896 0 _102_
rlabel metal1 9752 27574 9752 27574 0 _103_
rlabel metal2 18722 29308 18722 29308 0 _104_
rlabel metal2 15502 31246 15502 31246 0 _105_
rlabel metal1 15778 29512 15778 29512 0 _106_
rlabel metal2 18906 26690 18906 26690 0 _107_
rlabel metal1 20332 29818 20332 29818 0 _108_
rlabel metal1 14582 34646 14582 34646 0 _109_
rlabel metal2 15410 34952 15410 34952 0 _110_
rlabel metal1 17434 28424 17434 28424 0 _111_
rlabel metal1 20194 31450 20194 31450 0 _112_
rlabel metal2 14122 33694 14122 33694 0 _113_
rlabel metal1 9522 24378 9522 24378 0 _114_
rlabel metal1 18078 28118 18078 28118 0 _115_
rlabel metal1 20010 28730 20010 28730 0 _116_
rlabel metal1 18768 33558 18768 33558 0 _117_
rlabel metal1 16790 32810 16790 32810 0 _118_
rlabel metal1 21114 29274 21114 29274 0 _119_
rlabel metal1 20240 28594 20240 28594 0 _120_
rlabel metal1 16928 34646 16928 34646 0 _121_
rlabel metal1 15686 34510 15686 34510 0 _122_
rlabel metal2 17066 21760 17066 21760 0 _123_
rlabel metal1 20010 24242 20010 24242 0 _124_
rlabel metal2 21390 25534 21390 25534 0 _125_
rlabel metal1 14122 27574 14122 27574 0 _126_
rlabel metal1 20746 27030 20746 27030 0 _127_
rlabel metal1 15088 23222 15088 23222 0 _128_
rlabel metal1 16192 34918 16192 34918 0 _129_
rlabel metal1 12558 23800 12558 23800 0 _130_
rlabel metal2 15410 25432 15410 25432 0 _131_
rlabel metal1 18906 28730 18906 28730 0 _132_
rlabel metal1 13754 29614 13754 29614 0 _133_
rlabel via2 14030 30379 14030 30379 0 _134_
rlabel metal1 16238 20026 16238 20026 0 _135_
rlabel metal1 21620 24106 21620 24106 0 _136_
rlabel metal1 14306 19448 14306 19448 0 _137_
rlabel metal1 16376 21590 16376 21590 0 _138_
rlabel metal2 12466 24514 12466 24514 0 _139_
rlabel metal1 18308 23222 18308 23222 0 _140_
rlabel metal1 16514 24072 16514 24072 0 _141_
rlabel metal1 20378 25160 20378 25160 0 _142_
rlabel metal1 12512 22134 12512 22134 0 _143_
rlabel metal2 17710 23851 17710 23851 0 _144_
rlabel metal1 15410 30124 15410 30124 0 _145_
rlabel metal1 14720 32742 14720 32742 0 _146_
rlabel metal1 19366 23766 19366 23766 0 _147_
rlabel metal2 18078 23528 18078 23528 0 _148_
rlabel metal2 20746 26554 20746 26554 0 _149_
rlabel metal1 15778 23290 15778 23290 0 _150_
rlabel metal1 13846 26350 13846 26350 0 _151_
rlabel metal1 17296 26010 17296 26010 0 _152_
rlabel metal1 18078 29206 18078 29206 0 _153_
rlabel metal1 12374 21624 12374 21624 0 _154_
rlabel metal1 12926 22746 12926 22746 0 _155_
rlabel metal1 14122 28458 14122 28458 0 _156_
rlabel metal1 16376 33558 16376 33558 0 _157_
rlabel metal1 14260 31110 14260 31110 0 _158_
rlabel metal1 21206 26010 21206 26010 0 _159_
rlabel metal2 22678 26792 22678 26792 0 _160_
rlabel metal2 12558 25704 12558 25704 0 _161_
rlabel metal2 13570 19618 13570 19618 0 _162_
rlabel metal2 23322 26792 23322 26792 0 _163_
rlabel metal1 22954 25942 22954 25942 0 _164_
rlabel metal1 17894 32504 17894 32504 0 _165_
rlabel metal1 19688 26282 19688 26282 0 _166_
rlabel metal2 15410 21216 15410 21216 0 _167_
rlabel metal1 15594 22678 15594 22678 0 _168_
rlabel metal1 9614 21862 9614 21862 0 _169_
rlabel metal1 7360 24650 7360 24650 0 _170_
rlabel metal1 10534 20026 10534 20026 0 _171_
rlabel metal2 8694 22882 8694 22882 0 _172_
rlabel metal2 11454 19516 11454 19516 0 _173_
rlabel metal1 9798 21590 9798 21590 0 _174_
rlabel metal2 7958 25364 7958 25364 0 _175_
rlabel metal1 10626 25976 10626 25976 0 _176_
rlabel metal1 7590 24718 7590 24718 0 _177_
rlabel metal1 12949 28118 12949 28118 0 _178_
rlabel metal1 13202 18938 13202 18938 0 _179_
rlabel metal2 12466 26792 12466 26792 0 _180_
rlabel metal1 9292 27098 9292 27098 0 _181_
rlabel metal1 11040 23630 11040 23630 0 _182_
rlabel metal1 13938 30226 13938 30226 0 _183_
rlabel metal2 12558 23766 12558 23766 0 _184_
rlabel metal2 13202 29784 13202 29784 0 _185_
rlabel metal1 10304 22950 10304 22950 0 _186_
rlabel metal1 13202 24072 13202 24072 0 _187_
rlabel metal1 11914 19720 11914 19720 0 _188_
rlabel metal1 9154 25670 9154 25670 0 _189_
rlabel metal1 14398 29546 14398 29546 0 _190_
rlabel metal1 11776 22678 11776 22678 0 _191_
rlabel metal2 16422 28016 16422 28016 0 _192_
rlabel metal1 15686 31722 15686 31722 0 _193_
rlabel metal1 19826 33558 19826 33558 0 _194_
rlabel metal1 18630 26010 18630 26010 0 _195_
rlabel metal2 13754 29614 13754 29614 0 _196_
rlabel metal1 18446 24922 18446 24922 0 _197_
rlabel metal2 15778 30158 15778 30158 0 _198_
rlabel metal2 15502 33966 15502 33966 0 _199_
rlabel metal1 10902 26282 10902 26282 0 _200_
rlabel metal1 10626 24310 10626 24310 0 _201_
rlabel metal2 38226 26673 38226 26673 0 bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal2 38226 37179 38226 37179 0 bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal1 38456 36346 38456 36346 0 bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal2 38042 1792 38042 1792 0 bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal2 38226 19737 38226 19737 0 bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_
rlabel metal1 35604 37094 35604 37094 0 bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_
rlabel metal3 1188 3468 1188 3468 0 bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_
rlabel metal3 1188 19108 1188 19108 0 bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_
rlabel metal2 31786 1989 31786 1989 0 ccff_head
rlabel metal2 38226 12461 38226 12461 0 ccff_tail
rlabel metal1 20838 37230 20838 37230 0 chanx_left_in[0]
rlabel metal1 2944 21114 2944 21114 0 chanx_left_in[10]
rlabel metal1 37490 2414 37490 2414 0 chanx_left_in[11]
rlabel metal1 14950 2346 14950 2346 0 chanx_left_in[12]
rlabel via2 1610 4811 1610 4811 0 chanx_left_in[13]
rlabel metal2 38226 33439 38226 33439 0 chanx_left_in[14]
rlabel metal1 14490 37298 14490 37298 0 chanx_left_in[15]
rlabel metal3 1556 38828 1556 38828 0 chanx_left_in[16]
rlabel via2 23690 33371 23690 33371 0 chanx_left_in[17]
rlabel metal2 38226 5559 38226 5559 0 chanx_left_in[18]
rlabel metal1 9752 2414 9752 2414 0 chanx_left_in[1]
rlabel via2 38318 28645 38318 28645 0 chanx_left_in[2]
rlabel metal1 16928 37230 16928 37230 0 chanx_left_in[3]
rlabel metal2 38226 32215 38226 32215 0 chanx_left_in[4]
rlabel metal1 1748 22066 1748 22066 0 chanx_left_in[5]
rlabel metal1 23920 37434 23920 37434 0 chanx_left_in[6]
rlabel metal2 38318 29903 38318 29903 0 chanx_left_in[7]
rlabel metal2 46 38430 46 38430 0 chanx_left_in[8]
rlabel metal2 1702 2227 1702 2227 0 chanx_left_in[9]
rlabel metal3 1188 15708 1188 15708 0 chanx_left_out[0]
rlabel metal2 8418 1520 8418 1520 0 chanx_left_out[10]
rlabel metal1 19228 37094 19228 37094 0 chanx_left_out[11]
rlabel metal1 15594 37094 15594 37094 0 chanx_left_out[12]
rlabel metal2 38226 8857 38226 8857 0 chanx_left_out[13]
rlabel metal1 25346 37094 25346 37094 0 chanx_left_out[14]
rlabel metal1 27232 37094 27232 37094 0 chanx_left_out[15]
rlabel metal2 34822 1520 34822 1520 0 chanx_left_out[16]
rlabel metal3 1188 17748 1188 17748 0 chanx_left_out[17]
rlabel via2 38226 35445 38226 35445 0 chanx_left_out[18]
rlabel metal2 25162 1520 25162 1520 0 chanx_left_out[1]
rlabel metal3 1188 21148 1188 21148 0 chanx_left_out[2]
rlabel metal2 35834 2193 35834 2193 0 chanx_left_out[3]
rlabel metal2 38226 15793 38226 15793 0 chanx_left_out[4]
rlabel metal2 4554 1520 4554 1520 0 chanx_left_out[5]
rlabel metal3 1188 13668 1188 13668 0 chanx_left_out[6]
rlabel metal3 1188 31348 1188 31348 0 chanx_left_out[7]
rlabel metal2 28382 1520 28382 1520 0 chanx_left_out[8]
rlabel metal3 1188 29988 1188 29988 0 chanx_left_out[9]
rlabel metal2 15226 35207 15226 35207 0 chanx_right_in[0]
rlabel metal1 3312 2278 3312 2278 0 chanx_right_in[10]
rlabel metal1 11730 2346 11730 2346 0 chanx_right_in[11]
rlabel metal1 33672 2346 33672 2346 0 chanx_right_in[12]
rlabel via2 38318 14365 38318 14365 0 chanx_right_in[13]
rlabel metal3 38740 6868 38740 6868 0 chanx_right_in[14]
rlabel metal3 1142 6868 1142 6868 0 chanx_right_in[15]
rlabel via2 25346 35581 25346 35581 0 chanx_right_in[16]
rlabel metal1 37628 2822 37628 2822 0 chanx_right_in[17]
rlabel via2 1702 8891 1702 8891 0 chanx_right_in[18]
rlabel metal2 38226 10999 38226 10999 0 chanx_right_in[1]
rlabel metal2 1610 24667 1610 24667 0 chanx_right_in[2]
rlabel metal1 29716 2414 29716 2414 0 chanx_right_in[3]
rlabel metal2 38318 24633 38318 24633 0 chanx_right_in[4]
rlabel metal2 13294 36295 13294 36295 0 chanx_right_in[5]
rlabel metal1 4232 35598 4232 35598 0 chanx_right_in[6]
rlabel metal1 18170 2346 18170 2346 0 chanx_right_in[7]
rlabel metal2 2438 1836 2438 1836 0 chanx_right_in[8]
rlabel metal1 23368 2346 23368 2346 0 chanx_right_in[9]
rlabel metal2 12282 37784 12282 37784 0 chanx_right_out[0]
rlabel metal1 22172 37094 22172 37094 0 chanx_right_out[10]
rlabel metal1 33672 37094 33672 37094 0 chanx_right_out[11]
rlabel metal3 1188 26588 1188 26588 0 chanx_right_out[12]
rlabel metal3 1188 22508 1188 22508 0 chanx_right_out[13]
rlabel metal2 1334 1520 1334 1520 0 chanx_right_out[14]
rlabel metal1 37582 37094 37582 37094 0 chanx_right_out[15]
rlabel metal1 29072 37094 29072 37094 0 chanx_right_out[16]
rlabel metal2 16790 1520 16790 1520 0 chanx_right_out[17]
rlabel metal2 36754 38131 36754 38131 0 chanx_right_out[18]
rlabel metal2 38226 3417 38226 3417 0 chanx_right_out[1]
rlabel metal3 1188 10268 1188 10268 0 chanx_right_out[2]
rlabel metal2 38226 21233 38226 21233 0 chanx_right_out[3]
rlabel metal2 6486 1520 6486 1520 0 chanx_right_out[4]
rlabel metal2 12926 1520 12926 1520 0 chanx_right_out[5]
rlabel metal2 20010 1520 20010 1520 0 chanx_right_out[6]
rlabel metal2 38226 23341 38226 23341 0 chanx_right_out[7]
rlabel metal2 21298 823 21298 823 0 chanx_right_out[8]
rlabel metal1 32384 37094 32384 37094 0 chanx_right_out[9]
rlabel metal1 16882 29138 16882 29138 0 mem_bottom_ipin_0.DFFR_0_.Q
rlabel metal1 15364 19346 15364 19346 0 mem_bottom_ipin_0.DFFR_1_.Q
rlabel metal1 20148 21522 20148 21522 0 mem_bottom_ipin_0.DFFR_2_.Q
rlabel metal1 3818 31858 3818 31858 0 mem_bottom_ipin_0.DFFR_3_.Q
rlabel metal1 7636 28934 7636 28934 0 mem_bottom_ipin_0.DFFR_4_.Q
rlabel metal1 6026 31110 6026 31110 0 mem_bottom_ipin_0.DFFR_5_.Q
rlabel metal1 14030 20026 14030 20026 0 mem_bottom_ipin_1.DFFR_0_.Q
rlabel metal1 8602 24786 8602 24786 0 mem_bottom_ipin_1.DFFR_1_.Q
rlabel metal2 13938 17748 13938 17748 0 mem_bottom_ipin_1.DFFR_2_.Q
rlabel metal1 5290 35734 5290 35734 0 mem_bottom_ipin_1.DFFR_3_.Q
rlabel metal2 3588 32300 3588 32300 0 mem_bottom_ipin_1.DFFR_4_.Q
rlabel metal1 6614 34374 6614 34374 0 mem_bottom_ipin_1.DFFR_5_.Q
rlabel metal1 8556 34510 8556 34510 0 mem_bottom_ipin_2.DFFR_0_.Q
rlabel metal1 18308 25874 18308 25874 0 mem_bottom_ipin_2.DFFR_1_.Q
rlabel metal1 10902 27982 10902 27982 0 mem_bottom_ipin_2.DFFR_2_.Q
rlabel metal1 14352 35666 14352 35666 0 mem_bottom_ipin_2.DFFR_3_.Q
rlabel metal2 1978 35258 1978 35258 0 mem_bottom_ipin_2.DFFR_4_.Q
rlabel metal2 8142 35632 8142 35632 0 mem_bottom_ipin_2.DFFR_5_.Q
rlabel metal1 23368 32198 23368 32198 0 mem_top_ipin_0.DFFR_0_.Q
rlabel metal2 13018 18224 13018 18224 0 mem_top_ipin_0.DFFR_1_.Q
rlabel metal1 16146 26316 16146 26316 0 mem_top_ipin_0.DFFR_2_.Q
rlabel metal1 1794 36040 1794 36040 0 mem_top_ipin_0.DFFR_3_.Q
rlabel metal2 24610 34782 24610 34782 0 mem_top_ipin_0.DFFR_4_.Q
rlabel metal2 6762 37009 6762 37009 0 mem_top_ipin_0.DFFR_5_.Q
rlabel metal1 20838 34612 20838 34612 0 mem_top_ipin_1.DFFR_0_.Q
rlabel metal1 16146 28118 16146 28118 0 mem_top_ipin_1.DFFR_1_.Q
rlabel metal2 20562 36992 20562 36992 0 mem_top_ipin_1.DFFR_2_.Q
rlabel metal1 9338 37128 9338 37128 0 mem_top_ipin_1.DFFR_3_.Q
rlabel metal1 14398 36618 14398 36618 0 mem_top_ipin_1.DFFR_4_.Q
rlabel metal1 12466 36210 12466 36210 0 mem_top_ipin_1.DFFR_5_.Q
rlabel metal1 23230 32742 23230 32742 0 mem_top_ipin_2.DFFR_0_.Q
rlabel metal2 21390 27472 21390 27472 0 mem_top_ipin_2.DFFR_1_.Q
rlabel metal1 20608 24174 20608 24174 0 mem_top_ipin_2.DFFR_2_.Q
rlabel metal1 13340 34510 13340 34510 0 mem_top_ipin_2.DFFR_3_.Q
rlabel metal2 12834 35530 12834 35530 0 mem_top_ipin_2.DFFR_4_.Q
rlabel metal1 13110 35224 13110 35224 0 mem_top_ipin_2.DFFR_5_.Q
rlabel metal1 18308 21862 18308 21862 0 mem_top_ipin_3.DFFR_0_.Q
rlabel metal1 17204 19210 17204 19210 0 mem_top_ipin_3.DFFR_1_.Q
rlabel metal1 17250 21556 17250 21556 0 mem_top_ipin_3.DFFR_2_.Q
rlabel metal1 2208 29682 2208 29682 0 mem_top_ipin_3.DFFR_3_.Q
rlabel metal1 3542 29682 3542 29682 0 mem_top_ipin_3.DFFR_4_.Q
rlabel metal1 9384 32334 9384 32334 0 mem_top_ipin_3.DFFR_5_.Q
rlabel metal1 13018 22542 13018 22542 0 mem_top_ipin_4.DFFR_0_.Q
rlabel metal2 20654 24786 20654 24786 0 mem_top_ipin_4.DFFR_1_.Q
rlabel metal1 18170 21046 18170 21046 0 mem_top_ipin_4.DFFR_2_.Q
rlabel metal1 1978 36822 1978 36822 0 mem_top_ipin_4.DFFR_3_.Q
rlabel metal1 23828 34986 23828 34986 0 mem_top_ipin_4.DFFR_4_.Q
rlabel metal1 13662 32980 13662 32980 0 mem_top_ipin_4.DFFR_5_.Q
rlabel metal1 18952 20570 18952 20570 0 mem_top_ipin_5.DFFR_0_.Q
rlabel metal1 21482 25908 21482 25908 0 mem_top_ipin_5.DFFR_1_.Q
rlabel metal2 22770 37570 22770 37570 0 mem_top_ipin_5.DFFR_2_.Q
rlabel metal1 13570 32912 13570 32912 0 mem_top_ipin_5.DFFR_3_.Q
rlabel via2 12926 37077 12926 37077 0 mem_top_ipin_5.DFFR_4_.Q
rlabel metal2 8694 34408 8694 34408 0 mem_top_ipin_5.DFFR_5_.Q
rlabel metal2 13570 18530 13570 18530 0 mem_top_ipin_6.DFFR_0_.Q
rlabel metal2 20102 34068 20102 34068 0 mem_top_ipin_6.DFFR_1_.Q
rlabel metal1 8694 21522 8694 21522 0 mem_top_ipin_6.DFFR_2_.Q
rlabel metal1 4278 29512 4278 29512 0 mem_top_ipin_6.DFFR_3_.Q
rlabel metal1 4961 34374 4961 34374 0 mem_top_ipin_6.DFFR_4_.Q
rlabel metal1 6532 33898 6532 33898 0 mem_top_ipin_6.DFFR_5_.Q
rlabel metal1 15272 32878 15272 32878 0 mem_top_ipin_7.DFFR_0_.Q
rlabel metal2 10994 25568 10994 25568 0 mem_top_ipin_7.DFFR_1_.Q
rlabel metal2 17986 35139 17986 35139 0 mem_top_ipin_7.DFFR_2_.Q
rlabel metal1 3910 34918 3910 34918 0 mem_top_ipin_7.DFFR_3_.Q
rlabel metal1 8924 33558 8924 33558 0 mem_top_ipin_7.DFFR_4_.Q
rlabel metal1 15042 28594 15042 28594 0 mux_bottom_ipin_0.INVTX1_0_.out
rlabel metal2 7222 25534 7222 25534 0 mux_bottom_ipin_0.INVTX1_1_.out
rlabel metal2 17618 27676 17618 27676 0 mux_bottom_ipin_0.INVTX1_2_.out
rlabel metal1 12558 23630 12558 23630 0 mux_bottom_ipin_0.INVTX1_3_.out
rlabel metal2 14214 19890 14214 19890 0 mux_bottom_ipin_0.INVTX1_4_.out
rlabel metal2 15686 21216 15686 21216 0 mux_bottom_ipin_0.INVTX1_5_.out
rlabel metal1 20516 24718 20516 24718 0 mux_bottom_ipin_0.INVTX1_6_.out
rlabel metal1 18124 22066 18124 22066 0 mux_bottom_ipin_0.INVTX1_7_.out
rlabel metal1 16376 26962 16376 26962 0 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 14582 20978 14582 20978 0 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 20424 24650 20424 24650 0 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 20516 9622 20516 9622 0 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 12926 20332 12926 20332 0 mux_bottom_ipin_1.INVTX1_2_.out
rlabel metal1 19918 16558 19918 16558 0 mux_bottom_ipin_1.INVTX1_3_.out
rlabel metal2 22678 25636 22678 25636 0 mux_bottom_ipin_1.INVTX1_4_.out
rlabel metal1 15318 21930 15318 21930 0 mux_bottom_ipin_1.INVTX1_5_.out
rlabel metal1 11178 20366 11178 20366 0 mux_bottom_ipin_1.INVTX1_6_.out
rlabel metal1 16008 19890 16008 19890 0 mux_bottom_ipin_1.INVTX1_7_.out
rlabel metal1 12190 25160 12190 25160 0 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 17204 23154 17204 23154 0 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 14858 18734 14858 18734 0 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 10258 19652 10258 19652 0 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 15088 29070 15088 29070 0 mux_bottom_ipin_2.INVTX1_2_.out
rlabel metal2 9154 25636 9154 25636 0 mux_bottom_ipin_2.INVTX1_3_.out
rlabel metal1 21068 26418 21068 26418 0 mux_bottom_ipin_2.INVTX1_4_.out
rlabel metal1 13846 29240 13846 29240 0 mux_bottom_ipin_2.INVTX1_5_.out
rlabel metal3 15686 32028 15686 32028 0 mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 15134 28934 15134 28934 0 mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 19826 33082 19826 33082 0 mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 18814 30158 18814 30158 0 mux_top_ipin_0.INVTX1_2_.out
rlabel metal1 21620 11866 21620 11866 0 mux_top_ipin_0.INVTX1_3_.out
rlabel metal2 12650 20094 12650 20094 0 mux_top_ipin_0.INVTX1_4_.out
rlabel via1 13018 21947 13018 21947 0 mux_top_ipin_0.INVTX1_5_.out
rlabel metal1 14674 36006 14674 36006 0 mux_top_ipin_0.INVTX1_6_.out
rlabel metal1 11086 21896 11086 21896 0 mux_top_ipin_0.INVTX1_7_.out
rlabel metal1 15364 27914 15364 27914 0 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 13754 21471 13754 21471 0 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 16376 29546 16376 29546 0 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 21390 30770 21390 30770 0 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 21160 29206 21160 29206 0 mux_top_ipin_1.INVTX1_2_.out
rlabel metal2 20286 28101 20286 28101 0 mux_top_ipin_1.INVTX1_3_.out
rlabel metal1 14030 32300 14030 32300 0 mux_top_ipin_1.INVTX1_4_.out
rlabel metal1 9982 10234 9982 10234 0 mux_top_ipin_1.INVTX1_5_.out
rlabel metal2 16514 34204 16514 34204 0 mux_top_ipin_1.INVTX1_6_.out
rlabel metal1 15088 33286 15088 33286 0 mux_top_ipin_1.INVTX1_7_.out
rlabel metal1 19274 33388 19274 33388 0 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 20010 34918 20010 34918 0 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 18584 31858 18584 31858 0 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 32108 36754 32108 36754 0 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 13110 26520 13110 26520 0 mux_top_ipin_2.INVTX1_2_.out
rlabel metal1 9453 24786 9453 24786 0 mux_top_ipin_2.INVTX1_3_.out
rlabel metal1 14214 23290 14214 23290 0 mux_top_ipin_2.INVTX1_6_.out
rlabel metal2 15502 21080 15502 21080 0 mux_top_ipin_2.INVTX1_7_.out
rlabel metal1 19734 26792 19734 26792 0 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 16836 31858 16836 31858 0 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 14214 21454 14214 21454 0 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 34362 36482 34362 36482 0 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 16146 24106 16146 24106 0 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 15042 20366 15042 20366 0 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 19550 22712 19550 22712 0 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 32660 6290 32660 6290 0 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 17112 29070 17112 29070 0 mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 19550 29682 19550 29682 0 mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 12834 21216 12834 21216 0 mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 21252 30226 21252 30226 0 mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 10902 25806 10902 25806 0 mux_top_ipin_5.INVTX1_4_.out
rlabel metal1 12834 20978 12834 20978 0 mux_top_ipin_5.INVTX1_5_.out
rlabel metal1 19458 26452 19458 26452 0 mux_top_ipin_5.INVTX1_6_.out
rlabel metal1 20056 27506 20056 27506 0 mux_top_ipin_5.INVTX1_7_.out
rlabel metal1 22862 32266 22862 32266 0 mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 14168 19890 14168 19890 0 mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 20194 31382 20194 31382 0 mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 26220 35700 26220 35700 0 mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 11178 26418 11178 26418 0 mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 11960 20774 11960 20774 0 mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 10396 27030 10396 27030 0 mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 6831 6766 6831 6766 0 mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 12466 27370 12466 27370 0 mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 11086 27370 11086 27370 0 mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 14674 29886 14674 29886 0 mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 7314 19856 7314 19856 0 mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 26220 37332 26220 37332 0 net1
rlabel metal1 15548 12206 15548 12206 0 net10
rlabel metal1 12282 24684 12282 24684 0 net100
rlabel metal1 19320 33558 19320 33558 0 net101
rlabel metal1 37996 5814 37996 5814 0 net11
rlabel metal1 13110 3026 13110 3026 0 net12
rlabel metal2 38042 28764 38042 28764 0 net13
rlabel metal2 16836 36652 16836 36652 0 net14
rlabel metal1 19412 12954 19412 12954 0 net15
rlabel via2 12742 10251 12742 10251 0 net16
rlabel metal1 20102 13294 20102 13294 0 net17
rlabel metal1 37950 30158 37950 30158 0 net18
rlabel metal1 10074 24786 10074 24786 0 net19
rlabel metal1 17066 36720 17066 36720 0 net2
rlabel metal1 6716 2890 6716 2890 0 net20
rlabel metal1 5934 18938 5934 18938 0 net21
rlabel metal2 8602 2754 8602 2754 0 net22
rlabel metal3 11431 2652 11431 2652 0 net23
rlabel metal1 19872 19890 19872 19890 0 net24
rlabel metal1 37950 12206 37950 12206 0 net25
rlabel metal1 37904 7446 37904 7446 0 net26
rlabel metal2 20010 21488 20010 21488 0 net27
rlabel metal1 25392 17170 25392 17170 0 net28
rlabel metal1 19826 19754 19826 19754 0 net29
rlabel metal1 15456 36754 15456 36754 0 net3
rlabel metal1 18078 21522 18078 21522 0 net30
rlabel metal1 24196 6766 24196 6766 0 net31
rlabel metal2 1978 24174 1978 24174 0 net32
rlabel metal1 24748 11730 24748 11730 0 net33
rlabel metal1 37996 24718 37996 24718 0 net34
rlabel metal1 9384 36142 9384 36142 0 net35
rlabel metal1 4232 21998 4232 21998 0 net36
rlabel metal1 17434 2618 17434 2618 0 net37
rlabel metal1 20332 3026 20332 3026 0 net38
rlabel metal2 23322 11254 23322 11254 0 net39
rlabel metal2 37582 13328 37582 13328 0 net4
rlabel metal2 30682 37060 30682 37060 0 net40
rlabel metal2 36662 27982 36662 27982 0 net41
rlabel metal1 36961 36754 36961 36754 0 net42
rlabel metal2 34454 36346 34454 36346 0 net43
rlabel metal2 34546 4590 34546 4590 0 net44
rlabel metal2 36570 22202 36570 22202 0 net45
rlabel metal1 31602 36822 31602 36822 0 net46
rlabel metal1 2346 3502 2346 3502 0 net47
rlabel metal2 1886 19516 1886 19516 0 net48
rlabel via2 37490 12733 37490 12733 0 net49
rlabel metal2 14674 18938 14674 18938 0 net5
rlabel metal2 4002 17340 4002 17340 0 net50
rlabel metal2 8326 2618 8326 2618 0 net51
rlabel metal2 19550 35649 19550 35649 0 net52
rlabel via3 15893 35972 15893 35972 0 net53
rlabel metal2 38042 10506 38042 10506 0 net54
rlabel metal1 24288 37162 24288 37162 0 net55
rlabel metal2 16054 21658 16054 21658 0 net56
rlabel metal1 34960 3162 34960 3162 0 net57
rlabel metal1 2162 18258 2162 18258 0 net58
rlabel metal1 37766 35666 37766 35666 0 net59
rlabel metal2 1794 6119 1794 6119 0 net6
rlabel metal1 23874 6664 23874 6664 0 net60
rlabel metal1 1840 23494 1840 23494 0 net61
rlabel metal2 35926 2652 35926 2652 0 net62
rlabel metal1 38088 20230 38088 20230 0 net63
rlabel metal2 5566 2788 5566 2788 0 net64
rlabel metal2 5290 17884 5290 17884 0 net65
rlabel metal1 5980 26554 5980 26554 0 net66
rlabel metal2 27370 2652 27370 2652 0 net67
rlabel metal2 2070 23647 2070 23647 0 net68
rlabel metal1 13386 36108 13386 36108 0 net69
rlabel metal1 18860 20910 18860 20910 0 net7
rlabel metal1 18768 36890 18768 36890 0 net70
rlabel metal2 33626 30804 33626 30804 0 net71
rlabel metal1 1886 26894 1886 26894 0 net72
rlabel metal1 2116 22610 2116 22610 0 net73
rlabel metal1 1932 2414 1932 2414 0 net74
rlabel metal1 24886 36618 24886 36618 0 net75
rlabel metal2 28934 36924 28934 36924 0 net76
rlabel metal2 16882 7378 16882 7378 0 net77
rlabel metal1 37628 21862 37628 21862 0 net78
rlabel metal2 37490 3162 37490 3162 0 net79
rlabel metal1 14858 37196 14858 37196 0 net8
rlabel metal1 1886 10676 1886 10676 0 net80
rlabel metal2 38042 22236 38042 22236 0 net81
rlabel metal1 8740 2346 8740 2346 0 net82
rlabel metal2 13294 6154 13294 6154 0 net83
rlabel metal1 20010 13158 20010 13158 0 net84
rlabel metal2 38042 23868 38042 23868 0 net85
rlabel metal1 21712 2414 21712 2414 0 net86
rlabel metal1 32062 37230 32062 37230 0 net87
rlabel metal1 14490 36788 14490 36788 0 net88
rlabel metal1 23092 9350 23092 9350 0 net89
rlabel metal1 25760 36754 25760 36754 0 net9
rlabel metal2 3358 15436 3358 15436 0 net90
rlabel metal2 20102 22746 20102 22746 0 net91
rlabel metal1 14076 17578 14076 17578 0 net92
rlabel metal1 17526 28152 17526 28152 0 net93
rlabel metal2 20102 32096 20102 32096 0 net94
rlabel metal2 16514 25874 16514 25874 0 net95
rlabel metal2 21942 24480 21942 24480 0 net96
rlabel metal2 17342 24242 17342 24242 0 net97
rlabel metal2 21850 27064 21850 27064 0 net98
rlabel metal2 9430 23392 9430 23392 0 net99
rlabel metal1 30360 37298 30360 37298 0 pReset
rlabel metal2 22218 36482 22218 36482 0 prog_clk
rlabel metal1 14306 36652 14306 36652 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_
rlabel metal2 26450 1520 26450 1520 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_
rlabel metal3 1188 12308 1188 12308 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
