magic
tech sky130A
magscale 1 2
timestamp 1674174155
<< viali >>
rect 4524 37417 4558 37451
rect 24777 37417 24811 37451
rect 35081 37417 35115 37451
rect 9137 37281 9171 37315
rect 10609 37281 10643 37315
rect 15577 37281 15611 37315
rect 29929 37281 29963 37315
rect 1593 37213 1627 37247
rect 4261 37213 4295 37247
rect 6561 37213 6595 37247
rect 10885 37213 10919 37247
rect 11713 37213 11747 37247
rect 12541 37213 12575 37247
rect 13093 37213 13127 37247
rect 14933 37213 14967 37247
rect 17049 37213 17083 37247
rect 17509 37213 17543 37247
rect 18153 37213 18187 37247
rect 20085 37213 20119 37247
rect 22017 37213 22051 37247
rect 23489 37213 23523 37247
rect 23949 37213 23983 37247
rect 25421 37213 25455 37247
rect 27445 37213 27479 37247
rect 28457 37213 28491 37247
rect 30389 37213 30423 37247
rect 32321 37213 32355 37247
rect 33609 37213 33643 37247
rect 35725 37213 35759 37247
rect 1869 37145 1903 37179
rect 6837 37145 6871 37179
rect 16129 37145 16163 37179
rect 27997 37145 28031 37179
rect 35541 37145 35575 37179
rect 3341 37077 3375 37111
rect 6009 37077 6043 37111
rect 8309 37077 8343 37111
rect 11897 37077 11931 37111
rect 13185 37077 13219 37111
rect 14289 37077 14323 37111
rect 15117 37077 15151 37111
rect 16865 37077 16899 37111
rect 18337 37077 18371 37111
rect 20269 37077 20303 37111
rect 22201 37077 22235 37111
rect 23305 37077 23339 37111
rect 25329 37077 25363 37111
rect 27261 37077 27295 37111
rect 28641 37077 28675 37111
rect 30573 37077 30607 37111
rect 32505 37077 32539 37111
rect 33793 37077 33827 37111
rect 5273 36873 5307 36907
rect 6745 36873 6779 36907
rect 7757 36873 7791 36907
rect 11713 36873 11747 36907
rect 12449 36873 12483 36907
rect 14289 36873 14323 36907
rect 35449 36873 35483 36907
rect 36277 36873 36311 36907
rect 2973 36805 3007 36839
rect 10149 36805 10183 36839
rect 2237 36737 2271 36771
rect 2697 36737 2731 36771
rect 5457 36737 5491 36771
rect 6561 36737 6595 36771
rect 7941 36737 7975 36771
rect 11069 36737 11103 36771
rect 11897 36737 11931 36771
rect 13093 36737 13127 36771
rect 14105 36737 14139 36771
rect 16865 36737 16899 36771
rect 35633 36737 35667 36771
rect 36093 36737 36127 36771
rect 2053 36669 2087 36703
rect 4721 36669 4755 36703
rect 8401 36669 8435 36703
rect 10425 36669 10459 36703
rect 13553 36669 13587 36703
rect 14749 36669 14783 36703
rect 15301 36669 15335 36703
rect 15853 36669 15887 36703
rect 6009 36533 6043 36567
rect 10885 36533 10919 36567
rect 13001 36533 13035 36567
rect 17049 36533 17083 36567
rect 11989 36329 12023 36363
rect 13645 36329 13679 36363
rect 14841 36329 14875 36363
rect 36277 36329 36311 36363
rect 3341 36261 3375 36295
rect 15393 36261 15427 36295
rect 16589 36261 16623 36295
rect 1593 36193 1627 36227
rect 1869 36193 1903 36227
rect 4537 36193 4571 36227
rect 9137 36193 9171 36227
rect 9413 36193 9447 36227
rect 4813 36125 4847 36159
rect 5457 36125 5491 36159
rect 7941 36125 7975 36159
rect 8401 36125 8435 36159
rect 13093 36125 13127 36159
rect 36093 36125 36127 36159
rect 5365 36057 5399 36091
rect 5917 36057 5951 36091
rect 7665 36057 7699 36091
rect 11529 36057 11563 36091
rect 8493 35989 8527 36023
rect 10885 35989 10919 36023
rect 13001 35989 13035 36023
rect 14289 35989 14323 36023
rect 15945 35989 15979 36023
rect 35541 35989 35575 36023
rect 13553 35785 13587 35819
rect 14657 35785 14691 35819
rect 15209 35785 15243 35819
rect 15761 35785 15795 35819
rect 1869 35717 1903 35751
rect 9137 35717 9171 35751
rect 12357 35717 12391 35751
rect 12449 35717 12483 35751
rect 1593 35649 1627 35683
rect 9781 35649 9815 35683
rect 10609 35649 10643 35683
rect 11069 35649 11103 35683
rect 14105 35649 14139 35683
rect 36093 35649 36127 35683
rect 3985 35581 4019 35615
rect 4261 35581 4295 35615
rect 6009 35581 6043 35615
rect 7113 35581 7147 35615
rect 7389 35581 7423 35615
rect 11989 35581 12023 35615
rect 3341 35445 3375 35479
rect 6561 35445 6595 35479
rect 9965 35445 9999 35479
rect 10425 35445 10459 35479
rect 13001 35445 13035 35479
rect 35541 35445 35575 35479
rect 36277 35445 36311 35479
rect 8585 35241 8619 35275
rect 13093 35241 13127 35275
rect 14289 35241 14323 35275
rect 14841 35241 14875 35275
rect 28089 35241 28123 35275
rect 3341 35105 3375 35139
rect 5089 35105 5123 35139
rect 8033 35105 8067 35139
rect 9137 35105 9171 35139
rect 11529 35105 11563 35139
rect 11805 35105 11839 35139
rect 4445 35037 4479 35071
rect 5365 35037 5399 35071
rect 15577 35037 15611 35071
rect 27905 35037 27939 35071
rect 28641 35037 28675 35071
rect 3065 34969 3099 35003
rect 4169 34969 4203 35003
rect 6009 34969 6043 35003
rect 7757 34969 7791 35003
rect 9413 34969 9447 35003
rect 11621 34969 11655 35003
rect 1593 34901 1627 34935
rect 10885 34901 10919 34935
rect 13553 34901 13587 34935
rect 15669 34901 15703 34935
rect 16405 34901 16439 34935
rect 2237 34697 2271 34731
rect 6653 34697 6687 34731
rect 7297 34697 7331 34731
rect 14013 34697 14047 34731
rect 14657 34697 14691 34731
rect 15117 34697 15151 34731
rect 3709 34629 3743 34663
rect 11805 34629 11839 34663
rect 12725 34629 12759 34663
rect 13461 34629 13495 34663
rect 17049 34629 17083 34663
rect 1777 34561 1811 34595
rect 3985 34561 4019 34595
rect 4905 34561 4939 34595
rect 5549 34561 5583 34595
rect 6745 34561 6779 34595
rect 7389 34561 7423 34595
rect 10977 34561 11011 34595
rect 13369 34561 13403 34595
rect 1685 34493 1719 34527
rect 4721 34493 4755 34527
rect 5365 34493 5399 34527
rect 8309 34493 8343 34527
rect 9781 34493 9815 34527
rect 10057 34493 10091 34527
rect 12817 34493 12851 34527
rect 16957 34493 16991 34527
rect 17233 34493 17267 34527
rect 11069 34357 11103 34391
rect 3985 34153 4019 34187
rect 7113 34153 7147 34187
rect 7757 34153 7791 34187
rect 13001 34153 13035 34187
rect 14381 34153 14415 34187
rect 14933 34153 14967 34187
rect 15393 34153 15427 34187
rect 9137 34085 9171 34119
rect 15945 34085 15979 34119
rect 3433 34017 3467 34051
rect 6561 34017 6595 34051
rect 8401 34017 8435 34051
rect 7205 33949 7239 33983
rect 7849 33949 7883 33983
rect 8309 33949 8343 33983
rect 9689 33949 9723 33983
rect 10241 33949 10275 33983
rect 12909 33949 12943 33983
rect 13737 33949 13771 33983
rect 34897 33949 34931 33983
rect 35541 33949 35575 33983
rect 3157 33881 3191 33915
rect 4537 33881 4571 33915
rect 6285 33881 6319 33915
rect 11437 33881 11471 33915
rect 11529 33881 11563 33915
rect 12449 33881 12483 33915
rect 1685 33813 1719 33847
rect 10793 33813 10827 33847
rect 13645 33813 13679 33847
rect 34989 33813 35023 33847
rect 6653 33609 6687 33643
rect 7297 33609 7331 33643
rect 11989 33609 12023 33643
rect 14841 33609 14875 33643
rect 15301 33609 15335 33643
rect 31493 33609 31527 33643
rect 5733 33541 5767 33575
rect 10057 33541 10091 33575
rect 12541 33541 12575 33575
rect 1961 33473 1995 33507
rect 6561 33473 6595 33507
rect 7389 33473 7423 33507
rect 11897 33473 11931 33507
rect 13277 33473 13311 33507
rect 14105 33473 14139 33507
rect 31309 33473 31343 33507
rect 36093 33473 36127 33507
rect 2237 33405 2271 33439
rect 3709 33405 3743 33439
rect 6009 33405 6043 33439
rect 8309 33405 8343 33439
rect 10333 33405 10367 33439
rect 10793 33405 10827 33439
rect 36277 33337 36311 33371
rect 4261 33269 4295 33303
rect 13369 33269 13403 33303
rect 14197 33269 14231 33303
rect 5457 33065 5491 33099
rect 6101 33065 6135 33099
rect 14289 33065 14323 33099
rect 1685 32929 1719 32963
rect 1961 32929 1995 32963
rect 8585 32929 8619 32963
rect 13369 32929 13403 32963
rect 3985 32861 4019 32895
rect 4721 32861 4755 32895
rect 4813 32861 4847 32895
rect 5549 32861 5583 32895
rect 6009 32861 6043 32895
rect 10977 32861 11011 32895
rect 11437 32861 11471 32895
rect 12357 32861 12391 32895
rect 8309 32793 8343 32827
rect 10701 32793 10735 32827
rect 13553 32793 13587 32827
rect 13645 32793 13679 32827
rect 3433 32725 3467 32759
rect 4169 32725 4203 32759
rect 6837 32725 6871 32759
rect 9229 32725 9263 32759
rect 12449 32725 12483 32759
rect 36369 32725 36403 32759
rect 6653 32521 6687 32555
rect 7297 32521 7331 32555
rect 13645 32453 13679 32487
rect 14197 32453 14231 32487
rect 1777 32385 1811 32419
rect 4445 32385 4479 32419
rect 5089 32385 5123 32419
rect 5733 32385 5767 32419
rect 6561 32385 6595 32419
rect 7389 32385 7423 32419
rect 10149 32385 10183 32419
rect 12173 32385 12207 32419
rect 12817 32385 12851 32419
rect 2237 32317 2271 32351
rect 3709 32317 3743 32351
rect 3985 32317 4019 32351
rect 5825 32317 5859 32351
rect 8125 32317 8159 32351
rect 9873 32317 9907 32351
rect 13553 32317 13587 32351
rect 36093 32317 36127 32351
rect 36369 32317 36403 32351
rect 5181 32249 5215 32283
rect 10701 32249 10735 32283
rect 12265 32249 12299 32283
rect 1685 32181 1719 32215
rect 4537 32181 4571 32215
rect 12909 32181 12943 32215
rect 4077 31977 4111 32011
rect 4721 31977 4755 32011
rect 5365 31977 5399 32011
rect 9137 31977 9171 32011
rect 35909 31977 35943 32011
rect 2973 31909 3007 31943
rect 6009 31909 6043 31943
rect 8493 31909 8527 31943
rect 2421 31841 2455 31875
rect 6745 31841 6779 31875
rect 11529 31841 11563 31875
rect 13553 31841 13587 31875
rect 2145 31773 2179 31807
rect 2881 31773 2915 31807
rect 4169 31773 4203 31807
rect 4813 31773 4847 31807
rect 5273 31773 5307 31807
rect 5917 31773 5951 31807
rect 9873 31773 9907 31807
rect 9965 31773 9999 31807
rect 10793 31773 10827 31807
rect 10885 31773 10919 31807
rect 11437 31773 11471 31807
rect 12081 31773 12115 31807
rect 12817 31773 12851 31807
rect 13645 31773 13679 31807
rect 14657 31773 14691 31807
rect 14749 31773 14783 31807
rect 22753 31773 22787 31807
rect 22845 31773 22879 31807
rect 23397 31773 23431 31807
rect 36093 31773 36127 31807
rect 7021 31705 7055 31739
rect 12173 31637 12207 31671
rect 12909 31637 12943 31671
rect 6653 31433 6687 31467
rect 7297 31433 7331 31467
rect 7941 31433 7975 31467
rect 4445 31365 4479 31399
rect 12265 31365 12299 31399
rect 12817 31365 12851 31399
rect 14197 31365 14231 31399
rect 15393 31365 15427 31399
rect 15485 31365 15519 31399
rect 1961 31297 1995 31331
rect 6561 31297 6595 31331
rect 7205 31297 7239 31331
rect 7849 31297 7883 31331
rect 10793 31297 10827 31331
rect 2237 31229 2271 31263
rect 4169 31229 4203 31263
rect 8493 31229 8527 31263
rect 8769 31229 8803 31263
rect 12173 31229 12207 31263
rect 13277 31229 13311 31263
rect 14289 31229 14323 31263
rect 5917 31161 5951 31195
rect 14933 31161 14967 31195
rect 3709 31093 3743 31127
rect 10241 31093 10275 31127
rect 10885 31093 10919 31127
rect 4077 30889 4111 30923
rect 8327 30889 8361 30923
rect 9137 30889 9171 30923
rect 1869 30753 1903 30787
rect 3065 30753 3099 30787
rect 8585 30753 8619 30787
rect 10885 30753 10919 30787
rect 14381 30753 14415 30787
rect 2329 30685 2363 30719
rect 2973 30685 3007 30719
rect 5825 30685 5859 30719
rect 13277 30685 13311 30719
rect 15669 30685 15703 30719
rect 1685 30617 1719 30651
rect 5549 30617 5583 30651
rect 10609 30617 10643 30651
rect 11805 30617 11839 30651
rect 11897 30617 11931 30651
rect 12817 30617 12851 30651
rect 14473 30617 14507 30651
rect 15025 30617 15059 30651
rect 2421 30549 2455 30583
rect 6837 30549 6871 30583
rect 13369 30549 13403 30583
rect 15577 30549 15611 30583
rect 16129 30549 16163 30583
rect 3341 30345 3375 30379
rect 13461 30277 13495 30311
rect 15485 30277 15519 30311
rect 1593 30209 1627 30243
rect 4261 30209 4295 30243
rect 6561 30209 6595 30243
rect 10333 30209 10367 30243
rect 12173 30209 12207 30243
rect 12817 30209 12851 30243
rect 13369 30209 13403 30243
rect 14197 30209 14231 30243
rect 14841 30209 14875 30243
rect 36093 30209 36127 30243
rect 1869 30141 1903 30175
rect 4537 30141 4571 30175
rect 6009 30141 6043 30175
rect 7665 30141 7699 30175
rect 7941 30141 7975 30175
rect 11161 30141 11195 30175
rect 15393 30141 15427 30175
rect 16037 30141 16071 30175
rect 36369 30141 36403 30175
rect 10425 30073 10459 30107
rect 6653 30005 6687 30039
rect 9413 30005 9447 30039
rect 12081 30005 12115 30039
rect 12725 30005 12759 30039
rect 14105 30005 14139 30039
rect 14749 30005 14783 30039
rect 16957 30005 16991 30039
rect 1685 29801 1719 29835
rect 2329 29801 2363 29835
rect 4077 29801 4111 29835
rect 5273 29801 5307 29835
rect 9137 29801 9171 29835
rect 36369 29801 36403 29835
rect 4721 29733 4755 29767
rect 8585 29733 8619 29767
rect 6837 29665 6871 29699
rect 12357 29665 12391 29699
rect 13277 29665 13311 29699
rect 14381 29665 14415 29699
rect 14657 29665 14691 29699
rect 16221 29665 16255 29699
rect 1777 29597 1811 29631
rect 2237 29597 2271 29631
rect 2881 29597 2915 29631
rect 4169 29597 4203 29631
rect 4813 29597 4847 29631
rect 5825 29597 5859 29631
rect 10896 29597 10930 29631
rect 2973 29529 3007 29563
rect 7113 29529 7147 29563
rect 10609 29529 10643 29563
rect 11437 29529 11471 29563
rect 11529 29529 11563 29563
rect 13001 29529 13035 29563
rect 13093 29529 13127 29563
rect 14473 29529 14507 29563
rect 16405 29529 16439 29563
rect 16497 29529 16531 29563
rect 5917 29461 5951 29495
rect 17233 29461 17267 29495
rect 2973 29257 3007 29291
rect 5457 29257 5491 29291
rect 6009 29257 6043 29291
rect 8861 29257 8895 29291
rect 9505 29257 9539 29291
rect 6837 29189 6871 29223
rect 10241 29189 10275 29223
rect 10793 29189 10827 29223
rect 12449 29189 12483 29223
rect 13645 29189 13679 29223
rect 15209 29189 15243 29223
rect 16129 29189 16163 29223
rect 16865 29189 16899 29223
rect 17417 29189 17451 29223
rect 17509 29189 17543 29223
rect 1869 29121 1903 29155
rect 4721 29121 4755 29155
rect 6561 29121 6595 29155
rect 8769 29121 8803 29155
rect 9413 29121 9447 29155
rect 18061 29121 18095 29155
rect 1593 29053 1627 29087
rect 10149 29053 10183 29087
rect 12357 29053 12391 29087
rect 13001 29053 13035 29087
rect 13553 29053 13587 29087
rect 14565 29053 14599 29087
rect 15117 29053 15151 29087
rect 18153 29053 18187 29087
rect 8309 28985 8343 29019
rect 4463 28917 4497 28951
rect 18705 28917 18739 28951
rect 4077 28713 4111 28747
rect 4721 28713 4755 28747
rect 5825 28713 5859 28747
rect 18153 28713 18187 28747
rect 2329 28645 2363 28679
rect 8125 28577 8159 28611
rect 9413 28577 9447 28611
rect 10701 28577 10735 28611
rect 13001 28577 13035 28611
rect 13656 28589 13690 28623
rect 15301 28577 15335 28611
rect 16221 28577 16255 28611
rect 1777 28509 1811 28543
rect 2237 28509 2271 28543
rect 2881 28509 2915 28543
rect 9321 28509 9355 28543
rect 9965 28509 9999 28543
rect 14289 28509 14323 28543
rect 17417 28509 17451 28543
rect 18245 28509 18279 28543
rect 30481 28509 30515 28543
rect 2973 28441 3007 28475
rect 7849 28441 7883 28475
rect 10793 28441 10827 28475
rect 11345 28441 11379 28475
rect 11897 28441 11931 28475
rect 11989 28441 12023 28475
rect 12541 28441 12575 28475
rect 13553 28441 13587 28475
rect 15485 28441 15519 28475
rect 15577 28441 15611 28475
rect 16773 28441 16807 28475
rect 16865 28441 16899 28475
rect 30389 28441 30423 28475
rect 1685 28373 1719 28407
rect 5273 28373 5307 28407
rect 6377 28373 6411 28407
rect 10057 28373 10091 28407
rect 14381 28373 14415 28407
rect 17509 28373 17543 28407
rect 18705 28373 18739 28407
rect 2973 28169 3007 28203
rect 3617 28169 3651 28203
rect 4077 28169 4111 28203
rect 11069 28169 11103 28203
rect 11805 28169 11839 28203
rect 12357 28169 12391 28203
rect 18613 28169 18647 28203
rect 9505 28101 9539 28135
rect 13461 28101 13495 28135
rect 13553 28101 13587 28135
rect 14933 28101 14967 28135
rect 15761 28101 15795 28135
rect 16313 28101 16347 28135
rect 19717 28101 19751 28135
rect 1777 28033 1811 28067
rect 2237 28033 2271 28067
rect 2881 28033 2915 28067
rect 6561 28033 6595 28067
rect 7205 28033 7239 28067
rect 7849 28033 7883 28067
rect 8677 28033 8711 28067
rect 11161 28033 11195 28067
rect 12265 28033 12299 28067
rect 18061 28033 18095 28067
rect 18705 28033 18739 28067
rect 36093 28033 36127 28067
rect 2329 27965 2363 27999
rect 5917 27965 5951 27999
rect 9413 27965 9447 27999
rect 10057 27965 10091 27999
rect 14381 27965 14415 27999
rect 15025 27965 15059 27999
rect 15669 27965 15703 27999
rect 17233 27965 17267 27999
rect 36369 27965 36403 27999
rect 13001 27897 13035 27931
rect 1593 27829 1627 27863
rect 4905 27829 4939 27863
rect 5457 27829 5491 27863
rect 6653 27829 6687 27863
rect 7297 27829 7331 27863
rect 7941 27829 7975 27863
rect 8769 27829 8803 27863
rect 17969 27829 18003 27863
rect 19257 27829 19291 27863
rect 4077 27625 4111 27659
rect 4537 27625 4571 27659
rect 5089 27625 5123 27659
rect 18613 27625 18647 27659
rect 36369 27625 36403 27659
rect 1685 27557 1719 27591
rect 3157 27557 3191 27591
rect 11069 27557 11103 27591
rect 14933 27557 14967 27591
rect 2513 27489 2547 27523
rect 7849 27489 7883 27523
rect 8493 27489 8527 27523
rect 12357 27489 12391 27523
rect 13277 27489 13311 27523
rect 15485 27489 15519 27523
rect 16129 27489 16163 27523
rect 17969 27489 18003 27523
rect 19441 27489 19475 27523
rect 2421 27421 2455 27455
rect 3065 27421 3099 27455
rect 6561 27421 6595 27455
rect 7205 27421 7239 27455
rect 10977 27421 11011 27455
rect 11621 27421 11655 27455
rect 12265 27421 12299 27455
rect 14841 27421 14875 27455
rect 18061 27421 18095 27455
rect 18705 27421 18739 27455
rect 27261 27421 27295 27455
rect 6653 27353 6687 27387
rect 8401 27353 8435 27387
rect 9689 27353 9723 27387
rect 9781 27353 9815 27387
rect 10333 27353 10367 27387
rect 11713 27353 11747 27387
rect 13001 27353 13035 27387
rect 13093 27353 13127 27387
rect 16037 27353 16071 27387
rect 16681 27353 16715 27387
rect 17233 27353 17267 27387
rect 17325 27353 17359 27387
rect 27169 27353 27203 27387
rect 5917 27285 5951 27319
rect 7297 27285 7331 27319
rect 14381 27285 14415 27319
rect 2513 27081 2547 27115
rect 3893 27081 3927 27115
rect 4353 27081 4387 27115
rect 9137 27081 9171 27115
rect 10425 27081 10459 27115
rect 18797 27081 18831 27115
rect 36185 27081 36219 27115
rect 7757 27013 7791 27047
rect 7849 27013 7883 27047
rect 12725 27013 12759 27047
rect 12817 27013 12851 27047
rect 13829 27013 13863 27047
rect 14381 27013 14415 27047
rect 16129 27013 16163 27047
rect 16221 27013 16255 27047
rect 17049 27013 17083 27047
rect 17969 27013 18003 27047
rect 1593 26945 1627 26979
rect 2329 26945 2363 26979
rect 9045 26945 9079 26979
rect 9689 26945 9723 26979
rect 10517 26945 10551 26979
rect 11989 26945 12023 26979
rect 15025 26945 15059 26979
rect 18613 26945 18647 26979
rect 35725 26945 35759 26979
rect 36369 26945 36403 26979
rect 7205 26877 7239 26911
rect 8585 26877 8619 26911
rect 14473 26877 14507 26911
rect 15945 26877 15979 26911
rect 18061 26877 18095 26911
rect 11069 26809 11103 26843
rect 13277 26809 13311 26843
rect 1777 26741 1811 26775
rect 9781 26741 9815 26775
rect 12081 26741 12115 26775
rect 19257 26741 19291 26775
rect 1593 26537 1627 26571
rect 2237 26537 2271 26571
rect 6285 26537 6319 26571
rect 8401 26537 8435 26571
rect 15025 26469 15059 26503
rect 11437 26401 11471 26435
rect 12081 26401 12115 26435
rect 14381 26401 14415 26435
rect 15577 26401 15611 26435
rect 16589 26401 16623 26435
rect 17233 26401 17267 26435
rect 17509 26401 17543 26435
rect 19441 26401 19475 26435
rect 6193 26333 6227 26367
rect 8309 26333 8343 26367
rect 9781 26333 9815 26367
rect 10701 26333 10735 26367
rect 14289 26333 14323 26367
rect 16497 26333 16531 26367
rect 18521 26333 18555 26367
rect 7113 26265 7147 26299
rect 7665 26265 7699 26299
rect 7757 26265 7791 26299
rect 9689 26265 9723 26299
rect 10793 26265 10827 26299
rect 11529 26265 11563 26299
rect 13001 26265 13035 26299
rect 13553 26265 13587 26299
rect 13645 26265 13679 26299
rect 15485 26265 15519 26299
rect 17325 26265 17359 26299
rect 18429 26265 18463 26299
rect 19993 26197 20027 26231
rect 9137 25993 9171 26027
rect 17233 25993 17267 26027
rect 17877 25993 17911 26027
rect 12173 25925 12207 25959
rect 12265 25925 12299 25959
rect 14105 25925 14139 25959
rect 15301 25925 15335 25959
rect 18521 25925 18555 25959
rect 10241 25857 10275 25891
rect 10977 25857 11011 25891
rect 17141 25857 17175 25891
rect 17969 25857 18003 25891
rect 18613 25857 18647 25891
rect 19073 25857 19107 25891
rect 19625 25857 19659 25891
rect 13185 25789 13219 25823
rect 14013 25789 14047 25823
rect 15209 25789 15243 25823
rect 15485 25789 15519 25823
rect 10333 25721 10367 25755
rect 14565 25721 14599 25755
rect 20177 25721 20211 25755
rect 9781 25653 9815 25687
rect 11069 25653 11103 25687
rect 11069 25449 11103 25483
rect 18245 25449 18279 25483
rect 9781 25381 9815 25415
rect 12909 25381 12943 25415
rect 15209 25381 15243 25415
rect 16405 25381 16439 25415
rect 19441 25381 19475 25415
rect 12265 25313 12299 25347
rect 15761 25313 15795 25347
rect 1593 25245 1627 25279
rect 2237 25245 2271 25279
rect 10333 25245 10367 25279
rect 10977 25245 11011 25279
rect 14473 25245 14507 25279
rect 17693 25245 17727 25279
rect 18337 25245 18371 25279
rect 18797 25245 18831 25279
rect 9229 25177 9263 25211
rect 9321 25177 9355 25211
rect 10425 25177 10459 25211
rect 11621 25177 11655 25211
rect 12173 25177 12207 25211
rect 13369 25177 13403 25211
rect 13461 25177 13495 25211
rect 15669 25177 15703 25211
rect 16865 25177 16899 25211
rect 16957 25177 16991 25211
rect 1777 25109 1811 25143
rect 14565 25109 14599 25143
rect 17601 25109 17635 25143
rect 9045 24905 9079 24939
rect 11805 24905 11839 24939
rect 10609 24837 10643 24871
rect 12449 24837 12483 24871
rect 16129 24837 16163 24871
rect 17417 24837 17451 24871
rect 8493 24769 8527 24803
rect 9137 24769 9171 24803
rect 9781 24769 9815 24803
rect 14289 24769 14323 24803
rect 14933 24769 14967 24803
rect 18337 24769 18371 24803
rect 18429 24769 18463 24803
rect 25881 24769 25915 24803
rect 26525 24769 26559 24803
rect 33425 24769 33459 24803
rect 35541 24769 35575 24803
rect 36093 24769 36127 24803
rect 10517 24701 10551 24735
rect 12357 24701 12391 24735
rect 13185 24701 13219 24735
rect 16221 24701 16255 24735
rect 17509 24701 17543 24735
rect 11069 24633 11103 24667
rect 15669 24633 15703 24667
rect 16957 24633 16991 24667
rect 18981 24633 19015 24667
rect 26065 24633 26099 24667
rect 33609 24633 33643 24667
rect 9873 24565 9907 24599
rect 14381 24565 14415 24599
rect 15025 24565 15059 24599
rect 19533 24565 19567 24599
rect 36277 24565 36311 24599
rect 17417 24361 17451 24395
rect 17969 24361 18003 24395
rect 28825 24361 28859 24395
rect 9965 24293 9999 24327
rect 11069 24225 11103 24259
rect 11713 24225 11747 24259
rect 12173 24225 12207 24259
rect 13645 24225 13679 24259
rect 14933 24225 14967 24259
rect 15485 24225 15519 24259
rect 18521 24225 18555 24259
rect 12357 24157 12391 24191
rect 13553 24157 13587 24191
rect 16865 24157 16899 24191
rect 17509 24157 17543 24191
rect 28917 24157 28951 24191
rect 7849 24089 7883 24123
rect 8401 24089 8435 24123
rect 8493 24089 8527 24123
rect 9413 24089 9447 24123
rect 9505 24089 9539 24123
rect 11161 24089 11195 24123
rect 14289 24089 14323 24123
rect 14841 24089 14875 24123
rect 16037 24089 16071 24123
rect 16129 24089 16163 24123
rect 12817 24021 12851 24055
rect 16773 24021 16807 24055
rect 6653 23817 6687 23851
rect 9873 23817 9907 23851
rect 11069 23817 11103 23851
rect 16865 23817 16899 23851
rect 17509 23817 17543 23851
rect 36093 23817 36127 23851
rect 10425 23749 10459 23783
rect 12265 23749 12299 23783
rect 13185 23749 13219 23783
rect 13829 23749 13863 23783
rect 15393 23749 15427 23783
rect 1869 23681 1903 23715
rect 2513 23681 2547 23715
rect 6561 23681 6595 23715
rect 7205 23681 7239 23715
rect 10333 23681 10367 23715
rect 10977 23681 11011 23715
rect 22385 23681 22419 23715
rect 35909 23681 35943 23715
rect 12173 23613 12207 23647
rect 13737 23613 13771 23647
rect 14013 23613 14047 23647
rect 15301 23613 15335 23647
rect 15577 23613 15611 23647
rect 1685 23477 1719 23511
rect 2329 23477 2363 23511
rect 22477 23477 22511 23511
rect 13461 23273 13495 23307
rect 11713 23205 11747 23239
rect 15209 23205 15243 23239
rect 10609 23137 10643 23171
rect 12265 23137 12299 23171
rect 31125 23137 31159 23171
rect 6101 23069 6135 23103
rect 12449 23069 12483 23103
rect 13369 23069 13403 23103
rect 14381 23069 14415 23103
rect 16405 23069 16439 23103
rect 17049 23069 17083 23103
rect 17601 23069 17635 23103
rect 22201 23069 22235 23103
rect 31217 23069 31251 23103
rect 11161 23001 11195 23035
rect 11253 23001 11287 23035
rect 15669 23001 15703 23035
rect 15761 23001 15795 23035
rect 16589 23001 16623 23035
rect 6009 22933 6043 22967
rect 12909 22933 12943 22967
rect 14565 22933 14599 22967
rect 1961 22729 1995 22763
rect 12357 22729 12391 22763
rect 13001 22729 13035 22763
rect 8217 22661 8251 22695
rect 9045 22661 9079 22695
rect 9597 22661 9631 22695
rect 10609 22661 10643 22695
rect 11161 22661 11195 22695
rect 13553 22661 13587 22695
rect 14749 22661 14783 22695
rect 14841 22661 14875 22695
rect 15393 22661 15427 22695
rect 2145 22593 2179 22627
rect 12265 22593 12299 22627
rect 12909 22593 12943 22627
rect 14013 22593 14047 22627
rect 16037 22593 16071 22627
rect 16865 22593 16899 22627
rect 36093 22593 36127 22627
rect 7849 22525 7883 22559
rect 8309 22525 8343 22559
rect 8953 22525 8987 22559
rect 10517 22525 10551 22559
rect 14197 22525 14231 22559
rect 15945 22525 15979 22559
rect 11713 22457 11747 22491
rect 36277 22457 36311 22491
rect 2697 22389 2731 22423
rect 9229 22185 9263 22219
rect 10885 22185 10919 22219
rect 11529 22185 11563 22219
rect 7021 22049 7055 22083
rect 12633 22049 12667 22083
rect 13645 22049 13679 22083
rect 14841 22049 14875 22083
rect 5733 21981 5767 22015
rect 6929 21981 6963 22015
rect 7573 21981 7607 22015
rect 9321 21981 9355 22015
rect 10977 21981 11011 22015
rect 11437 21981 11471 22015
rect 12541 21981 12575 22015
rect 13737 21981 13771 22015
rect 16221 21981 16255 22015
rect 16681 21981 16715 22015
rect 31953 21981 31987 22015
rect 8585 21913 8619 21947
rect 10333 21913 10367 21947
rect 15393 21913 15427 21947
rect 15485 21913 15519 21947
rect 5917 21845 5951 21879
rect 6377 21845 6411 21879
rect 14289 21845 14323 21879
rect 16129 21845 16163 21879
rect 31769 21845 31803 21879
rect 32505 21845 32539 21879
rect 12633 21641 12667 21675
rect 13277 21641 13311 21675
rect 7941 21573 7975 21607
rect 13921 21573 13955 21607
rect 15669 21573 15703 21607
rect 1869 21505 1903 21539
rect 13369 21505 13403 21539
rect 13829 21505 13863 21539
rect 36093 21505 36127 21539
rect 7389 21437 7423 21471
rect 8033 21437 8067 21471
rect 14657 21437 14691 21471
rect 15761 21437 15795 21471
rect 15209 21369 15243 21403
rect 1685 21301 1719 21335
rect 12081 21301 12115 21335
rect 36277 21301 36311 21335
rect 12173 21097 12207 21131
rect 30573 21097 30607 21131
rect 36093 21097 36127 21131
rect 13737 21029 13771 21063
rect 14749 20961 14783 20995
rect 30665 20893 30699 20927
rect 31217 20893 31251 20927
rect 35449 20893 35483 20927
rect 35909 20893 35943 20927
rect 14841 20825 14875 20859
rect 15393 20825 15427 20859
rect 13001 20757 13035 20791
rect 14381 20553 14415 20587
rect 16221 20553 16255 20587
rect 14289 20417 14323 20451
rect 14933 20417 14967 20451
rect 15577 20417 15611 20451
rect 15669 20281 15703 20315
rect 3065 20009 3099 20043
rect 8217 20009 8251 20043
rect 9229 20009 9263 20043
rect 21833 20009 21867 20043
rect 1869 19805 1903 19839
rect 2513 19805 2547 19839
rect 7665 19805 7699 19839
rect 9137 19805 9171 19839
rect 9781 19805 9815 19839
rect 21373 19805 21407 19839
rect 1685 19669 1719 19703
rect 2329 19669 2363 19703
rect 7573 19669 7607 19703
rect 21189 19669 21223 19703
rect 2513 18785 2547 18819
rect 8125 18785 8159 18819
rect 16405 18785 16439 18819
rect 1961 18717 1995 18751
rect 7481 18649 7515 18683
rect 7573 18649 7607 18683
rect 16957 18649 16991 18683
rect 17049 18649 17083 18683
rect 1777 18581 1811 18615
rect 17693 18581 17727 18615
rect 1685 18241 1719 18275
rect 1777 18037 1811 18071
rect 1593 17765 1627 17799
rect 27353 17289 27387 17323
rect 27169 17153 27203 17187
rect 27813 17153 27847 17187
rect 36093 17153 36127 17187
rect 36277 17017 36311 17051
rect 1869 16065 1903 16099
rect 13829 16065 13863 16099
rect 25421 16065 25455 16099
rect 26065 16065 26099 16099
rect 36093 16065 36127 16099
rect 36369 15997 36403 16031
rect 13645 15929 13679 15963
rect 14381 15929 14415 15963
rect 1685 15861 1719 15895
rect 25605 15861 25639 15895
rect 36369 15657 36403 15691
rect 24869 14365 24903 14399
rect 25513 14365 25547 14399
rect 31401 14365 31435 14399
rect 1685 14297 1719 14331
rect 1869 14297 1903 14331
rect 31309 14297 31343 14331
rect 25053 14229 25087 14263
rect 1685 14025 1719 14059
rect 13185 14025 13219 14059
rect 13369 13889 13403 13923
rect 13829 13889 13863 13923
rect 36093 13889 36127 13923
rect 36277 13685 36311 13719
rect 1961 13277 1995 13311
rect 1869 13141 1903 13175
rect 1869 12801 1903 12835
rect 1685 12597 1719 12631
rect 35725 11713 35759 11747
rect 36369 11713 36403 11747
rect 36185 11509 36219 11543
rect 1869 10625 1903 10659
rect 36093 10625 36127 10659
rect 36369 10557 36403 10591
rect 1685 10421 1719 10455
rect 36369 10217 36403 10251
rect 5365 9605 5399 9639
rect 5273 9537 5307 9571
rect 36001 9537 36035 9571
rect 35449 9333 35483 9367
rect 36093 9333 36127 9367
rect 1869 8993 1903 9027
rect 1593 8925 1627 8959
rect 1593 8585 1627 8619
rect 10885 8585 10919 8619
rect 15209 8585 15243 8619
rect 24501 8585 24535 8619
rect 10977 8449 11011 8483
rect 15117 8449 15151 8483
rect 15761 8449 15795 8483
rect 24593 8449 24627 8483
rect 35449 8449 35483 8483
rect 36093 8449 36127 8483
rect 35633 8313 35667 8347
rect 36277 8313 36311 8347
rect 15761 8041 15795 8075
rect 15853 7837 15887 7871
rect 1869 7361 1903 7395
rect 1685 7157 1719 7191
rect 6377 6749 6411 6783
rect 7021 6749 7055 6783
rect 6561 6613 6595 6647
rect 15025 6409 15059 6443
rect 36185 6409 36219 6443
rect 15117 6273 15151 6307
rect 15577 6273 15611 6307
rect 35725 6273 35759 6307
rect 36369 6273 36403 6307
rect 1593 5185 1627 5219
rect 2237 5185 2271 5219
rect 36093 5185 36127 5219
rect 1777 4981 1811 5015
rect 36277 4981 36311 5015
rect 36369 3893 36403 3927
rect 2329 3689 2363 3723
rect 15577 3689 15611 3723
rect 1869 3485 1903 3519
rect 2513 3485 2547 3519
rect 15117 3485 15151 3519
rect 36093 3485 36127 3519
rect 1685 3349 1719 3383
rect 14933 3349 14967 3383
rect 35541 3349 35575 3383
rect 36277 3349 36311 3383
rect 11713 3145 11747 3179
rect 12449 3145 12483 3179
rect 14473 3077 14507 3111
rect 23673 3077 23707 3111
rect 1869 3009 1903 3043
rect 3985 3009 4019 3043
rect 11897 3009 11931 3043
rect 15853 3009 15887 3043
rect 19349 3009 19383 3043
rect 19993 3009 20027 3043
rect 23029 3009 23063 3043
rect 33057 3009 33091 3043
rect 34805 3009 34839 3043
rect 36093 3009 36127 3043
rect 23121 2941 23155 2975
rect 36369 2941 36403 2975
rect 14657 2873 14691 2907
rect 33241 2873 33275 2907
rect 1685 2805 1719 2839
rect 2329 2805 2363 2839
rect 4169 2805 4203 2839
rect 10241 2805 10275 2839
rect 15669 2805 15703 2839
rect 19441 2805 19475 2839
rect 32321 2805 32355 2839
rect 34989 2805 35023 2839
rect 2513 2601 2547 2635
rect 3249 2601 3283 2635
rect 19441 2601 19475 2635
rect 20821 2601 20855 2635
rect 22201 2601 22235 2635
rect 32413 2601 32447 2635
rect 34161 2601 34195 2635
rect 10701 2533 10735 2567
rect 13737 2533 13771 2567
rect 16221 2533 16255 2567
rect 9413 2465 9447 2499
rect 24869 2465 24903 2499
rect 30021 2465 30055 2499
rect 35817 2465 35851 2499
rect 1869 2397 1903 2431
rect 2329 2397 2363 2431
rect 4629 2397 4663 2431
rect 6561 2397 6595 2431
rect 9137 2397 9171 2431
rect 11989 2397 12023 2431
rect 15209 2397 15243 2431
rect 16865 2397 16899 2431
rect 19625 2397 19659 2431
rect 20361 2397 20395 2431
rect 24593 2397 24627 2431
rect 25881 2397 25915 2431
rect 27169 2397 27203 2431
rect 29745 2397 29779 2431
rect 31033 2397 31067 2431
rect 33609 2397 33643 2431
rect 35541 2397 35575 2431
rect 3341 2329 3375 2363
rect 3985 2329 4019 2363
rect 10517 2329 10551 2363
rect 13553 2329 13587 2363
rect 14289 2329 14323 2363
rect 21465 2329 21499 2363
rect 22109 2329 22143 2363
rect 32505 2329 32539 2363
rect 34253 2329 34287 2363
rect 34897 2329 34931 2363
rect 1685 2261 1719 2295
rect 4813 2261 4847 2295
rect 6745 2261 6779 2295
rect 8493 2261 8527 2295
rect 11805 2261 11839 2295
rect 15025 2261 15059 2295
rect 17049 2261 17083 2295
rect 18797 2261 18831 2295
rect 20177 2261 20211 2295
rect 23949 2261 23983 2295
rect 26065 2261 26099 2295
rect 27353 2261 27387 2295
rect 29101 2261 29135 2295
rect 31217 2261 31251 2295
<< metal1 >>
rect 658 37612 664 37664
rect 716 37652 722 37664
rect 5166 37652 5172 37664
rect 716 37624 5172 37652
rect 716 37612 722 37624
rect 5166 37612 5172 37624
rect 5224 37612 5230 37664
rect 1104 37562 36892 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 36892 37562
rect 1104 37488 36892 37510
rect 4512 37451 4570 37457
rect 4512 37417 4524 37451
rect 4558 37448 4570 37451
rect 24765 37451 24823 37457
rect 4558 37420 9168 37448
rect 4558 37417 4570 37420
rect 4512 37411 4570 37417
rect 3418 37272 3424 37324
rect 3476 37312 3482 37324
rect 4522 37312 4528 37324
rect 3476 37284 4528 37312
rect 3476 37272 3482 37284
rect 4522 37272 4528 37284
rect 4580 37272 4586 37324
rect 9140 37321 9168 37420
rect 24765 37417 24777 37451
rect 24811 37448 24823 37451
rect 25130 37448 25136 37460
rect 24811 37420 25136 37448
rect 24811 37417 24823 37420
rect 24765 37411 24823 37417
rect 25130 37408 25136 37420
rect 25188 37408 25194 37460
rect 35069 37451 35127 37457
rect 35069 37417 35081 37451
rect 35115 37448 35127 37451
rect 35434 37448 35440 37460
rect 35115 37420 35440 37448
rect 35115 37417 35127 37420
rect 35069 37411 35127 37417
rect 35434 37408 35440 37420
rect 35492 37408 35498 37460
rect 9125 37315 9183 37321
rect 9125 37281 9137 37315
rect 9171 37312 9183 37315
rect 9306 37312 9312 37324
rect 9171 37284 9312 37312
rect 9171 37281 9183 37284
rect 9125 37275 9183 37281
rect 9306 37272 9312 37284
rect 9364 37272 9370 37324
rect 10594 37312 10600 37324
rect 10555 37284 10600 37312
rect 10594 37272 10600 37284
rect 10652 37272 10658 37324
rect 15565 37315 15623 37321
rect 15565 37312 15577 37315
rect 14936 37284 15577 37312
rect 1581 37247 1639 37253
rect 1581 37213 1593 37247
rect 1627 37213 1639 37247
rect 1581 37207 1639 37213
rect 4249 37247 4307 37253
rect 4249 37213 4261 37247
rect 4295 37213 4307 37247
rect 4249 37207 4307 37213
rect 1596 37120 1624 37207
rect 1762 37136 1768 37188
rect 1820 37176 1826 37188
rect 1857 37179 1915 37185
rect 1857 37176 1869 37179
rect 1820 37148 1869 37176
rect 1820 37136 1826 37148
rect 1857 37145 1869 37148
rect 1903 37145 1915 37179
rect 3142 37176 3148 37188
rect 3082 37148 3148 37176
rect 1857 37139 1915 37145
rect 3142 37136 3148 37148
rect 3200 37136 3206 37188
rect 4264 37176 4292 37207
rect 5626 37204 5632 37256
rect 5684 37204 5690 37256
rect 6549 37247 6607 37253
rect 6549 37244 6561 37247
rect 5828 37216 6561 37244
rect 3252 37148 4292 37176
rect 1578 37108 1584 37120
rect 1491 37080 1584 37108
rect 1578 37068 1584 37080
rect 1636 37108 1642 37120
rect 2590 37108 2596 37120
rect 1636 37080 2596 37108
rect 1636 37068 1642 37080
rect 2590 37068 2596 37080
rect 2648 37108 2654 37120
rect 3252 37108 3280 37148
rect 2648 37080 3280 37108
rect 2648 37068 2654 37080
rect 3326 37068 3332 37120
rect 3384 37108 3390 37120
rect 4264 37108 4292 37148
rect 5828 37108 5856 37216
rect 6549 37213 6561 37216
rect 6595 37213 6607 37247
rect 6549 37207 6607 37213
rect 10870 37204 10876 37256
rect 10928 37244 10934 37256
rect 11698 37244 11704 37256
rect 10928 37216 10973 37244
rect 11659 37216 11704 37244
rect 10928 37204 10934 37216
rect 11698 37204 11704 37216
rect 11756 37204 11762 37256
rect 12529 37247 12587 37253
rect 12529 37213 12541 37247
rect 12575 37244 12587 37247
rect 12894 37244 12900 37256
rect 12575 37216 12900 37244
rect 12575 37213 12587 37216
rect 12529 37207 12587 37213
rect 12894 37204 12900 37216
rect 12952 37244 12958 37256
rect 13081 37247 13139 37253
rect 13081 37244 13093 37247
rect 12952 37216 13093 37244
rect 12952 37204 12958 37216
rect 13081 37213 13093 37216
rect 13127 37213 13139 37247
rect 13081 37207 13139 37213
rect 14826 37204 14832 37256
rect 14884 37244 14890 37256
rect 14936 37253 14964 37284
rect 15565 37281 15577 37284
rect 15611 37281 15623 37315
rect 15565 37275 15623 37281
rect 29917 37315 29975 37321
rect 29917 37281 29929 37315
rect 29963 37312 29975 37315
rect 30282 37312 30288 37324
rect 29963 37284 30288 37312
rect 29963 37281 29975 37284
rect 29917 37275 29975 37281
rect 30282 37272 30288 37284
rect 30340 37312 30346 37324
rect 30340 37284 30420 37312
rect 30340 37272 30346 37284
rect 14921 37247 14979 37253
rect 14921 37244 14933 37247
rect 14884 37216 14933 37244
rect 14884 37204 14890 37216
rect 14921 37213 14933 37216
rect 14967 37213 14979 37247
rect 14921 37207 14979 37213
rect 16574 37204 16580 37256
rect 16632 37244 16638 37256
rect 17037 37247 17095 37253
rect 17037 37244 17049 37247
rect 16632 37216 17049 37244
rect 16632 37204 16638 37216
rect 17037 37213 17049 37216
rect 17083 37244 17095 37247
rect 17497 37247 17555 37253
rect 17497 37244 17509 37247
rect 17083 37216 17509 37244
rect 17083 37213 17095 37216
rect 17037 37207 17095 37213
rect 17497 37213 17509 37216
rect 17543 37213 17555 37247
rect 18138 37244 18144 37256
rect 18099 37216 18144 37244
rect 17497 37207 17555 37213
rect 18138 37204 18144 37216
rect 18196 37204 18202 37256
rect 18782 37204 18788 37256
rect 18840 37244 18846 37256
rect 20073 37247 20131 37253
rect 20073 37244 20085 37247
rect 18840 37216 20085 37244
rect 18840 37204 18846 37216
rect 20073 37213 20085 37216
rect 20119 37213 20131 37247
rect 22002 37244 22008 37256
rect 21963 37216 22008 37244
rect 20073 37207 20131 37213
rect 22002 37204 22008 37216
rect 22060 37204 22066 37256
rect 23474 37244 23480 37256
rect 23435 37216 23480 37244
rect 23474 37204 23480 37216
rect 23532 37244 23538 37256
rect 23937 37247 23995 37253
rect 23937 37244 23949 37247
rect 23532 37216 23949 37244
rect 23532 37204 23538 37216
rect 23937 37213 23949 37216
rect 23983 37213 23995 37247
rect 23937 37207 23995 37213
rect 25130 37204 25136 37256
rect 25188 37244 25194 37256
rect 25409 37247 25467 37253
rect 25409 37244 25421 37247
rect 25188 37216 25421 37244
rect 25188 37204 25194 37216
rect 25409 37213 25421 37216
rect 25455 37213 25467 37247
rect 25409 37207 25467 37213
rect 27433 37247 27491 37253
rect 27433 37213 27445 37247
rect 27479 37244 27491 37247
rect 28442 37244 28448 37256
rect 27479 37216 28028 37244
rect 28403 37216 28448 37244
rect 27479 37213 27491 37216
rect 27433 37207 27491 37213
rect 6825 37179 6883 37185
rect 6825 37176 6837 37179
rect 6656 37148 6837 37176
rect 6656 37120 6684 37148
rect 6825 37145 6837 37148
rect 6871 37145 6883 37179
rect 6825 37139 6883 37145
rect 7834 37136 7840 37188
rect 7892 37136 7898 37188
rect 8570 37136 8576 37188
rect 8628 37176 8634 37188
rect 11790 37176 11796 37188
rect 8628 37148 9430 37176
rect 10244 37148 11796 37176
rect 8628 37136 8634 37148
rect 3384 37080 3429 37108
rect 4264 37080 5856 37108
rect 5997 37111 6055 37117
rect 3384 37068 3390 37080
rect 5997 37077 6009 37111
rect 6043 37108 6055 37111
rect 6638 37108 6644 37120
rect 6043 37080 6644 37108
rect 6043 37077 6055 37080
rect 5997 37071 6055 37077
rect 6638 37068 6644 37080
rect 6696 37068 6702 37120
rect 8294 37108 8300 37120
rect 8255 37080 8300 37108
rect 8294 37068 8300 37080
rect 8352 37068 8358 37120
rect 8662 37068 8668 37120
rect 8720 37108 8726 37120
rect 10244 37108 10272 37148
rect 11790 37136 11796 37148
rect 11848 37136 11854 37188
rect 16114 37176 16120 37188
rect 16075 37148 16120 37176
rect 16114 37136 16120 37148
rect 16172 37136 16178 37188
rect 21818 37136 21824 37188
rect 21876 37176 21882 37188
rect 28000 37185 28028 37216
rect 28442 37204 28448 37216
rect 28500 37204 28506 37256
rect 30392 37253 30420 37284
rect 30377 37247 30435 37253
rect 30377 37213 30389 37247
rect 30423 37213 30435 37247
rect 30377 37207 30435 37213
rect 31478 37204 31484 37256
rect 31536 37244 31542 37256
rect 32309 37247 32367 37253
rect 32309 37244 32321 37247
rect 31536 37216 32321 37244
rect 31536 37204 31542 37216
rect 32309 37213 32321 37216
rect 32355 37213 32367 37247
rect 33594 37244 33600 37256
rect 33555 37216 33600 37244
rect 32309 37207 32367 37213
rect 33594 37204 33600 37216
rect 33652 37204 33658 37256
rect 35434 37204 35440 37256
rect 35492 37244 35498 37256
rect 35713 37247 35771 37253
rect 35713 37244 35725 37247
rect 35492 37216 35725 37244
rect 35492 37204 35498 37216
rect 35713 37213 35725 37216
rect 35759 37213 35771 37247
rect 35713 37207 35771 37213
rect 27985 37179 28043 37185
rect 21876 37148 23336 37176
rect 21876 37136 21882 37148
rect 8720 37080 10272 37108
rect 8720 37068 8726 37080
rect 11054 37068 11060 37120
rect 11112 37108 11118 37120
rect 11885 37111 11943 37117
rect 11885 37108 11897 37111
rect 11112 37080 11897 37108
rect 11112 37068 11118 37080
rect 11885 37077 11897 37080
rect 11931 37077 11943 37111
rect 13170 37108 13176 37120
rect 13131 37080 13176 37108
rect 11885 37071 11943 37077
rect 13170 37068 13176 37080
rect 13228 37068 13234 37120
rect 13538 37068 13544 37120
rect 13596 37108 13602 37120
rect 14277 37111 14335 37117
rect 14277 37108 14289 37111
rect 13596 37080 14289 37108
rect 13596 37068 13602 37080
rect 14277 37077 14289 37080
rect 14323 37077 14335 37111
rect 15102 37108 15108 37120
rect 15063 37080 15108 37108
rect 14277 37071 14335 37077
rect 15102 37068 15108 37080
rect 15160 37068 15166 37120
rect 15194 37068 15200 37120
rect 15252 37108 15258 37120
rect 16853 37111 16911 37117
rect 16853 37108 16865 37111
rect 15252 37080 16865 37108
rect 15252 37068 15258 37080
rect 16853 37077 16865 37080
rect 16899 37077 16911 37111
rect 16853 37071 16911 37077
rect 18046 37068 18052 37120
rect 18104 37108 18110 37120
rect 18325 37111 18383 37117
rect 18325 37108 18337 37111
rect 18104 37080 18337 37108
rect 18104 37068 18110 37080
rect 18325 37077 18337 37080
rect 18371 37077 18383 37111
rect 18325 37071 18383 37077
rect 19978 37068 19984 37120
rect 20036 37108 20042 37120
rect 20257 37111 20315 37117
rect 20257 37108 20269 37111
rect 20036 37080 20269 37108
rect 20036 37068 20042 37080
rect 20257 37077 20269 37080
rect 20303 37077 20315 37111
rect 20257 37071 20315 37077
rect 21266 37068 21272 37120
rect 21324 37108 21330 37120
rect 23308 37117 23336 37148
rect 27985 37145 27997 37179
rect 28031 37176 28043 37179
rect 31846 37176 31852 37188
rect 28031 37148 31852 37176
rect 28031 37145 28043 37148
rect 27985 37139 28043 37145
rect 31846 37136 31852 37148
rect 31904 37136 31910 37188
rect 35526 37176 35532 37188
rect 35487 37148 35532 37176
rect 35526 37136 35532 37148
rect 35584 37136 35590 37188
rect 22189 37111 22247 37117
rect 22189 37108 22201 37111
rect 21324 37080 22201 37108
rect 21324 37068 21330 37080
rect 22189 37077 22201 37080
rect 22235 37077 22247 37111
rect 22189 37071 22247 37077
rect 23293 37111 23351 37117
rect 23293 37077 23305 37111
rect 23339 37077 23351 37111
rect 25314 37108 25320 37120
rect 25275 37080 25320 37108
rect 23293 37071 23351 37077
rect 25314 37068 25320 37080
rect 25372 37068 25378 37120
rect 26418 37068 26424 37120
rect 26476 37108 26482 37120
rect 27249 37111 27307 37117
rect 27249 37108 27261 37111
rect 26476 37080 27261 37108
rect 26476 37068 26482 37080
rect 27249 37077 27261 37080
rect 27295 37077 27307 37111
rect 27249 37071 27307 37077
rect 28350 37068 28356 37120
rect 28408 37108 28414 37120
rect 28629 37111 28687 37117
rect 28629 37108 28641 37111
rect 28408 37080 28641 37108
rect 28408 37068 28414 37080
rect 28629 37077 28641 37080
rect 28675 37077 28687 37111
rect 30558 37108 30564 37120
rect 30519 37080 30564 37108
rect 28629 37071 28687 37077
rect 30558 37068 30564 37080
rect 30616 37068 30622 37120
rect 31754 37068 31760 37120
rect 31812 37108 31818 37120
rect 32493 37111 32551 37117
rect 32493 37108 32505 37111
rect 31812 37080 32505 37108
rect 31812 37068 31818 37080
rect 32493 37077 32505 37080
rect 32539 37077 32551 37111
rect 32493 37071 32551 37077
rect 33502 37068 33508 37120
rect 33560 37108 33566 37120
rect 33781 37111 33839 37117
rect 33781 37108 33793 37111
rect 33560 37080 33793 37108
rect 33560 37068 33566 37080
rect 33781 37077 33793 37080
rect 33827 37077 33839 37111
rect 33781 37071 33839 37077
rect 1104 37018 36892 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 36892 37018
rect 1104 36944 36892 36966
rect 4614 36864 4620 36916
rect 4672 36904 4678 36916
rect 5261 36907 5319 36913
rect 5261 36904 5273 36907
rect 4672 36876 5273 36904
rect 4672 36864 4678 36876
rect 5261 36873 5273 36876
rect 5307 36873 5319 36907
rect 5261 36867 5319 36873
rect 5810 36864 5816 36916
rect 5868 36904 5874 36916
rect 6733 36907 6791 36913
rect 6733 36904 6745 36907
rect 5868 36876 6745 36904
rect 5868 36864 5874 36876
rect 6733 36873 6745 36876
rect 6779 36873 6791 36907
rect 7742 36904 7748 36916
rect 7703 36876 7748 36904
rect 6733 36867 6791 36873
rect 7742 36864 7748 36876
rect 7800 36864 7806 36916
rect 11698 36904 11704 36916
rect 7944 36876 11008 36904
rect 11659 36876 11704 36904
rect 2958 36836 2964 36848
rect 2919 36808 2964 36836
rect 2958 36796 2964 36808
rect 3016 36796 3022 36848
rect 6822 36836 6828 36848
rect 4186 36808 6828 36836
rect 6822 36796 6828 36808
rect 6880 36796 6886 36848
rect 2222 36768 2228 36780
rect 2183 36740 2228 36768
rect 2222 36728 2228 36740
rect 2280 36728 2286 36780
rect 2590 36728 2596 36780
rect 2648 36768 2654 36780
rect 2685 36771 2743 36777
rect 2685 36768 2697 36771
rect 2648 36740 2697 36768
rect 2648 36728 2654 36740
rect 2685 36737 2697 36740
rect 2731 36737 2743 36771
rect 2685 36731 2743 36737
rect 5445 36771 5503 36777
rect 5445 36737 5457 36771
rect 5491 36768 5503 36771
rect 6546 36768 6552 36780
rect 5491 36740 6408 36768
rect 6507 36740 6552 36768
rect 5491 36737 5503 36740
rect 5445 36731 5503 36737
rect 2041 36703 2099 36709
rect 2041 36669 2053 36703
rect 2087 36700 2099 36703
rect 4706 36700 4712 36712
rect 2087 36672 4568 36700
rect 4667 36672 4712 36700
rect 2087 36669 2099 36672
rect 2041 36663 2099 36669
rect 4540 36632 4568 36672
rect 4706 36660 4712 36672
rect 4764 36660 4770 36712
rect 4890 36632 4896 36644
rect 4540 36604 4896 36632
rect 4890 36592 4896 36604
rect 4948 36592 4954 36644
rect 6380 36632 6408 36740
rect 6546 36728 6552 36740
rect 6604 36728 6610 36780
rect 7944 36777 7972 36876
rect 10137 36839 10195 36845
rect 10137 36805 10149 36839
rect 10183 36836 10195 36839
rect 10778 36836 10784 36848
rect 10183 36808 10784 36836
rect 10183 36805 10195 36808
rect 10137 36799 10195 36805
rect 10778 36796 10784 36808
rect 10836 36796 10842 36848
rect 7929 36771 7987 36777
rect 7929 36737 7941 36771
rect 7975 36737 7987 36771
rect 7929 36731 7987 36737
rect 8036 36740 9062 36768
rect 6454 36660 6460 36712
rect 6512 36700 6518 36712
rect 8036 36700 8064 36740
rect 8386 36700 8392 36712
rect 6512 36672 8064 36700
rect 8347 36672 8392 36700
rect 6512 36660 6518 36672
rect 8386 36660 8392 36672
rect 8444 36660 8450 36712
rect 8496 36672 10364 36700
rect 8496 36632 8524 36672
rect 6380 36604 8524 36632
rect 10336 36632 10364 36672
rect 10410 36660 10416 36712
rect 10468 36700 10474 36712
rect 10870 36700 10876 36712
rect 10468 36672 10876 36700
rect 10468 36660 10474 36672
rect 10870 36660 10876 36672
rect 10928 36660 10934 36712
rect 10980 36632 11008 36876
rect 11698 36864 11704 36876
rect 11756 36864 11762 36916
rect 11790 36864 11796 36916
rect 11848 36904 11854 36916
rect 12437 36907 12495 36913
rect 12437 36904 12449 36907
rect 11848 36876 12449 36904
rect 11848 36864 11854 36876
rect 12437 36873 12449 36876
rect 12483 36904 12495 36907
rect 13814 36904 13820 36916
rect 12483 36876 13820 36904
rect 12483 36873 12495 36876
rect 12437 36867 12495 36873
rect 13814 36864 13820 36876
rect 13872 36864 13878 36916
rect 14277 36907 14335 36913
rect 14277 36873 14289 36907
rect 14323 36904 14335 36907
rect 18138 36904 18144 36916
rect 14323 36876 18144 36904
rect 14323 36873 14335 36876
rect 14277 36867 14335 36873
rect 18138 36864 18144 36876
rect 18196 36864 18202 36916
rect 35437 36907 35495 36913
rect 35437 36873 35449 36907
rect 35483 36904 35495 36907
rect 35618 36904 35624 36916
rect 35483 36876 35624 36904
rect 35483 36873 35495 36876
rect 35437 36867 35495 36873
rect 35618 36864 35624 36876
rect 35676 36864 35682 36916
rect 35802 36864 35808 36916
rect 35860 36904 35866 36916
rect 36265 36907 36323 36913
rect 36265 36904 36277 36907
rect 35860 36876 36277 36904
rect 35860 36864 35866 36876
rect 36265 36873 36277 36876
rect 36311 36873 36323 36907
rect 36265 36867 36323 36873
rect 13354 36836 13360 36848
rect 12406 36808 13360 36836
rect 11054 36728 11060 36780
rect 11112 36768 11118 36780
rect 11885 36771 11943 36777
rect 11112 36740 11157 36768
rect 11112 36728 11118 36740
rect 11885 36737 11897 36771
rect 11931 36768 11943 36771
rect 12406 36768 12434 36808
rect 13354 36796 13360 36808
rect 13412 36836 13418 36848
rect 15194 36836 15200 36848
rect 13412 36808 15200 36836
rect 13412 36796 13418 36808
rect 15194 36796 15200 36808
rect 15252 36796 15258 36848
rect 13078 36768 13084 36780
rect 11931 36740 12434 36768
rect 13039 36740 13084 36768
rect 11931 36737 11943 36740
rect 11885 36731 11943 36737
rect 13078 36728 13084 36740
rect 13136 36728 13142 36780
rect 13998 36728 14004 36780
rect 14056 36768 14062 36780
rect 14093 36771 14151 36777
rect 14093 36768 14105 36771
rect 14056 36740 14105 36768
rect 14056 36728 14062 36740
rect 14093 36737 14105 36740
rect 14139 36737 14151 36771
rect 14093 36731 14151 36737
rect 15102 36728 15108 36780
rect 15160 36768 15166 36780
rect 16853 36771 16911 36777
rect 16853 36768 16865 36771
rect 15160 36740 16865 36768
rect 15160 36728 15166 36740
rect 16853 36737 16865 36740
rect 16899 36737 16911 36771
rect 35618 36768 35624 36780
rect 35579 36740 35624 36768
rect 16853 36731 16911 36737
rect 35618 36728 35624 36740
rect 35676 36728 35682 36780
rect 36081 36771 36139 36777
rect 36081 36737 36093 36771
rect 36127 36768 36139 36771
rect 36170 36768 36176 36780
rect 36127 36740 36176 36768
rect 36127 36737 36139 36740
rect 36081 36731 36139 36737
rect 36170 36728 36176 36740
rect 36228 36728 36234 36780
rect 11974 36660 11980 36712
rect 12032 36700 12038 36712
rect 13538 36700 13544 36712
rect 12032 36672 13544 36700
rect 12032 36660 12038 36672
rect 13538 36660 13544 36672
rect 13596 36700 13602 36712
rect 14737 36703 14795 36709
rect 14737 36700 14749 36703
rect 13596 36672 14749 36700
rect 13596 36660 13602 36672
rect 14737 36669 14749 36672
rect 14783 36700 14795 36703
rect 15289 36703 15347 36709
rect 15289 36700 15301 36703
rect 14783 36672 15301 36700
rect 14783 36669 14795 36672
rect 14737 36663 14795 36669
rect 15289 36669 15301 36672
rect 15335 36700 15347 36703
rect 15841 36703 15899 36709
rect 15841 36700 15853 36703
rect 15335 36672 15853 36700
rect 15335 36669 15347 36672
rect 15289 36663 15347 36669
rect 15841 36669 15853 36672
rect 15887 36700 15899 36703
rect 16114 36700 16120 36712
rect 15887 36672 16120 36700
rect 15887 36669 15899 36672
rect 15841 36663 15899 36669
rect 16114 36660 16120 36672
rect 16172 36660 16178 36712
rect 10336 36604 10916 36632
rect 10980 36604 13032 36632
rect 3142 36524 3148 36576
rect 3200 36564 3206 36576
rect 5810 36564 5816 36576
rect 3200 36536 5816 36564
rect 3200 36524 3206 36536
rect 5810 36524 5816 36536
rect 5868 36524 5874 36576
rect 5997 36567 6055 36573
rect 5997 36533 6009 36567
rect 6043 36564 6055 36567
rect 6362 36564 6368 36576
rect 6043 36536 6368 36564
rect 6043 36533 6055 36536
rect 5997 36527 6055 36533
rect 6362 36524 6368 36536
rect 6420 36524 6426 36576
rect 7650 36524 7656 36576
rect 7708 36564 7714 36576
rect 9030 36564 9036 36576
rect 7708 36536 9036 36564
rect 7708 36524 7714 36536
rect 9030 36524 9036 36536
rect 9088 36524 9094 36576
rect 9122 36524 9128 36576
rect 9180 36564 9186 36576
rect 10410 36564 10416 36576
rect 9180 36536 10416 36564
rect 9180 36524 9186 36536
rect 10410 36524 10416 36536
rect 10468 36524 10474 36576
rect 10888 36573 10916 36604
rect 13004 36573 13032 36604
rect 14366 36592 14372 36644
rect 14424 36632 14430 36644
rect 35526 36632 35532 36644
rect 14424 36604 35532 36632
rect 14424 36592 14430 36604
rect 35526 36592 35532 36604
rect 35584 36592 35590 36644
rect 10873 36567 10931 36573
rect 10873 36533 10885 36567
rect 10919 36533 10931 36567
rect 10873 36527 10931 36533
rect 12989 36567 13047 36573
rect 12989 36533 13001 36567
rect 13035 36533 13047 36567
rect 12989 36527 13047 36533
rect 17037 36567 17095 36573
rect 17037 36533 17049 36567
rect 17083 36564 17095 36567
rect 22002 36564 22008 36576
rect 17083 36536 22008 36564
rect 17083 36533 17095 36536
rect 17037 36527 17095 36533
rect 22002 36524 22008 36536
rect 22060 36524 22066 36576
rect 1104 36474 36892 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 36892 36474
rect 1104 36400 36892 36422
rect 2222 36320 2228 36372
rect 2280 36360 2286 36372
rect 2280 36332 5120 36360
rect 2280 36320 2286 36332
rect 3329 36295 3387 36301
rect 3329 36261 3341 36295
rect 3375 36292 3387 36295
rect 4982 36292 4988 36304
rect 3375 36264 4988 36292
rect 3375 36261 3387 36264
rect 3329 36255 3387 36261
rect 4982 36252 4988 36264
rect 5040 36252 5046 36304
rect 5092 36292 5120 36332
rect 5166 36320 5172 36372
rect 5224 36360 5230 36372
rect 5224 36332 10824 36360
rect 5224 36320 5230 36332
rect 5092 36264 5212 36292
rect 1578 36224 1584 36236
rect 1539 36196 1584 36224
rect 1578 36184 1584 36196
rect 1636 36184 1642 36236
rect 1857 36227 1915 36233
rect 1857 36193 1869 36227
rect 1903 36224 1915 36227
rect 2406 36224 2412 36236
rect 1903 36196 2412 36224
rect 1903 36193 1915 36196
rect 1857 36187 1915 36193
rect 2406 36184 2412 36196
rect 2464 36184 2470 36236
rect 4525 36227 4583 36233
rect 4525 36193 4537 36227
rect 4571 36224 4583 36227
rect 5074 36224 5080 36236
rect 4571 36196 5080 36224
rect 4571 36193 4583 36196
rect 4525 36187 4583 36193
rect 5074 36184 5080 36196
rect 5132 36184 5138 36236
rect 5184 36224 5212 36264
rect 8294 36252 8300 36304
rect 8352 36292 8358 36304
rect 10796 36292 10824 36332
rect 10870 36320 10876 36372
rect 10928 36360 10934 36372
rect 11974 36360 11980 36372
rect 10928 36332 11980 36360
rect 10928 36320 10934 36332
rect 11974 36320 11980 36332
rect 12032 36320 12038 36372
rect 13633 36363 13691 36369
rect 13633 36329 13645 36363
rect 13679 36360 13691 36363
rect 13814 36360 13820 36372
rect 13679 36332 13820 36360
rect 13679 36329 13691 36332
rect 13633 36323 13691 36329
rect 13814 36320 13820 36332
rect 13872 36360 13878 36372
rect 14826 36360 14832 36372
rect 13872 36332 14832 36360
rect 13872 36320 13878 36332
rect 14826 36320 14832 36332
rect 14884 36360 14890 36372
rect 36265 36363 36323 36369
rect 14884 36332 15516 36360
rect 14884 36320 14890 36332
rect 8352 36264 9260 36292
rect 10796 36264 11100 36292
rect 8352 36252 8358 36264
rect 9122 36224 9128 36236
rect 5184 36196 8524 36224
rect 9083 36196 9128 36224
rect 5460 36168 5488 36196
rect 4801 36159 4859 36165
rect 4801 36125 4813 36159
rect 4847 36156 4859 36159
rect 5166 36156 5172 36168
rect 4847 36128 5172 36156
rect 4847 36125 4859 36128
rect 4801 36119 4859 36125
rect 5166 36116 5172 36128
rect 5224 36116 5230 36168
rect 5442 36156 5448 36168
rect 5355 36128 5448 36156
rect 5442 36116 5448 36128
rect 5500 36116 5506 36168
rect 7929 36159 7987 36165
rect 7929 36125 7941 36159
rect 7975 36156 7987 36159
rect 8294 36156 8300 36168
rect 7975 36128 8300 36156
rect 7975 36125 7987 36128
rect 7929 36119 7987 36125
rect 8294 36116 8300 36128
rect 8352 36116 8358 36168
rect 8389 36159 8447 36165
rect 8389 36125 8401 36159
rect 8435 36156 8447 36159
rect 8496 36156 8524 36196
rect 9122 36184 9128 36196
rect 9180 36184 9186 36236
rect 9232 36224 9260 36264
rect 9401 36227 9459 36233
rect 9401 36224 9413 36227
rect 9232 36196 9413 36224
rect 9401 36193 9413 36196
rect 9447 36224 9459 36227
rect 10962 36224 10968 36236
rect 9447 36196 10968 36224
rect 9447 36193 9459 36196
rect 9401 36187 9459 36193
rect 10962 36184 10968 36196
rect 11020 36184 11026 36236
rect 8662 36156 8668 36168
rect 8435 36128 8668 36156
rect 8435 36125 8447 36128
rect 8389 36119 8447 36125
rect 8662 36116 8668 36128
rect 8720 36116 8726 36168
rect 11072 36156 11100 36264
rect 12526 36252 12532 36304
rect 12584 36292 12590 36304
rect 15381 36295 15439 36301
rect 15381 36292 15393 36295
rect 12584 36264 15393 36292
rect 12584 36252 12590 36264
rect 15381 36261 15393 36264
rect 15427 36261 15439 36295
rect 15488 36292 15516 36332
rect 36265 36329 36277 36363
rect 36311 36360 36323 36363
rect 36722 36360 36728 36372
rect 36311 36332 36728 36360
rect 36311 36329 36323 36332
rect 36265 36323 36323 36329
rect 36722 36320 36728 36332
rect 36780 36320 36786 36372
rect 16577 36295 16635 36301
rect 16577 36292 16589 36295
rect 15488 36264 16589 36292
rect 15381 36255 15439 36261
rect 16577 36261 16589 36264
rect 16623 36292 16635 36295
rect 30558 36292 30564 36304
rect 16623 36264 30564 36292
rect 16623 36261 16635 36264
rect 16577 36255 16635 36261
rect 30558 36252 30564 36264
rect 30616 36252 30622 36304
rect 12526 36156 12532 36168
rect 11072 36128 12532 36156
rect 12526 36116 12532 36128
rect 12584 36116 12590 36168
rect 13081 36159 13139 36165
rect 13081 36125 13093 36159
rect 13127 36156 13139 36159
rect 15102 36156 15108 36168
rect 13127 36128 15108 36156
rect 13127 36125 13139 36128
rect 13081 36119 13139 36125
rect 15102 36116 15108 36128
rect 15160 36116 15166 36168
rect 36081 36159 36139 36165
rect 36081 36156 36093 36159
rect 35866 36128 36093 36156
rect 5353 36091 5411 36097
rect 5353 36088 5365 36091
rect 3082 36060 5365 36088
rect 5353 36057 5365 36060
rect 5399 36057 5411 36091
rect 5902 36088 5908 36100
rect 5863 36060 5908 36088
rect 5353 36051 5411 36057
rect 5902 36048 5908 36060
rect 5960 36048 5966 36100
rect 6270 36048 6276 36100
rect 6328 36088 6334 36100
rect 7650 36088 7656 36100
rect 6328 36060 6486 36088
rect 7611 36060 7656 36088
rect 6328 36048 6334 36060
rect 7650 36048 7656 36060
rect 7708 36048 7714 36100
rect 8404 36060 9812 36088
rect 4062 35980 4068 36032
rect 4120 36020 4126 36032
rect 8404 36020 8432 36060
rect 4120 35992 8432 36020
rect 8481 36023 8539 36029
rect 4120 35980 4126 35992
rect 8481 35989 8493 36023
rect 8527 36020 8539 36023
rect 9674 36020 9680 36032
rect 8527 35992 9680 36020
rect 8527 35989 8539 35992
rect 8481 35983 8539 35989
rect 9674 35980 9680 35992
rect 9732 35980 9738 36032
rect 9784 36020 9812 36060
rect 9858 36048 9864 36100
rect 9916 36048 9922 36100
rect 11054 36048 11060 36100
rect 11112 36088 11118 36100
rect 11517 36091 11575 36097
rect 11517 36088 11529 36091
rect 11112 36060 11529 36088
rect 11112 36048 11118 36060
rect 11517 36057 11529 36060
rect 11563 36088 11575 36091
rect 14366 36088 14372 36100
rect 11563 36060 14372 36088
rect 11563 36057 11575 36060
rect 11517 36051 11575 36057
rect 14366 36048 14372 36060
rect 14424 36048 14430 36100
rect 10410 36020 10416 36032
rect 9784 35992 10416 36020
rect 10410 35980 10416 35992
rect 10468 35980 10474 36032
rect 10870 36020 10876 36032
rect 10831 35992 10876 36020
rect 10870 35980 10876 35992
rect 10928 35980 10934 36032
rect 12434 35980 12440 36032
rect 12492 36020 12498 36032
rect 12989 36023 13047 36029
rect 12989 36020 13001 36023
rect 12492 35992 13001 36020
rect 12492 35980 12498 35992
rect 12989 35989 13001 35992
rect 13035 35989 13047 36023
rect 12989 35983 13047 35989
rect 13538 35980 13544 36032
rect 13596 36020 13602 36032
rect 14277 36023 14335 36029
rect 14277 36020 14289 36023
rect 13596 35992 14289 36020
rect 13596 35980 13602 35992
rect 14277 35989 14289 35992
rect 14323 35989 14335 36023
rect 15930 36020 15936 36032
rect 15891 35992 15936 36020
rect 14277 35983 14335 35989
rect 15930 35980 15936 35992
rect 15988 35980 15994 36032
rect 35342 35980 35348 36032
rect 35400 36020 35406 36032
rect 35529 36023 35587 36029
rect 35529 36020 35541 36023
rect 35400 35992 35541 36020
rect 35400 35980 35406 35992
rect 35529 35989 35541 35992
rect 35575 36020 35587 36023
rect 35866 36020 35894 36128
rect 36081 36125 36093 36128
rect 36127 36125 36139 36159
rect 36081 36119 36139 36125
rect 35575 35992 35894 36020
rect 35575 35989 35587 35992
rect 35529 35983 35587 35989
rect 1104 35930 36892 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 36892 35930
rect 1104 35856 36892 35878
rect 3326 35816 3332 35828
rect 1872 35788 3332 35816
rect 1872 35757 1900 35788
rect 3326 35776 3332 35788
rect 3384 35816 3390 35828
rect 3786 35816 3792 35828
rect 3384 35788 3792 35816
rect 3384 35776 3390 35788
rect 3786 35776 3792 35788
rect 3844 35776 3850 35828
rect 6730 35816 6736 35828
rect 4632 35788 6736 35816
rect 1857 35751 1915 35757
rect 1857 35717 1869 35751
rect 1903 35717 1915 35751
rect 4632 35748 4660 35788
rect 6730 35776 6736 35788
rect 6788 35776 6794 35828
rect 12986 35816 12992 35828
rect 6932 35788 11192 35816
rect 6178 35748 6184 35760
rect 3082 35720 4660 35748
rect 5474 35720 6184 35748
rect 1857 35711 1915 35717
rect 6178 35708 6184 35720
rect 6236 35708 6242 35760
rect 1578 35680 1584 35692
rect 1539 35652 1584 35680
rect 1578 35640 1584 35652
rect 1636 35640 1642 35692
rect 5718 35640 5724 35692
rect 5776 35680 5782 35692
rect 6932 35680 6960 35788
rect 7098 35708 7104 35760
rect 7156 35748 7162 35760
rect 7156 35720 7866 35748
rect 7156 35708 7162 35720
rect 9030 35708 9036 35760
rect 9088 35748 9094 35760
rect 9125 35751 9183 35757
rect 9125 35748 9137 35751
rect 9088 35720 9137 35748
rect 9088 35708 9094 35720
rect 9125 35717 9137 35720
rect 9171 35717 9183 35751
rect 9125 35711 9183 35717
rect 5776 35652 6960 35680
rect 5776 35640 5782 35652
rect 2590 35572 2596 35624
rect 2648 35612 2654 35624
rect 3973 35615 4031 35621
rect 3973 35612 3985 35615
rect 2648 35584 3985 35612
rect 2648 35572 2654 35584
rect 3973 35581 3985 35584
rect 4019 35581 4031 35615
rect 3973 35575 4031 35581
rect 4249 35615 4307 35621
rect 4249 35581 4261 35615
rect 4295 35612 4307 35615
rect 4706 35612 4712 35624
rect 4295 35584 4712 35612
rect 4295 35581 4307 35584
rect 4249 35575 4307 35581
rect 4706 35572 4712 35584
rect 4764 35612 4770 35624
rect 5997 35615 6055 35621
rect 4764 35584 5672 35612
rect 4764 35572 4770 35584
rect 5644 35544 5672 35584
rect 5997 35581 6009 35615
rect 6043 35612 6055 35615
rect 6362 35612 6368 35624
rect 6043 35584 6368 35612
rect 6043 35581 6055 35584
rect 5997 35575 6055 35581
rect 6362 35572 6368 35584
rect 6420 35572 6426 35624
rect 6546 35572 6552 35624
rect 6604 35612 6610 35624
rect 7101 35615 7159 35621
rect 7101 35612 7113 35615
rect 6604 35584 7113 35612
rect 6604 35572 6610 35584
rect 7101 35581 7113 35584
rect 7147 35581 7159 35615
rect 7101 35575 7159 35581
rect 7377 35615 7435 35621
rect 7377 35581 7389 35615
rect 7423 35612 7435 35615
rect 8662 35612 8668 35624
rect 7423 35584 8668 35612
rect 7423 35581 7435 35584
rect 7377 35575 7435 35581
rect 8662 35572 8668 35584
rect 8720 35572 8726 35624
rect 9140 35612 9168 35711
rect 9766 35680 9772 35692
rect 9727 35652 9772 35680
rect 9766 35640 9772 35652
rect 9824 35640 9830 35692
rect 10410 35640 10416 35692
rect 10468 35680 10474 35692
rect 10597 35683 10655 35689
rect 10597 35680 10609 35683
rect 10468 35652 10609 35680
rect 10468 35640 10474 35652
rect 10597 35649 10609 35652
rect 10643 35680 10655 35683
rect 11057 35683 11115 35689
rect 11057 35680 11069 35683
rect 10643 35652 11069 35680
rect 10643 35649 10655 35652
rect 10597 35643 10655 35649
rect 11057 35649 11069 35652
rect 11103 35649 11115 35683
rect 11057 35643 11115 35649
rect 9214 35612 9220 35624
rect 9127 35584 9220 35612
rect 9214 35572 9220 35584
rect 9272 35612 9278 35624
rect 9272 35584 10732 35612
rect 9272 35572 9278 35584
rect 10502 35544 10508 35556
rect 5644 35516 6684 35544
rect 2958 35436 2964 35488
rect 3016 35476 3022 35488
rect 3329 35479 3387 35485
rect 3329 35476 3341 35479
rect 3016 35448 3341 35476
rect 3016 35436 3022 35448
rect 3329 35445 3341 35448
rect 3375 35476 3387 35479
rect 5718 35476 5724 35488
rect 3375 35448 5724 35476
rect 3375 35445 3387 35448
rect 3329 35439 3387 35445
rect 5718 35436 5724 35448
rect 5776 35436 5782 35488
rect 6546 35476 6552 35488
rect 6507 35448 6552 35476
rect 6546 35436 6552 35448
rect 6604 35436 6610 35488
rect 6656 35476 6684 35516
rect 9646 35516 10508 35544
rect 9646 35476 9674 35516
rect 10502 35504 10508 35516
rect 10560 35504 10566 35556
rect 9950 35476 9956 35488
rect 6656 35448 9674 35476
rect 9911 35448 9956 35476
rect 9950 35436 9956 35448
rect 10008 35436 10014 35488
rect 10410 35476 10416 35488
rect 10371 35448 10416 35476
rect 10410 35436 10416 35448
rect 10468 35436 10474 35488
rect 10704 35476 10732 35584
rect 11164 35544 11192 35788
rect 12360 35788 12992 35816
rect 12360 35757 12388 35788
rect 12986 35776 12992 35788
rect 13044 35776 13050 35828
rect 13538 35816 13544 35828
rect 13499 35788 13544 35816
rect 13538 35776 13544 35788
rect 13596 35816 13602 35828
rect 14645 35819 14703 35825
rect 14645 35816 14657 35819
rect 13596 35788 14657 35816
rect 13596 35776 13602 35788
rect 14645 35785 14657 35788
rect 14691 35816 14703 35819
rect 15102 35816 15108 35828
rect 14691 35788 15108 35816
rect 14691 35785 14703 35788
rect 14645 35779 14703 35785
rect 15102 35776 15108 35788
rect 15160 35816 15166 35828
rect 15197 35819 15255 35825
rect 15197 35816 15209 35819
rect 15160 35788 15209 35816
rect 15160 35776 15166 35788
rect 15197 35785 15209 35788
rect 15243 35816 15255 35819
rect 15749 35819 15807 35825
rect 15749 35816 15761 35819
rect 15243 35788 15761 35816
rect 15243 35785 15255 35788
rect 15197 35779 15255 35785
rect 15749 35785 15761 35788
rect 15795 35816 15807 35819
rect 15930 35816 15936 35828
rect 15795 35788 15936 35816
rect 15795 35785 15807 35788
rect 15749 35779 15807 35785
rect 15930 35776 15936 35788
rect 15988 35776 15994 35828
rect 12345 35751 12403 35757
rect 12345 35717 12357 35751
rect 12391 35717 12403 35751
rect 12345 35711 12403 35717
rect 12434 35708 12440 35760
rect 12492 35748 12498 35760
rect 12492 35720 12537 35748
rect 12492 35708 12498 35720
rect 12618 35640 12624 35692
rect 12676 35680 12682 35692
rect 14093 35683 14151 35689
rect 14093 35680 14105 35683
rect 12676 35652 14105 35680
rect 12676 35640 12682 35652
rect 14093 35649 14105 35652
rect 14139 35680 14151 35683
rect 15470 35680 15476 35692
rect 14139 35652 15476 35680
rect 14139 35649 14151 35652
rect 14093 35643 14151 35649
rect 15470 35640 15476 35652
rect 15528 35640 15534 35692
rect 36081 35683 36139 35689
rect 36081 35680 36093 35683
rect 35866 35652 36093 35680
rect 11974 35612 11980 35624
rect 11935 35584 11980 35612
rect 11974 35572 11980 35584
rect 12032 35572 12038 35624
rect 15562 35612 15568 35624
rect 12406 35584 15568 35612
rect 12406 35544 12434 35584
rect 15562 35572 15568 35584
rect 15620 35572 15626 35624
rect 11164 35516 12434 35544
rect 12989 35479 13047 35485
rect 12989 35476 13001 35479
rect 10704 35448 13001 35476
rect 12989 35445 13001 35448
rect 13035 35445 13047 35479
rect 12989 35439 13047 35445
rect 35434 35436 35440 35488
rect 35492 35476 35498 35488
rect 35529 35479 35587 35485
rect 35529 35476 35541 35479
rect 35492 35448 35541 35476
rect 35492 35436 35498 35448
rect 35529 35445 35541 35448
rect 35575 35476 35587 35479
rect 35866 35476 35894 35652
rect 36081 35649 36093 35652
rect 36127 35649 36139 35683
rect 36081 35643 36139 35649
rect 36262 35476 36268 35488
rect 35575 35448 35894 35476
rect 36223 35448 36268 35476
rect 35575 35445 35587 35448
rect 35529 35439 35587 35445
rect 36262 35436 36268 35448
rect 36320 35436 36326 35488
rect 1104 35386 36892 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 36892 35386
rect 1104 35312 36892 35334
rect 1762 35232 1768 35284
rect 1820 35272 1826 35284
rect 7282 35272 7288 35284
rect 1820 35244 4016 35272
rect 1820 35232 1826 35244
rect 2590 35096 2596 35148
rect 2648 35136 2654 35148
rect 3329 35139 3387 35145
rect 3329 35136 3341 35139
rect 2648 35108 3341 35136
rect 2648 35096 2654 35108
rect 3329 35105 3341 35108
rect 3375 35105 3387 35139
rect 3329 35099 3387 35105
rect 3878 35096 3884 35148
rect 3936 35136 3942 35148
rect 3988 35136 4016 35244
rect 5552 35244 7288 35272
rect 5077 35139 5135 35145
rect 5077 35136 5089 35139
rect 3936 35108 5089 35136
rect 3936 35096 3942 35108
rect 5077 35105 5089 35108
rect 5123 35105 5135 35139
rect 5077 35099 5135 35105
rect 4433 35071 4491 35077
rect 4433 35037 4445 35071
rect 4479 35068 4491 35071
rect 4982 35068 4988 35080
rect 4479 35040 4988 35068
rect 4479 35037 4491 35040
rect 4433 35031 4491 35037
rect 4982 35028 4988 35040
rect 5040 35068 5046 35080
rect 5353 35071 5411 35077
rect 5353 35068 5365 35071
rect 5040 35040 5365 35068
rect 5040 35028 5046 35040
rect 5353 35037 5365 35040
rect 5399 35068 5411 35071
rect 5442 35068 5448 35080
rect 5399 35040 5448 35068
rect 5399 35037 5411 35040
rect 5353 35031 5411 35037
rect 5442 35028 5448 35040
rect 5500 35028 5506 35080
rect 3053 35003 3111 35009
rect 2622 34972 2774 35000
rect 1578 34932 1584 34944
rect 1539 34904 1584 34932
rect 1578 34892 1584 34904
rect 1636 34892 1642 34944
rect 2746 34932 2774 34972
rect 3053 34969 3065 35003
rect 3099 35000 3111 35003
rect 4062 35000 4068 35012
rect 3099 34972 4068 35000
rect 3099 34969 3111 34972
rect 3053 34963 3111 34969
rect 4062 34960 4068 34972
rect 4120 34960 4126 35012
rect 4157 35003 4215 35009
rect 4157 34969 4169 35003
rect 4203 35000 4215 35003
rect 4706 35000 4712 35012
rect 4203 34972 4712 35000
rect 4203 34969 4215 34972
rect 4157 34963 4215 34969
rect 4706 34960 4712 34972
rect 4764 34960 4770 35012
rect 5552 35000 5580 35244
rect 7282 35232 7288 35244
rect 7340 35232 7346 35284
rect 7374 35232 7380 35284
rect 7432 35272 7438 35284
rect 8573 35275 8631 35281
rect 7432 35244 7972 35272
rect 7432 35232 7438 35244
rect 7944 35204 7972 35244
rect 8573 35241 8585 35275
rect 8619 35272 8631 35275
rect 9766 35272 9772 35284
rect 8619 35244 9772 35272
rect 8619 35241 8631 35244
rect 8573 35235 8631 35241
rect 9766 35232 9772 35244
rect 9824 35232 9830 35284
rect 9950 35232 9956 35284
rect 10008 35272 10014 35284
rect 13081 35275 13139 35281
rect 10008 35244 12848 35272
rect 10008 35232 10014 35244
rect 12820 35204 12848 35244
rect 13081 35241 13093 35275
rect 13127 35272 13139 35275
rect 13538 35272 13544 35284
rect 13127 35244 13544 35272
rect 13127 35241 13139 35244
rect 13081 35235 13139 35241
rect 13538 35232 13544 35244
rect 13596 35272 13602 35284
rect 14277 35275 14335 35281
rect 14277 35272 14289 35275
rect 13596 35244 14289 35272
rect 13596 35232 13602 35244
rect 14277 35241 14289 35244
rect 14323 35241 14335 35275
rect 14826 35272 14832 35284
rect 14787 35244 14832 35272
rect 14277 35235 14335 35241
rect 14826 35232 14832 35244
rect 14884 35232 14890 35284
rect 28077 35275 28135 35281
rect 28077 35241 28089 35275
rect 28123 35272 28135 35275
rect 28442 35272 28448 35284
rect 28123 35244 28448 35272
rect 28123 35241 28135 35244
rect 28077 35235 28135 35241
rect 28442 35232 28448 35244
rect 28500 35232 28506 35284
rect 13998 35204 14004 35216
rect 7944 35176 9260 35204
rect 12820 35176 14004 35204
rect 6546 35096 6552 35148
rect 6604 35136 6610 35148
rect 8021 35139 8079 35145
rect 8021 35136 8033 35139
rect 6604 35108 8033 35136
rect 6604 35096 6610 35108
rect 8021 35105 8033 35108
rect 8067 35136 8079 35139
rect 8294 35136 8300 35148
rect 8067 35108 8300 35136
rect 8067 35105 8079 35108
rect 8021 35099 8079 35105
rect 8294 35096 8300 35108
rect 8352 35136 8358 35148
rect 8754 35136 8760 35148
rect 8352 35108 8760 35136
rect 8352 35096 8358 35108
rect 8754 35096 8760 35108
rect 8812 35136 8818 35148
rect 9122 35136 9128 35148
rect 8812 35108 9128 35136
rect 8812 35096 8818 35108
rect 9122 35096 9128 35108
rect 9180 35096 9186 35148
rect 9232 35136 9260 35176
rect 13998 35164 14004 35176
rect 14056 35164 14062 35216
rect 10686 35136 10692 35148
rect 9232 35108 10692 35136
rect 10686 35096 10692 35108
rect 10744 35096 10750 35148
rect 11517 35139 11575 35145
rect 11517 35105 11529 35139
rect 11563 35136 11575 35139
rect 11698 35136 11704 35148
rect 11563 35108 11704 35136
rect 11563 35105 11575 35108
rect 11517 35099 11575 35105
rect 11698 35096 11704 35108
rect 11756 35096 11762 35148
rect 11790 35096 11796 35148
rect 11848 35136 11854 35148
rect 11848 35108 11893 35136
rect 11848 35096 11854 35108
rect 12894 35096 12900 35148
rect 12952 35136 12958 35148
rect 13170 35136 13176 35148
rect 12952 35108 13176 35136
rect 12952 35096 12958 35108
rect 13170 35096 13176 35108
rect 13228 35096 13234 35148
rect 15562 35068 15568 35080
rect 15523 35040 15568 35068
rect 15562 35028 15568 35040
rect 15620 35028 15626 35080
rect 27890 35068 27896 35080
rect 27803 35040 27896 35068
rect 27890 35028 27896 35040
rect 27948 35068 27954 35080
rect 28629 35071 28687 35077
rect 28629 35068 28641 35071
rect 27948 35040 28641 35068
rect 27948 35028 27954 35040
rect 28629 35037 28641 35040
rect 28675 35068 28687 35071
rect 35894 35068 35900 35080
rect 28675 35040 35900 35068
rect 28675 35037 28687 35040
rect 28629 35031 28687 35037
rect 35894 35028 35900 35040
rect 35952 35028 35958 35080
rect 5092 34972 5580 35000
rect 5092 34932 5120 34972
rect 5626 34960 5632 35012
rect 5684 35000 5690 35012
rect 5997 35003 6055 35009
rect 5997 35000 6009 35003
rect 5684 34972 6009 35000
rect 5684 34960 5690 34972
rect 5997 34969 6009 34972
rect 6043 34969 6055 35003
rect 7466 35000 7472 35012
rect 7314 34972 7472 35000
rect 5997 34963 6055 34969
rect 7466 34960 7472 34972
rect 7524 34960 7530 35012
rect 7745 35003 7803 35009
rect 7745 34969 7757 35003
rect 7791 34969 7803 35003
rect 7745 34963 7803 34969
rect 2746 34904 5120 34932
rect 6178 34892 6184 34944
rect 6236 34932 6242 34944
rect 7006 34932 7012 34944
rect 6236 34904 7012 34932
rect 6236 34892 6242 34904
rect 7006 34892 7012 34904
rect 7064 34892 7070 34944
rect 7760 34932 7788 34963
rect 8478 34960 8484 35012
rect 8536 35000 8542 35012
rect 9030 35000 9036 35012
rect 8536 34972 9036 35000
rect 8536 34960 8542 34972
rect 9030 34960 9036 34972
rect 9088 35000 9094 35012
rect 9401 35003 9459 35009
rect 9401 35000 9413 35003
rect 9088 34972 9413 35000
rect 9088 34960 9094 34972
rect 9401 34969 9413 34972
rect 9447 34969 9459 35003
rect 9401 34963 9459 34969
rect 9674 34960 9680 35012
rect 9732 35000 9738 35012
rect 9732 34972 9890 35000
rect 10704 34972 11008 35000
rect 9732 34960 9738 34972
rect 8386 34932 8392 34944
rect 7760 34904 8392 34932
rect 8386 34892 8392 34904
rect 8444 34932 8450 34944
rect 10704 34932 10732 34972
rect 8444 34904 10732 34932
rect 8444 34892 8450 34904
rect 10778 34892 10784 34944
rect 10836 34932 10842 34944
rect 10873 34935 10931 34941
rect 10873 34932 10885 34935
rect 10836 34904 10885 34932
rect 10836 34892 10842 34904
rect 10873 34901 10885 34904
rect 10919 34901 10931 34935
rect 10980 34932 11008 34972
rect 11606 34960 11612 35012
rect 11664 35000 11670 35012
rect 11664 34972 11709 35000
rect 11664 34960 11670 34972
rect 12526 34932 12532 34944
rect 10980 34904 12532 34932
rect 10873 34895 10931 34901
rect 12526 34892 12532 34904
rect 12584 34932 12590 34944
rect 13541 34935 13599 34941
rect 13541 34932 13553 34935
rect 12584 34904 13553 34932
rect 12584 34892 12590 34904
rect 13541 34901 13553 34904
rect 13587 34901 13599 34935
rect 15654 34932 15660 34944
rect 15615 34904 15660 34932
rect 13541 34895 13599 34901
rect 15654 34892 15660 34904
rect 15712 34892 15718 34944
rect 16393 34935 16451 34941
rect 16393 34901 16405 34935
rect 16439 34932 16451 34935
rect 16942 34932 16948 34944
rect 16439 34904 16948 34932
rect 16439 34901 16451 34904
rect 16393 34895 16451 34901
rect 16942 34892 16948 34904
rect 17000 34892 17006 34944
rect 1104 34842 36892 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 36892 34842
rect 1104 34768 36892 34790
rect 2225 34731 2283 34737
rect 2225 34697 2237 34731
rect 2271 34728 2283 34731
rect 2406 34728 2412 34740
rect 2271 34700 2412 34728
rect 2271 34697 2283 34700
rect 2225 34691 2283 34697
rect 2406 34688 2412 34700
rect 2464 34688 2470 34740
rect 2682 34688 2688 34740
rect 2740 34728 2746 34740
rect 2740 34700 4016 34728
rect 2740 34688 2746 34700
rect 3234 34620 3240 34672
rect 3292 34620 3298 34672
rect 3694 34660 3700 34672
rect 3655 34632 3700 34660
rect 3694 34620 3700 34632
rect 3752 34620 3758 34672
rect 3988 34604 4016 34700
rect 5718 34688 5724 34740
rect 5776 34728 5782 34740
rect 6641 34731 6699 34737
rect 6641 34728 6653 34731
rect 5776 34700 6653 34728
rect 5776 34688 5782 34700
rect 6641 34697 6653 34700
rect 6687 34697 6699 34731
rect 6641 34691 6699 34697
rect 6822 34688 6828 34740
rect 6880 34728 6886 34740
rect 7285 34731 7343 34737
rect 7285 34728 7297 34731
rect 6880 34700 7297 34728
rect 6880 34688 6886 34700
rect 7285 34697 7297 34700
rect 7331 34697 7343 34731
rect 9858 34728 9864 34740
rect 7285 34691 7343 34697
rect 7392 34700 9864 34728
rect 5166 34660 5172 34672
rect 4816 34632 5172 34660
rect 1762 34592 1768 34604
rect 1723 34564 1768 34592
rect 1762 34552 1768 34564
rect 1820 34552 1826 34604
rect 3970 34552 3976 34604
rect 4028 34592 4034 34604
rect 4816 34592 4844 34632
rect 5166 34620 5172 34632
rect 5224 34620 5230 34672
rect 5350 34620 5356 34672
rect 5408 34660 5414 34672
rect 7392 34660 7420 34700
rect 9858 34688 9864 34700
rect 9916 34688 9922 34740
rect 9950 34688 9956 34740
rect 10008 34728 10014 34740
rect 14001 34731 14059 34737
rect 14001 34728 14013 34731
rect 10008 34700 14013 34728
rect 10008 34688 10014 34700
rect 14001 34697 14013 34700
rect 14047 34697 14059 34731
rect 14001 34691 14059 34697
rect 14645 34731 14703 34737
rect 14645 34697 14657 34731
rect 14691 34728 14703 34731
rect 14826 34728 14832 34740
rect 14691 34700 14832 34728
rect 14691 34697 14703 34700
rect 14645 34691 14703 34697
rect 14826 34688 14832 34700
rect 14884 34688 14890 34740
rect 15102 34728 15108 34740
rect 15063 34700 15108 34728
rect 15102 34688 15108 34700
rect 15160 34688 15166 34740
rect 5408 34632 7420 34660
rect 5408 34620 5414 34632
rect 8478 34620 8484 34672
rect 8536 34660 8542 34672
rect 8536 34632 8602 34660
rect 8536 34620 8542 34632
rect 9490 34620 9496 34672
rect 9548 34660 9554 34672
rect 10134 34660 10140 34672
rect 9548 34632 10140 34660
rect 9548 34620 9554 34632
rect 10134 34620 10140 34632
rect 10192 34660 10198 34672
rect 10594 34660 10600 34672
rect 10192 34632 10600 34660
rect 10192 34620 10198 34632
rect 10594 34620 10600 34632
rect 10652 34620 10658 34672
rect 11790 34660 11796 34672
rect 11751 34632 11796 34660
rect 11790 34620 11796 34632
rect 11848 34620 11854 34672
rect 12713 34663 12771 34669
rect 12713 34629 12725 34663
rect 12759 34660 12771 34663
rect 13449 34663 13507 34669
rect 13449 34660 13461 34663
rect 12759 34632 13461 34660
rect 12759 34629 12771 34632
rect 12713 34623 12771 34629
rect 13449 34629 13461 34632
rect 13495 34629 13507 34663
rect 13449 34623 13507 34629
rect 15654 34620 15660 34672
rect 15712 34660 15718 34672
rect 17037 34663 17095 34669
rect 17037 34660 17049 34663
rect 15712 34632 17049 34660
rect 15712 34620 15718 34632
rect 17037 34629 17049 34632
rect 17083 34629 17095 34663
rect 17037 34623 17095 34629
rect 4028 34564 4121 34592
rect 4632 34564 4844 34592
rect 4893 34595 4951 34601
rect 4028 34552 4034 34564
rect 1673 34527 1731 34533
rect 1673 34493 1685 34527
rect 1719 34524 1731 34527
rect 4632 34524 4660 34564
rect 4893 34561 4905 34595
rect 4939 34592 4951 34595
rect 4982 34592 4988 34604
rect 4939 34564 4988 34592
rect 4939 34561 4951 34564
rect 4893 34555 4951 34561
rect 4982 34552 4988 34564
rect 5040 34552 5046 34604
rect 5534 34592 5540 34604
rect 5495 34564 5540 34592
rect 5534 34552 5540 34564
rect 5592 34552 5598 34604
rect 6733 34595 6791 34601
rect 6733 34561 6745 34595
rect 6779 34592 6791 34595
rect 6822 34592 6828 34604
rect 6779 34564 6828 34592
rect 6779 34561 6791 34564
rect 6733 34555 6791 34561
rect 6822 34552 6828 34564
rect 6880 34592 6886 34604
rect 7377 34595 7435 34601
rect 7377 34592 7389 34595
rect 6880 34564 7389 34592
rect 6880 34552 6886 34564
rect 7377 34561 7389 34564
rect 7423 34561 7435 34595
rect 10962 34592 10968 34604
rect 10923 34564 10968 34592
rect 7377 34555 7435 34561
rect 10962 34552 10968 34564
rect 11020 34552 11026 34604
rect 13262 34552 13268 34604
rect 13320 34592 13326 34604
rect 13357 34595 13415 34601
rect 13357 34592 13369 34595
rect 13320 34564 13369 34592
rect 13320 34552 13326 34564
rect 13357 34561 13369 34564
rect 13403 34561 13415 34595
rect 13357 34555 13415 34561
rect 1719 34496 4660 34524
rect 4709 34527 4767 34533
rect 1719 34493 1731 34496
rect 1673 34487 1731 34493
rect 4709 34493 4721 34527
rect 4755 34493 4767 34527
rect 5350 34524 5356 34536
rect 5311 34496 5356 34524
rect 4709 34487 4767 34493
rect 4724 34456 4752 34487
rect 5350 34484 5356 34496
rect 5408 34484 5414 34536
rect 8297 34527 8355 34533
rect 8297 34493 8309 34527
rect 8343 34524 8355 34527
rect 9398 34524 9404 34536
rect 8343 34496 9404 34524
rect 8343 34493 8355 34496
rect 8297 34487 8355 34493
rect 9398 34484 9404 34496
rect 9456 34484 9462 34536
rect 9766 34524 9772 34536
rect 9727 34496 9772 34524
rect 9766 34484 9772 34496
rect 9824 34484 9830 34536
rect 10045 34527 10103 34533
rect 10045 34493 10057 34527
rect 10091 34493 10103 34527
rect 10045 34487 10103 34493
rect 5534 34456 5540 34468
rect 4724 34428 5540 34456
rect 5534 34416 5540 34428
rect 5592 34416 5598 34468
rect 5902 34416 5908 34468
rect 5960 34456 5966 34468
rect 6638 34456 6644 34468
rect 5960 34428 6644 34456
rect 5960 34416 5966 34428
rect 6638 34416 6644 34428
rect 6696 34416 6702 34468
rect 9582 34348 9588 34400
rect 9640 34388 9646 34400
rect 10060 34388 10088 34487
rect 11974 34484 11980 34536
rect 12032 34524 12038 34536
rect 12805 34527 12863 34533
rect 12805 34524 12817 34527
rect 12032 34496 12817 34524
rect 12032 34484 12038 34496
rect 12805 34493 12817 34496
rect 12851 34493 12863 34527
rect 12805 34487 12863 34493
rect 13170 34484 13176 34536
rect 13228 34524 13234 34536
rect 16942 34524 16948 34536
rect 13228 34496 16804 34524
rect 16903 34496 16948 34524
rect 13228 34484 13234 34496
rect 11790 34416 11796 34468
rect 11848 34456 11854 34468
rect 12342 34456 12348 34468
rect 11848 34428 12348 34456
rect 11848 34416 11854 34428
rect 12342 34416 12348 34428
rect 12400 34456 12406 34468
rect 16776 34456 16804 34496
rect 16942 34484 16948 34496
rect 17000 34484 17006 34536
rect 17221 34527 17279 34533
rect 17221 34524 17233 34527
rect 17052 34496 17233 34524
rect 17052 34456 17080 34496
rect 17221 34493 17233 34496
rect 17267 34493 17279 34527
rect 17221 34487 17279 34493
rect 12400 34428 16574 34456
rect 16776 34428 17080 34456
rect 12400 34416 12406 34428
rect 9640 34360 10088 34388
rect 11057 34391 11115 34397
rect 9640 34348 9646 34360
rect 11057 34357 11069 34391
rect 11103 34388 11115 34391
rect 11514 34388 11520 34400
rect 11103 34360 11520 34388
rect 11103 34357 11115 34360
rect 11057 34351 11115 34357
rect 11514 34348 11520 34360
rect 11572 34348 11578 34400
rect 16546 34388 16574 34428
rect 34790 34388 34796 34400
rect 16546 34360 34796 34388
rect 34790 34348 34796 34360
rect 34848 34348 34854 34400
rect 1104 34298 36892 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 36892 34298
rect 1104 34224 36892 34246
rect 3970 34184 3976 34196
rect 3931 34156 3976 34184
rect 3970 34144 3976 34156
rect 4028 34144 4034 34196
rect 5810 34144 5816 34196
rect 5868 34184 5874 34196
rect 7101 34187 7159 34193
rect 7101 34184 7113 34187
rect 5868 34156 7113 34184
rect 5868 34144 5874 34156
rect 7101 34153 7113 34156
rect 7147 34153 7159 34187
rect 7101 34147 7159 34153
rect 7745 34187 7803 34193
rect 7745 34153 7757 34187
rect 7791 34184 7803 34187
rect 7834 34184 7840 34196
rect 7791 34156 7840 34184
rect 7791 34153 7803 34156
rect 7745 34147 7803 34153
rect 7834 34144 7840 34156
rect 7892 34144 7898 34196
rect 12986 34184 12992 34196
rect 7944 34156 12434 34184
rect 12947 34156 12992 34184
rect 3421 34051 3479 34057
rect 3421 34017 3433 34051
rect 3467 34048 3479 34051
rect 3988 34048 4016 34144
rect 6638 34076 6644 34128
rect 6696 34116 6702 34128
rect 7944 34116 7972 34156
rect 6696 34088 7972 34116
rect 6696 34076 6702 34088
rect 8754 34076 8760 34128
rect 8812 34116 8818 34128
rect 9125 34119 9183 34125
rect 9125 34116 9137 34119
rect 8812 34088 9137 34116
rect 8812 34076 8818 34088
rect 9125 34085 9137 34088
rect 9171 34116 9183 34119
rect 9582 34116 9588 34128
rect 9171 34088 9588 34116
rect 9171 34085 9183 34088
rect 9125 34079 9183 34085
rect 9582 34076 9588 34088
rect 9640 34116 9646 34128
rect 12406 34116 12434 34156
rect 12986 34144 12992 34156
rect 13044 34144 13050 34196
rect 14366 34184 14372 34196
rect 14327 34156 14372 34184
rect 14366 34144 14372 34156
rect 14424 34144 14430 34196
rect 14921 34187 14979 34193
rect 14921 34153 14933 34187
rect 14967 34184 14979 34187
rect 15102 34184 15108 34196
rect 14967 34156 15108 34184
rect 14967 34153 14979 34156
rect 14921 34147 14979 34153
rect 15102 34144 15108 34156
rect 15160 34184 15166 34196
rect 15381 34187 15439 34193
rect 15381 34184 15393 34187
rect 15160 34156 15393 34184
rect 15160 34144 15166 34156
rect 15381 34153 15393 34156
rect 15427 34153 15439 34187
rect 15381 34147 15439 34153
rect 14458 34116 14464 34128
rect 9640 34088 9720 34116
rect 12406 34088 14464 34116
rect 9640 34076 9646 34088
rect 5902 34048 5908 34060
rect 3467 34020 4016 34048
rect 5092 34020 5908 34048
rect 3467 34017 3479 34020
rect 3421 34011 3479 34017
rect 5092 33980 5120 34020
rect 5902 34008 5908 34020
rect 5960 34008 5966 34060
rect 6178 34008 6184 34060
rect 6236 34048 6242 34060
rect 6546 34048 6552 34060
rect 6236 34020 6552 34048
rect 6236 34008 6242 34020
rect 6546 34008 6552 34020
rect 6604 34008 6610 34060
rect 6730 34008 6736 34060
rect 6788 34048 6794 34060
rect 8389 34051 8447 34057
rect 8389 34048 8401 34051
rect 6788 34020 8401 34048
rect 6788 34008 6794 34020
rect 8389 34017 8401 34020
rect 8435 34017 8447 34051
rect 8389 34011 8447 34017
rect 7190 33980 7196 33992
rect 4448 33952 5120 33980
rect 7151 33952 7196 33980
rect 3145 33915 3203 33921
rect 2714 33884 2774 33912
rect 1673 33847 1731 33853
rect 1673 33813 1685 33847
rect 1719 33844 1731 33847
rect 2222 33844 2228 33856
rect 1719 33816 2228 33844
rect 1719 33813 1731 33816
rect 1673 33807 1731 33813
rect 2222 33804 2228 33816
rect 2280 33804 2286 33856
rect 2746 33844 2774 33884
rect 3145 33881 3157 33915
rect 3191 33912 3203 33915
rect 4448 33912 4476 33952
rect 7190 33940 7196 33952
rect 7248 33940 7254 33992
rect 7374 33940 7380 33992
rect 7432 33980 7438 33992
rect 9692 33989 9720 34088
rect 14458 34076 14464 34088
rect 14516 34116 14522 34128
rect 15933 34119 15991 34125
rect 15933 34116 15945 34119
rect 14516 34088 15945 34116
rect 14516 34076 14522 34088
rect 15933 34085 15945 34088
rect 15979 34085 15991 34119
rect 15933 34079 15991 34085
rect 9766 34008 9772 34060
rect 9824 34048 9830 34060
rect 9824 34020 12940 34048
rect 9824 34008 9830 34020
rect 7837 33983 7895 33989
rect 7837 33980 7849 33983
rect 7432 33952 7849 33980
rect 7432 33940 7438 33952
rect 7837 33949 7849 33952
rect 7883 33949 7895 33983
rect 8297 33983 8355 33989
rect 8297 33980 8309 33983
rect 7837 33943 7895 33949
rect 8036 33952 8309 33980
rect 3191 33884 4476 33912
rect 4525 33915 4583 33921
rect 3191 33881 3203 33884
rect 3145 33875 3203 33881
rect 4525 33881 4537 33915
rect 4571 33912 4583 33915
rect 4798 33912 4804 33924
rect 4571 33884 4804 33912
rect 4571 33881 4583 33884
rect 4525 33875 4583 33881
rect 4798 33872 4804 33884
rect 4856 33872 4862 33924
rect 6273 33915 6331 33921
rect 5842 33884 6224 33912
rect 5902 33844 5908 33856
rect 2746 33816 5908 33844
rect 5902 33804 5908 33816
rect 5960 33804 5966 33856
rect 6196 33844 6224 33884
rect 6273 33881 6285 33915
rect 6319 33912 6331 33915
rect 6362 33912 6368 33924
rect 6319 33884 6368 33912
rect 6319 33881 6331 33884
rect 6273 33875 6331 33881
rect 6362 33872 6368 33884
rect 6420 33872 6426 33924
rect 7926 33912 7932 33924
rect 6472 33884 7932 33912
rect 6472 33844 6500 33884
rect 7926 33872 7932 33884
rect 7984 33872 7990 33924
rect 6196 33816 6500 33844
rect 7190 33804 7196 33856
rect 7248 33844 7254 33856
rect 8036 33844 8064 33952
rect 8297 33949 8309 33952
rect 8343 33949 8355 33983
rect 8297 33943 8355 33949
rect 9677 33983 9735 33989
rect 9677 33949 9689 33983
rect 9723 33980 9735 33983
rect 10229 33983 10287 33989
rect 10229 33980 10241 33983
rect 9723 33952 10241 33980
rect 9723 33949 9735 33952
rect 9677 33943 9735 33949
rect 10229 33949 10241 33952
rect 10275 33949 10287 33983
rect 10229 33943 10287 33949
rect 10778 33940 10784 33992
rect 10836 33940 10842 33992
rect 12912 33989 12940 34020
rect 12897 33983 12955 33989
rect 12897 33949 12909 33983
rect 12943 33949 12955 33983
rect 12897 33943 12955 33949
rect 13725 33983 13783 33989
rect 13725 33949 13737 33983
rect 13771 33980 13783 33983
rect 14366 33980 14372 33992
rect 13771 33952 14372 33980
rect 13771 33949 13783 33952
rect 13725 33943 13783 33949
rect 14366 33940 14372 33952
rect 14424 33940 14430 33992
rect 34790 33940 34796 33992
rect 34848 33980 34854 33992
rect 34885 33983 34943 33989
rect 34885 33980 34897 33983
rect 34848 33952 34897 33980
rect 34848 33940 34854 33952
rect 34885 33949 34897 33952
rect 34931 33980 34943 33983
rect 35529 33983 35587 33989
rect 35529 33980 35541 33983
rect 34931 33952 35541 33980
rect 34931 33949 34943 33952
rect 34885 33943 34943 33949
rect 35529 33949 35541 33952
rect 35575 33949 35587 33983
rect 35529 33943 35587 33949
rect 8202 33872 8208 33924
rect 8260 33912 8266 33924
rect 10796 33912 10824 33940
rect 11422 33912 11428 33924
rect 8260 33884 10824 33912
rect 11383 33884 11428 33912
rect 8260 33872 8266 33884
rect 11422 33872 11428 33884
rect 11480 33872 11486 33924
rect 11514 33872 11520 33924
rect 11572 33912 11578 33924
rect 11572 33884 11617 33912
rect 11572 33872 11578 33884
rect 12342 33872 12348 33924
rect 12400 33912 12406 33924
rect 12437 33915 12495 33921
rect 12437 33912 12449 33915
rect 12400 33884 12449 33912
rect 12400 33872 12406 33884
rect 12437 33881 12449 33884
rect 12483 33881 12495 33915
rect 12437 33875 12495 33881
rect 7248 33816 8064 33844
rect 7248 33804 7254 33816
rect 8662 33804 8668 33856
rect 8720 33844 8726 33856
rect 10781 33847 10839 33853
rect 10781 33844 10793 33847
rect 8720 33816 10793 33844
rect 8720 33804 8726 33816
rect 10781 33813 10793 33816
rect 10827 33813 10839 33847
rect 10781 33807 10839 33813
rect 10962 33804 10968 33856
rect 11020 33844 11026 33856
rect 13262 33844 13268 33856
rect 11020 33816 13268 33844
rect 11020 33804 11026 33816
rect 13262 33804 13268 33816
rect 13320 33804 13326 33856
rect 13630 33844 13636 33856
rect 13591 33816 13636 33844
rect 13630 33804 13636 33816
rect 13688 33804 13694 33856
rect 34974 33844 34980 33856
rect 34935 33816 34980 33844
rect 34974 33804 34980 33816
rect 35032 33804 35038 33856
rect 1104 33754 36892 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 36892 33754
rect 1104 33680 36892 33702
rect 2222 33600 2228 33652
rect 2280 33640 2286 33652
rect 4982 33640 4988 33652
rect 2280 33612 4988 33640
rect 2280 33600 2286 33612
rect 4982 33600 4988 33612
rect 5040 33600 5046 33652
rect 6641 33643 6699 33649
rect 6641 33609 6653 33643
rect 6687 33640 6699 33643
rect 7098 33640 7104 33652
rect 6687 33612 7104 33640
rect 6687 33609 6699 33612
rect 6641 33603 6699 33609
rect 7098 33600 7104 33612
rect 7156 33600 7162 33652
rect 7282 33640 7288 33652
rect 7243 33612 7288 33640
rect 7282 33600 7288 33612
rect 7340 33600 7346 33652
rect 9306 33600 9312 33652
rect 9364 33640 9370 33652
rect 9364 33612 10548 33640
rect 9364 33600 9370 33612
rect 2498 33572 2504 33584
rect 1964 33544 2504 33572
rect 1670 33464 1676 33516
rect 1728 33504 1734 33516
rect 1964 33513 1992 33544
rect 2498 33532 2504 33544
rect 2556 33532 2562 33584
rect 3602 33572 3608 33584
rect 3450 33544 3608 33572
rect 3602 33532 3608 33544
rect 3660 33532 3666 33584
rect 5442 33572 5448 33584
rect 5290 33544 5448 33572
rect 5442 33532 5448 33544
rect 5500 33532 5506 33584
rect 5721 33575 5779 33581
rect 5721 33541 5733 33575
rect 5767 33572 5779 33575
rect 8202 33572 8208 33584
rect 5767 33544 8208 33572
rect 5767 33541 5779 33544
rect 5721 33535 5779 33541
rect 8202 33532 8208 33544
rect 8260 33532 8266 33584
rect 8386 33532 8392 33584
rect 8444 33572 8450 33584
rect 10045 33575 10103 33581
rect 8444 33544 8878 33572
rect 8444 33532 8450 33544
rect 10045 33541 10057 33575
rect 10091 33572 10103 33575
rect 10410 33572 10416 33584
rect 10091 33544 10416 33572
rect 10091 33541 10103 33544
rect 10045 33535 10103 33541
rect 10410 33532 10416 33544
rect 10468 33532 10474 33584
rect 1949 33507 2007 33513
rect 1949 33504 1961 33507
rect 1728 33476 1961 33504
rect 1728 33464 1734 33476
rect 1949 33473 1961 33476
rect 1995 33473 2007 33507
rect 6546 33504 6552 33516
rect 6507 33476 6552 33504
rect 1949 33467 2007 33473
rect 6546 33464 6552 33476
rect 6604 33504 6610 33516
rect 6822 33504 6828 33516
rect 6604 33476 6828 33504
rect 6604 33464 6610 33476
rect 6822 33464 6828 33476
rect 6880 33464 6886 33516
rect 7190 33464 7196 33516
rect 7248 33504 7254 33516
rect 7377 33507 7435 33513
rect 7377 33504 7389 33507
rect 7248 33476 7389 33504
rect 7248 33464 7254 33476
rect 7377 33473 7389 33476
rect 7423 33473 7435 33507
rect 10520 33504 10548 33612
rect 11606 33600 11612 33652
rect 11664 33640 11670 33652
rect 11977 33643 12035 33649
rect 11977 33640 11989 33643
rect 11664 33612 11989 33640
rect 11664 33600 11670 33612
rect 11977 33609 11989 33612
rect 12023 33609 12035 33643
rect 11977 33603 12035 33609
rect 14829 33643 14887 33649
rect 14829 33609 14841 33643
rect 14875 33640 14887 33643
rect 15102 33640 15108 33652
rect 14875 33612 15108 33640
rect 14875 33609 14887 33612
rect 14829 33603 14887 33609
rect 15102 33600 15108 33612
rect 15160 33640 15166 33652
rect 15289 33643 15347 33649
rect 15289 33640 15301 33643
rect 15160 33612 15301 33640
rect 15160 33600 15166 33612
rect 15289 33609 15301 33612
rect 15335 33609 15347 33643
rect 31478 33640 31484 33652
rect 31439 33612 31484 33640
rect 15289 33603 15347 33609
rect 31478 33600 31484 33612
rect 31536 33600 31542 33652
rect 10778 33532 10784 33584
rect 10836 33572 10842 33584
rect 12250 33572 12256 33584
rect 10836 33544 12256 33572
rect 10836 33532 10842 33544
rect 12250 33532 12256 33544
rect 12308 33572 12314 33584
rect 12529 33575 12587 33581
rect 12529 33572 12541 33575
rect 12308 33544 12541 33572
rect 12308 33532 12314 33544
rect 12529 33541 12541 33544
rect 12575 33541 12587 33575
rect 12529 33535 12587 33541
rect 11885 33507 11943 33513
rect 11885 33504 11897 33507
rect 10520 33476 11897 33504
rect 7377 33467 7435 33473
rect 11885 33473 11897 33476
rect 11931 33473 11943 33507
rect 13262 33504 13268 33516
rect 13223 33476 13268 33504
rect 11885 33467 11943 33473
rect 13262 33464 13268 33476
rect 13320 33464 13326 33516
rect 13998 33464 14004 33516
rect 14056 33504 14062 33516
rect 14093 33507 14151 33513
rect 14093 33504 14105 33507
rect 14056 33476 14105 33504
rect 14056 33464 14062 33476
rect 14093 33473 14105 33476
rect 14139 33473 14151 33507
rect 14093 33467 14151 33473
rect 31297 33507 31355 33513
rect 31297 33473 31309 33507
rect 31343 33473 31355 33507
rect 31297 33467 31355 33473
rect 2222 33436 2228 33448
rect 2183 33408 2228 33436
rect 2222 33396 2228 33408
rect 2280 33396 2286 33448
rect 3694 33436 3700 33448
rect 3607 33408 3700 33436
rect 3694 33396 3700 33408
rect 3752 33436 3758 33448
rect 5997 33439 6055 33445
rect 3752 33408 5948 33436
rect 3752 33396 3758 33408
rect 5920 33368 5948 33408
rect 5997 33405 6009 33439
rect 6043 33436 6055 33439
rect 6086 33436 6092 33448
rect 6043 33408 6092 33436
rect 6043 33405 6055 33408
rect 5997 33399 6055 33405
rect 6086 33396 6092 33408
rect 6144 33396 6150 33448
rect 6840 33436 6868 33464
rect 7282 33436 7288 33448
rect 6840 33408 7288 33436
rect 7282 33396 7288 33408
rect 7340 33396 7346 33448
rect 8297 33439 8355 33445
rect 8297 33405 8309 33439
rect 8343 33436 8355 33439
rect 8846 33436 8852 33448
rect 8343 33408 8852 33436
rect 8343 33405 8355 33408
rect 8297 33399 8355 33405
rect 8846 33396 8852 33408
rect 8904 33396 8910 33448
rect 9582 33396 9588 33448
rect 9640 33436 9646 33448
rect 10321 33439 10379 33445
rect 10321 33436 10333 33439
rect 9640 33408 10333 33436
rect 9640 33396 9646 33408
rect 10321 33405 10333 33408
rect 10367 33436 10379 33439
rect 10781 33439 10839 33445
rect 10781 33436 10793 33439
rect 10367 33408 10793 33436
rect 10367 33405 10379 33408
rect 10321 33399 10379 33405
rect 10781 33405 10793 33408
rect 10827 33405 10839 33439
rect 31312 33436 31340 33467
rect 34974 33464 34980 33516
rect 35032 33504 35038 33516
rect 36081 33507 36139 33513
rect 36081 33504 36093 33507
rect 35032 33476 36093 33504
rect 35032 33464 35038 33476
rect 36081 33473 36093 33476
rect 36127 33473 36139 33507
rect 36081 33467 36139 33473
rect 36446 33436 36452 33448
rect 31312 33408 36452 33436
rect 10781 33399 10839 33405
rect 36446 33396 36452 33408
rect 36504 33396 36510 33448
rect 7834 33368 7840 33380
rect 5920 33340 7840 33368
rect 7834 33328 7840 33340
rect 7892 33328 7898 33380
rect 36262 33368 36268 33380
rect 36223 33340 36268 33368
rect 36262 33328 36268 33340
rect 36320 33328 36326 33380
rect 4154 33260 4160 33312
rect 4212 33300 4218 33312
rect 4249 33303 4307 33309
rect 4249 33300 4261 33303
rect 4212 33272 4261 33300
rect 4212 33260 4218 33272
rect 4249 33269 4261 33272
rect 4295 33300 4307 33303
rect 10962 33300 10968 33312
rect 4295 33272 10968 33300
rect 4295 33269 4307 33272
rect 4249 33263 4307 33269
rect 10962 33260 10968 33272
rect 11020 33260 11026 33312
rect 13357 33303 13415 33309
rect 13357 33269 13369 33303
rect 13403 33300 13415 33303
rect 13538 33300 13544 33312
rect 13403 33272 13544 33300
rect 13403 33269 13415 33272
rect 13357 33263 13415 33269
rect 13538 33260 13544 33272
rect 13596 33260 13602 33312
rect 14185 33303 14243 33309
rect 14185 33269 14197 33303
rect 14231 33300 14243 33303
rect 14366 33300 14372 33312
rect 14231 33272 14372 33300
rect 14231 33269 14243 33272
rect 14185 33263 14243 33269
rect 14366 33260 14372 33272
rect 14424 33260 14430 33312
rect 1104 33210 36892 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 36892 33210
rect 1104 33136 36892 33158
rect 1578 33056 1584 33108
rect 1636 33096 1642 33108
rect 5442 33096 5448 33108
rect 1636 33068 4936 33096
rect 5403 33068 5448 33096
rect 1636 33056 1642 33068
rect 4798 33028 4804 33040
rect 3344 33000 4804 33028
rect 1670 32960 1676 32972
rect 1631 32932 1676 32960
rect 1670 32920 1676 32932
rect 1728 32920 1734 32972
rect 1949 32963 2007 32969
rect 1949 32929 1961 32963
rect 1995 32960 2007 32963
rect 3344 32960 3372 33000
rect 4798 32988 4804 33000
rect 4856 32988 4862 33040
rect 4908 33028 4936 33068
rect 5442 33056 5448 33068
rect 5500 33056 5506 33108
rect 6089 33099 6147 33105
rect 6089 33065 6101 33099
rect 6135 33096 6147 33099
rect 6270 33096 6276 33108
rect 6135 33068 6276 33096
rect 6135 33065 6147 33068
rect 6089 33059 6147 33065
rect 6270 33056 6276 33068
rect 6328 33056 6334 33108
rect 6380 33068 12388 33096
rect 6380 33028 6408 33068
rect 4908 33000 6408 33028
rect 8496 33000 9260 33028
rect 4890 32960 4896 32972
rect 1995 32932 3372 32960
rect 4724 32932 4896 32960
rect 1995 32929 2007 32932
rect 1949 32923 2007 32929
rect 3326 32852 3332 32904
rect 3384 32892 3390 32904
rect 4724 32901 4752 32932
rect 4890 32920 4896 32932
rect 4948 32960 4954 32972
rect 5258 32960 5264 32972
rect 4948 32932 5264 32960
rect 4948 32920 4954 32932
rect 5258 32920 5264 32932
rect 5316 32920 5322 32972
rect 8496 32960 8524 33000
rect 6104 32932 8524 32960
rect 8573 32963 8631 32969
rect 3973 32895 4031 32901
rect 3973 32892 3985 32895
rect 3384 32864 3985 32892
rect 3384 32852 3390 32864
rect 3973 32861 3985 32864
rect 4019 32861 4031 32895
rect 3973 32855 4031 32861
rect 4709 32895 4767 32901
rect 4709 32861 4721 32895
rect 4755 32861 4767 32895
rect 4709 32855 4767 32861
rect 4801 32895 4859 32901
rect 4801 32861 4813 32895
rect 4847 32892 4859 32895
rect 5442 32892 5448 32904
rect 4847 32864 5448 32892
rect 4847 32861 4859 32864
rect 4801 32855 4859 32861
rect 5442 32852 5448 32864
rect 5500 32852 5506 32904
rect 5534 32852 5540 32904
rect 5592 32892 5598 32904
rect 5592 32864 5637 32892
rect 5592 32852 5598 32864
rect 5902 32852 5908 32904
rect 5960 32892 5966 32904
rect 5997 32895 6055 32901
rect 5997 32892 6009 32895
rect 5960 32864 6009 32892
rect 5960 32852 5966 32864
rect 5997 32861 6009 32864
rect 6043 32861 6055 32895
rect 5997 32855 6055 32861
rect 4614 32824 4620 32836
rect 3174 32796 4620 32824
rect 4614 32784 4620 32796
rect 4672 32784 4678 32836
rect 4890 32784 4896 32836
rect 4948 32824 4954 32836
rect 6104 32824 6132 32932
rect 8573 32929 8585 32963
rect 8619 32960 8631 32963
rect 8754 32960 8760 32972
rect 8619 32932 8760 32960
rect 8619 32929 8631 32932
rect 8573 32923 8631 32929
rect 8754 32920 8760 32932
rect 8812 32960 8818 32972
rect 9122 32960 9128 32972
rect 8812 32932 9128 32960
rect 8812 32920 8818 32932
rect 9122 32920 9128 32932
rect 9180 32920 9186 32972
rect 9232 32960 9260 33000
rect 10226 32960 10232 32972
rect 9232 32932 10232 32960
rect 10226 32920 10232 32932
rect 10284 32920 10290 32972
rect 10962 32852 10968 32904
rect 11020 32892 11026 32904
rect 12360 32901 12388 33068
rect 12710 33056 12716 33108
rect 12768 33096 12774 33108
rect 14277 33099 14335 33105
rect 14277 33096 14289 33099
rect 12768 33068 14289 33096
rect 12768 33056 12774 33068
rect 14277 33065 14289 33068
rect 14323 33096 14335 33099
rect 14734 33096 14740 33108
rect 14323 33068 14740 33096
rect 14323 33065 14335 33068
rect 14277 33059 14335 33065
rect 14734 33056 14740 33068
rect 14792 33056 14798 33108
rect 13722 33028 13728 33040
rect 13372 33000 13728 33028
rect 13372 32969 13400 33000
rect 13722 32988 13728 33000
rect 13780 32988 13786 33040
rect 13357 32963 13415 32969
rect 13357 32929 13369 32963
rect 13403 32929 13415 32963
rect 13357 32923 13415 32929
rect 11425 32895 11483 32901
rect 11425 32892 11437 32895
rect 11020 32864 11437 32892
rect 11020 32852 11026 32864
rect 11425 32861 11437 32864
rect 11471 32861 11483 32895
rect 11425 32855 11483 32861
rect 12345 32895 12403 32901
rect 12345 32861 12357 32895
rect 12391 32861 12403 32895
rect 12345 32855 12403 32861
rect 4948 32796 6132 32824
rect 4948 32784 4954 32796
rect 6638 32784 6644 32836
rect 6696 32824 6702 32836
rect 8297 32827 8355 32833
rect 6696 32796 7130 32824
rect 6696 32784 6702 32796
rect 8297 32793 8309 32827
rect 8343 32824 8355 32827
rect 8343 32796 8892 32824
rect 8343 32793 8355 32796
rect 8297 32787 8355 32793
rect 3421 32759 3479 32765
rect 3421 32725 3433 32759
rect 3467 32756 3479 32759
rect 3694 32756 3700 32768
rect 3467 32728 3700 32756
rect 3467 32725 3479 32728
rect 3421 32719 3479 32725
rect 3694 32716 3700 32728
rect 3752 32716 3758 32768
rect 4157 32759 4215 32765
rect 4157 32725 4169 32759
rect 4203 32756 4215 32759
rect 4522 32756 4528 32768
rect 4203 32728 4528 32756
rect 4203 32725 4215 32728
rect 4157 32719 4215 32725
rect 4522 32716 4528 32728
rect 4580 32716 4586 32768
rect 5258 32716 5264 32768
rect 5316 32756 5322 32768
rect 6546 32756 6552 32768
rect 5316 32728 6552 32756
rect 5316 32716 5322 32728
rect 6546 32716 6552 32728
rect 6604 32716 6610 32768
rect 6822 32756 6828 32768
rect 6783 32728 6828 32756
rect 6822 32716 6828 32728
rect 6880 32716 6886 32768
rect 8864 32756 8892 32796
rect 8938 32784 8944 32836
rect 8996 32824 9002 32836
rect 10686 32824 10692 32836
rect 8996 32796 9522 32824
rect 10647 32796 10692 32824
rect 8996 32784 9002 32796
rect 10686 32784 10692 32796
rect 10744 32824 10750 32836
rect 13538 32824 13544 32836
rect 10744 32796 13400 32824
rect 13499 32796 13544 32824
rect 10744 32784 10750 32796
rect 9217 32759 9275 32765
rect 9217 32756 9229 32759
rect 8864 32728 9229 32756
rect 9217 32725 9229 32728
rect 9263 32756 9275 32759
rect 12158 32756 12164 32768
rect 9263 32728 12164 32756
rect 9263 32725 9275 32728
rect 9217 32719 9275 32725
rect 12158 32716 12164 32728
rect 12216 32716 12222 32768
rect 12434 32756 12440 32768
rect 12395 32728 12440 32756
rect 12434 32716 12440 32728
rect 12492 32716 12498 32768
rect 13372 32756 13400 32796
rect 13538 32784 13544 32796
rect 13596 32784 13602 32836
rect 13630 32784 13636 32836
rect 13688 32824 13694 32836
rect 14826 32824 14832 32836
rect 13688 32796 13733 32824
rect 14200 32796 14832 32824
rect 13688 32784 13694 32796
rect 14200 32756 14228 32796
rect 14826 32784 14832 32796
rect 14884 32784 14890 32836
rect 36354 32756 36360 32768
rect 13372 32728 14228 32756
rect 36315 32728 36360 32756
rect 36354 32716 36360 32728
rect 36412 32716 36418 32768
rect 1104 32666 36892 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 36892 32666
rect 1104 32592 36892 32614
rect 1670 32512 1676 32564
rect 1728 32552 1734 32564
rect 1946 32552 1952 32564
rect 1728 32524 1952 32552
rect 1728 32512 1734 32524
rect 1946 32512 1952 32524
rect 2004 32552 2010 32564
rect 6638 32552 6644 32564
rect 2004 32524 4016 32552
rect 2004 32512 2010 32524
rect 1688 32456 2530 32484
rect 1688 32428 1716 32456
rect 1670 32376 1676 32428
rect 1728 32376 1734 32428
rect 1765 32419 1823 32425
rect 1765 32385 1777 32419
rect 1811 32416 1823 32419
rect 2406 32416 2412 32428
rect 1811 32388 2412 32416
rect 1811 32385 1823 32388
rect 1765 32379 1823 32385
rect 2406 32376 2412 32388
rect 2464 32376 2470 32428
rect 2225 32351 2283 32357
rect 2225 32317 2237 32351
rect 2271 32348 2283 32351
rect 3694 32348 3700 32360
rect 2271 32320 2636 32348
rect 3655 32320 3700 32348
rect 2271 32317 2283 32320
rect 2225 32311 2283 32317
rect 2608 32292 2636 32320
rect 3694 32308 3700 32320
rect 3752 32308 3758 32360
rect 3988 32357 4016 32524
rect 5368 32524 5856 32552
rect 6599 32524 6644 32552
rect 4154 32376 4160 32428
rect 4212 32416 4218 32428
rect 4433 32419 4491 32425
rect 4433 32416 4445 32419
rect 4212 32388 4445 32416
rect 4212 32376 4218 32388
rect 4433 32385 4445 32388
rect 4479 32416 4491 32419
rect 4890 32416 4896 32428
rect 4479 32388 4896 32416
rect 4479 32385 4491 32388
rect 4433 32379 4491 32385
rect 4890 32376 4896 32388
rect 4948 32416 4954 32428
rect 5077 32419 5135 32425
rect 5077 32416 5089 32419
rect 4948 32388 5089 32416
rect 4948 32376 4954 32388
rect 5077 32385 5089 32388
rect 5123 32385 5135 32419
rect 5077 32379 5135 32385
rect 3973 32351 4031 32357
rect 3973 32317 3985 32351
rect 4019 32348 4031 32351
rect 4062 32348 4068 32360
rect 4019 32320 4068 32348
rect 4019 32317 4031 32320
rect 3973 32311 4031 32317
rect 4062 32308 4068 32320
rect 4120 32308 4126 32360
rect 2590 32240 2596 32292
rect 2648 32240 2654 32292
rect 5169 32283 5227 32289
rect 5169 32249 5181 32283
rect 5215 32280 5227 32283
rect 5368 32280 5396 32524
rect 5828 32484 5856 32524
rect 6638 32512 6644 32524
rect 6696 32512 6702 32564
rect 7006 32512 7012 32564
rect 7064 32552 7070 32564
rect 7285 32555 7343 32561
rect 7285 32552 7297 32555
rect 7064 32524 7297 32552
rect 7064 32512 7070 32524
rect 7285 32521 7297 32524
rect 7331 32521 7343 32555
rect 8938 32552 8944 32564
rect 7285 32515 7343 32521
rect 7576 32524 8944 32552
rect 7466 32484 7472 32496
rect 5828 32456 7472 32484
rect 7466 32444 7472 32456
rect 7524 32444 7530 32496
rect 5534 32376 5540 32428
rect 5592 32416 5598 32428
rect 5721 32419 5779 32425
rect 5721 32416 5733 32419
rect 5592 32388 5733 32416
rect 5592 32376 5598 32388
rect 5721 32385 5733 32388
rect 5767 32416 5779 32419
rect 6549 32419 6607 32425
rect 6549 32416 6561 32419
rect 5767 32388 6561 32416
rect 5767 32385 5779 32388
rect 5721 32379 5779 32385
rect 6549 32385 6561 32388
rect 6595 32416 6607 32419
rect 7190 32416 7196 32428
rect 6595 32388 7196 32416
rect 6595 32385 6607 32388
rect 6549 32379 6607 32385
rect 7190 32376 7196 32388
rect 7248 32376 7254 32428
rect 7282 32376 7288 32428
rect 7340 32416 7346 32428
rect 7377 32419 7435 32425
rect 7377 32416 7389 32419
rect 7340 32388 7389 32416
rect 7340 32376 7346 32388
rect 7377 32385 7389 32388
rect 7423 32385 7435 32419
rect 7377 32379 7435 32385
rect 5813 32351 5871 32357
rect 5813 32317 5825 32351
rect 5859 32348 5871 32351
rect 7576 32348 7604 32524
rect 8938 32512 8944 32524
rect 8996 32512 9002 32564
rect 9122 32512 9128 32564
rect 9180 32552 9186 32564
rect 12710 32552 12716 32564
rect 9180 32524 10180 32552
rect 9180 32512 9186 32524
rect 7742 32444 7748 32496
rect 7800 32484 7806 32496
rect 7800 32456 8694 32484
rect 7800 32444 7806 32456
rect 10152 32425 10180 32524
rect 10704 32524 12716 32552
rect 10226 32444 10232 32496
rect 10284 32484 10290 32496
rect 10704 32484 10732 32524
rect 12710 32512 12716 32524
rect 12768 32512 12774 32564
rect 12802 32512 12808 32564
rect 12860 32552 12866 32564
rect 13170 32552 13176 32564
rect 12860 32524 13176 32552
rect 12860 32512 12866 32524
rect 13170 32512 13176 32524
rect 13228 32552 13234 32564
rect 13228 32524 14228 32552
rect 13228 32512 13234 32524
rect 10284 32456 10732 32484
rect 10284 32444 10290 32456
rect 12434 32444 12440 32496
rect 12492 32484 12498 32496
rect 14200 32493 14228 32524
rect 13633 32487 13691 32493
rect 13633 32484 13645 32487
rect 12492 32456 13645 32484
rect 12492 32444 12498 32456
rect 13633 32453 13645 32456
rect 13679 32453 13691 32487
rect 13633 32447 13691 32453
rect 14185 32487 14243 32493
rect 14185 32453 14197 32487
rect 14231 32453 14243 32487
rect 14185 32447 14243 32453
rect 10137 32419 10195 32425
rect 10137 32385 10149 32419
rect 10183 32416 10195 32419
rect 10318 32416 10324 32428
rect 10183 32388 10324 32416
rect 10183 32385 10195 32388
rect 10137 32379 10195 32385
rect 10318 32376 10324 32388
rect 10376 32376 10382 32428
rect 10778 32376 10784 32428
rect 10836 32416 10842 32428
rect 12161 32419 12219 32425
rect 12161 32416 12173 32419
rect 10836 32388 12173 32416
rect 10836 32376 10842 32388
rect 12161 32385 12173 32388
rect 12207 32385 12219 32419
rect 12161 32379 12219 32385
rect 12805 32419 12863 32425
rect 12805 32385 12817 32419
rect 12851 32385 12863 32419
rect 12805 32379 12863 32385
rect 5859 32320 7604 32348
rect 8113 32351 8171 32357
rect 5859 32317 5871 32320
rect 5813 32311 5871 32317
rect 8113 32317 8125 32351
rect 8159 32348 8171 32351
rect 8662 32348 8668 32360
rect 8159 32320 8668 32348
rect 8159 32317 8171 32320
rect 8113 32311 8171 32317
rect 8662 32308 8668 32320
rect 8720 32308 8726 32360
rect 9490 32308 9496 32360
rect 9548 32348 9554 32360
rect 9861 32351 9919 32357
rect 9861 32348 9873 32351
rect 9548 32320 9873 32348
rect 9548 32308 9554 32320
rect 9861 32317 9873 32320
rect 9907 32348 9919 32351
rect 12820 32348 12848 32379
rect 9907 32320 12848 32348
rect 13541 32351 13599 32357
rect 9907 32317 9919 32320
rect 9861 32311 9919 32317
rect 13541 32317 13553 32351
rect 13587 32348 13599 32351
rect 13722 32348 13728 32360
rect 13587 32320 13728 32348
rect 13587 32317 13599 32320
rect 13541 32311 13599 32317
rect 13722 32308 13728 32320
rect 13780 32308 13786 32360
rect 36078 32348 36084 32360
rect 36039 32320 36084 32348
rect 36078 32308 36084 32320
rect 36136 32308 36142 32360
rect 36354 32348 36360 32360
rect 36315 32320 36360 32348
rect 36354 32308 36360 32320
rect 36412 32308 36418 32360
rect 5215 32252 5396 32280
rect 5215 32249 5227 32252
rect 5169 32243 5227 32249
rect 10318 32240 10324 32292
rect 10376 32280 10382 32292
rect 10689 32283 10747 32289
rect 10689 32280 10701 32283
rect 10376 32252 10701 32280
rect 10376 32240 10382 32252
rect 10689 32249 10701 32252
rect 10735 32280 10747 32283
rect 10962 32280 10968 32292
rect 10735 32252 10968 32280
rect 10735 32249 10747 32252
rect 10689 32243 10747 32249
rect 10962 32240 10968 32252
rect 11020 32240 11026 32292
rect 12253 32283 12311 32289
rect 12253 32249 12265 32283
rect 12299 32280 12311 32283
rect 13998 32280 14004 32292
rect 12299 32252 14004 32280
rect 12299 32249 12311 32252
rect 12253 32243 12311 32249
rect 13998 32240 14004 32252
rect 14056 32240 14062 32292
rect 1673 32215 1731 32221
rect 1673 32181 1685 32215
rect 1719 32212 1731 32215
rect 3970 32212 3976 32224
rect 1719 32184 3976 32212
rect 1719 32181 1731 32184
rect 1673 32175 1731 32181
rect 3970 32172 3976 32184
rect 4028 32172 4034 32224
rect 4525 32215 4583 32221
rect 4525 32181 4537 32215
rect 4571 32212 4583 32215
rect 8478 32212 8484 32224
rect 4571 32184 8484 32212
rect 4571 32181 4583 32184
rect 4525 32175 4583 32181
rect 8478 32172 8484 32184
rect 8536 32172 8542 32224
rect 12897 32215 12955 32221
rect 12897 32181 12909 32215
rect 12943 32212 12955 32215
rect 14182 32212 14188 32224
rect 12943 32184 14188 32212
rect 12943 32181 12955 32184
rect 12897 32175 12955 32181
rect 14182 32172 14188 32184
rect 14240 32172 14246 32224
rect 1104 32122 36892 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 36892 32122
rect 1104 32048 36892 32070
rect 3234 31968 3240 32020
rect 3292 32008 3298 32020
rect 4065 32011 4123 32017
rect 4065 32008 4077 32011
rect 3292 31980 4077 32008
rect 3292 31968 3298 31980
rect 4065 31977 4077 31980
rect 4111 31977 4123 32011
rect 4065 31971 4123 31977
rect 4614 31968 4620 32020
rect 4672 32008 4678 32020
rect 4709 32011 4767 32017
rect 4709 32008 4721 32011
rect 4672 31980 4721 32008
rect 4672 31968 4678 31980
rect 4709 31977 4721 31980
rect 4755 31977 4767 32011
rect 4709 31971 4767 31977
rect 5353 32011 5411 32017
rect 5353 31977 5365 32011
rect 5399 32008 5411 32011
rect 8386 32008 8392 32020
rect 5399 31980 8392 32008
rect 5399 31977 5411 31980
rect 5353 31971 5411 31977
rect 8386 31968 8392 31980
rect 8444 31968 8450 32020
rect 9122 32008 9128 32020
rect 9083 31980 9128 32008
rect 9122 31968 9128 31980
rect 9180 31968 9186 32020
rect 10410 31968 10416 32020
rect 10468 32008 10474 32020
rect 10468 31980 12756 32008
rect 10468 31968 10474 31980
rect 2961 31943 3019 31949
rect 2961 31909 2973 31943
rect 3007 31940 3019 31943
rect 4798 31940 4804 31952
rect 3007 31912 4804 31940
rect 3007 31909 3019 31912
rect 2961 31903 3019 31909
rect 4798 31900 4804 31912
rect 4856 31900 4862 31952
rect 5258 31940 5264 31952
rect 5184 31912 5264 31940
rect 2222 31832 2228 31884
rect 2280 31872 2286 31884
rect 2409 31875 2467 31881
rect 2409 31872 2421 31875
rect 2280 31844 2421 31872
rect 2280 31832 2286 31844
rect 2409 31841 2421 31844
rect 2455 31841 2467 31875
rect 2409 31835 2467 31841
rect 3694 31832 3700 31884
rect 3752 31872 3758 31884
rect 4890 31872 4896 31884
rect 3752 31844 4896 31872
rect 3752 31832 3758 31844
rect 4890 31832 4896 31844
rect 4948 31832 4954 31884
rect 2130 31804 2136 31816
rect 2091 31776 2136 31804
rect 2130 31764 2136 31776
rect 2188 31764 2194 31816
rect 2869 31807 2927 31813
rect 2869 31773 2881 31807
rect 2915 31804 2927 31807
rect 2958 31804 2964 31816
rect 2915 31776 2964 31804
rect 2915 31773 2927 31776
rect 2869 31767 2927 31773
rect 2958 31764 2964 31776
rect 3016 31804 3022 31816
rect 3878 31804 3884 31816
rect 3016 31776 3884 31804
rect 3016 31764 3022 31776
rect 3878 31764 3884 31776
rect 3936 31764 3942 31816
rect 4157 31807 4215 31813
rect 4157 31773 4169 31807
rect 4203 31804 4215 31807
rect 4614 31804 4620 31816
rect 4203 31776 4620 31804
rect 4203 31773 4215 31776
rect 4157 31767 4215 31773
rect 4614 31764 4620 31776
rect 4672 31764 4678 31816
rect 4801 31807 4859 31813
rect 4801 31773 4813 31807
rect 4847 31804 4859 31807
rect 5074 31804 5080 31816
rect 4847 31776 5080 31804
rect 4847 31773 4859 31776
rect 4801 31767 4859 31773
rect 5074 31764 5080 31776
rect 5132 31804 5138 31816
rect 5184 31804 5212 31912
rect 5258 31900 5264 31912
rect 5316 31900 5322 31952
rect 5997 31943 6055 31949
rect 5997 31909 6009 31943
rect 6043 31940 6055 31943
rect 6454 31940 6460 31952
rect 6043 31912 6460 31940
rect 6043 31909 6055 31912
rect 5997 31903 6055 31909
rect 6454 31900 6460 31912
rect 6512 31900 6518 31952
rect 6546 31900 6552 31952
rect 6604 31940 6610 31952
rect 8481 31943 8539 31949
rect 6604 31912 6868 31940
rect 6604 31900 6610 31912
rect 5810 31832 5816 31884
rect 5868 31872 5874 31884
rect 6086 31872 6092 31884
rect 5868 31844 6092 31872
rect 5868 31832 5874 31844
rect 6086 31832 6092 31844
rect 6144 31872 6150 31884
rect 6733 31875 6791 31881
rect 6733 31872 6745 31875
rect 6144 31844 6745 31872
rect 6144 31832 6150 31844
rect 6733 31841 6745 31844
rect 6779 31841 6791 31875
rect 6840 31872 6868 31912
rect 8481 31909 8493 31943
rect 8527 31940 8539 31943
rect 10686 31940 10692 31952
rect 8527 31912 10692 31940
rect 8527 31909 8539 31912
rect 8481 31903 8539 31909
rect 10686 31900 10692 31912
rect 10744 31900 10750 31952
rect 12728 31940 12756 31980
rect 35618 31968 35624 32020
rect 35676 32008 35682 32020
rect 35897 32011 35955 32017
rect 35897 32008 35909 32011
rect 35676 31980 35909 32008
rect 35676 31968 35682 31980
rect 35897 31977 35909 31980
rect 35943 31977 35955 32011
rect 35897 31971 35955 31977
rect 12728 31912 12848 31940
rect 6840 31844 10180 31872
rect 6733 31835 6791 31841
rect 5132 31776 5212 31804
rect 5261 31807 5319 31813
rect 5132 31764 5138 31776
rect 5261 31773 5273 31807
rect 5307 31773 5319 31807
rect 5261 31767 5319 31773
rect 4632 31736 4660 31764
rect 5276 31736 5304 31767
rect 5442 31764 5448 31816
rect 5500 31804 5506 31816
rect 5905 31807 5963 31813
rect 5905 31804 5917 31807
rect 5500 31776 5917 31804
rect 5500 31764 5506 31776
rect 5905 31773 5917 31776
rect 5951 31804 5963 31807
rect 6546 31804 6552 31816
rect 5951 31776 6552 31804
rect 5951 31773 5963 31776
rect 5905 31767 5963 31773
rect 6546 31764 6552 31776
rect 6604 31764 6610 31816
rect 9766 31764 9772 31816
rect 9824 31804 9830 31816
rect 9861 31807 9919 31813
rect 9861 31804 9873 31807
rect 9824 31776 9873 31804
rect 9824 31764 9830 31776
rect 9861 31773 9873 31776
rect 9907 31773 9919 31807
rect 9861 31767 9919 31773
rect 9950 31764 9956 31816
rect 10008 31804 10014 31816
rect 10152 31804 10180 31844
rect 10594 31832 10600 31884
rect 10652 31872 10658 31884
rect 11517 31875 11575 31881
rect 10652 31844 11468 31872
rect 10652 31832 10658 31844
rect 10781 31807 10839 31813
rect 10781 31804 10793 31807
rect 10008 31776 10053 31804
rect 10152 31776 10793 31804
rect 10008 31764 10014 31776
rect 10781 31773 10793 31776
rect 10827 31773 10839 31807
rect 10781 31767 10839 31773
rect 10873 31807 10931 31813
rect 10873 31773 10885 31807
rect 10919 31804 10931 31807
rect 11330 31804 11336 31816
rect 10919 31776 11336 31804
rect 10919 31773 10931 31776
rect 10873 31767 10931 31773
rect 11330 31764 11336 31776
rect 11388 31764 11394 31816
rect 11440 31813 11468 31844
rect 11517 31841 11529 31875
rect 11563 31872 11575 31875
rect 12710 31872 12716 31884
rect 11563 31844 12716 31872
rect 11563 31841 11575 31844
rect 11517 31835 11575 31841
rect 12710 31832 12716 31844
rect 12768 31832 12774 31884
rect 12820 31813 12848 31912
rect 13538 31872 13544 31884
rect 13499 31844 13544 31872
rect 13538 31832 13544 31844
rect 13596 31832 13602 31884
rect 11425 31807 11483 31813
rect 11425 31773 11437 31807
rect 11471 31773 11483 31807
rect 11425 31767 11483 31773
rect 12069 31807 12127 31813
rect 12069 31773 12081 31807
rect 12115 31773 12127 31807
rect 12069 31767 12127 31773
rect 12805 31807 12863 31813
rect 12805 31773 12817 31807
rect 12851 31773 12863 31807
rect 12805 31767 12863 31773
rect 5994 31736 6000 31748
rect 4632 31708 6000 31736
rect 5994 31696 6000 31708
rect 6052 31696 6058 31748
rect 7006 31736 7012 31748
rect 6967 31708 7012 31736
rect 7006 31696 7012 31708
rect 7064 31696 7070 31748
rect 7282 31696 7288 31748
rect 7340 31736 7346 31748
rect 7340 31708 7498 31736
rect 7340 31696 7346 31708
rect 11054 31696 11060 31748
rect 11112 31736 11118 31748
rect 12084 31736 12112 31767
rect 13354 31764 13360 31816
rect 13412 31804 13418 31816
rect 13633 31807 13691 31813
rect 13633 31804 13645 31807
rect 13412 31776 13645 31804
rect 13412 31764 13418 31776
rect 13633 31773 13645 31776
rect 13679 31773 13691 31807
rect 13633 31767 13691 31773
rect 14090 31764 14096 31816
rect 14148 31804 14154 31816
rect 14645 31807 14703 31813
rect 14645 31804 14657 31807
rect 14148 31776 14657 31804
rect 14148 31764 14154 31776
rect 14645 31773 14657 31776
rect 14691 31773 14703 31807
rect 14645 31767 14703 31773
rect 14737 31807 14795 31813
rect 14737 31773 14749 31807
rect 14783 31804 14795 31807
rect 15378 31804 15384 31816
rect 14783 31776 15384 31804
rect 14783 31773 14795 31776
rect 14737 31767 14795 31773
rect 15378 31764 15384 31776
rect 15436 31764 15442 31816
rect 19426 31764 19432 31816
rect 19484 31804 19490 31816
rect 22741 31807 22799 31813
rect 22741 31804 22753 31807
rect 19484 31776 22753 31804
rect 19484 31764 19490 31776
rect 22741 31773 22753 31776
rect 22787 31773 22799 31807
rect 22741 31767 22799 31773
rect 22833 31807 22891 31813
rect 22833 31773 22845 31807
rect 22879 31804 22891 31807
rect 23385 31807 23443 31813
rect 23385 31804 23397 31807
rect 22879 31776 23397 31804
rect 22879 31773 22891 31776
rect 22833 31767 22891 31773
rect 23385 31773 23397 31776
rect 23431 31804 23443 31807
rect 27890 31804 27896 31816
rect 23431 31776 27896 31804
rect 23431 31773 23443 31776
rect 23385 31767 23443 31773
rect 27890 31764 27896 31776
rect 27948 31764 27954 31816
rect 35986 31764 35992 31816
rect 36044 31804 36050 31816
rect 36081 31807 36139 31813
rect 36081 31804 36093 31807
rect 36044 31776 36093 31804
rect 36044 31764 36050 31776
rect 36081 31773 36093 31776
rect 36127 31773 36139 31807
rect 36081 31767 36139 31773
rect 11112 31708 12112 31736
rect 11112 31696 11118 31708
rect 13446 31696 13452 31748
rect 13504 31736 13510 31748
rect 13814 31736 13820 31748
rect 13504 31708 13820 31736
rect 13504 31696 13510 31708
rect 13814 31696 13820 31708
rect 13872 31696 13878 31748
rect 4430 31628 4436 31680
rect 4488 31668 4494 31680
rect 9582 31668 9588 31680
rect 4488 31640 9588 31668
rect 4488 31628 4494 31640
rect 9582 31628 9588 31640
rect 9640 31628 9646 31680
rect 11882 31628 11888 31680
rect 11940 31668 11946 31680
rect 12161 31671 12219 31677
rect 12161 31668 12173 31671
rect 11940 31640 12173 31668
rect 11940 31628 11946 31640
rect 12161 31637 12173 31640
rect 12207 31637 12219 31671
rect 12161 31631 12219 31637
rect 12897 31671 12955 31677
rect 12897 31637 12909 31671
rect 12943 31668 12955 31671
rect 13722 31668 13728 31680
rect 12943 31640 13728 31668
rect 12943 31637 12955 31640
rect 12897 31631 12955 31637
rect 13722 31628 13728 31640
rect 13780 31628 13786 31680
rect 1104 31578 36892 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 36892 31578
rect 1104 31504 36892 31526
rect 4706 31424 4712 31476
rect 4764 31464 4770 31476
rect 5074 31464 5080 31476
rect 4764 31436 5080 31464
rect 4764 31424 4770 31436
rect 5074 31424 5080 31436
rect 5132 31424 5138 31476
rect 5166 31424 5172 31476
rect 5224 31464 5230 31476
rect 5350 31464 5356 31476
rect 5224 31436 5356 31464
rect 5224 31424 5230 31436
rect 5350 31424 5356 31436
rect 5408 31424 5414 31476
rect 5718 31424 5724 31476
rect 5776 31464 5782 31476
rect 6641 31467 6699 31473
rect 6641 31464 6653 31467
rect 5776 31436 6653 31464
rect 5776 31424 5782 31436
rect 6641 31433 6653 31436
rect 6687 31433 6699 31467
rect 7282 31464 7288 31476
rect 7243 31436 7288 31464
rect 6641 31427 6699 31433
rect 7282 31424 7288 31436
rect 7340 31424 7346 31476
rect 7926 31464 7932 31476
rect 7887 31436 7932 31464
rect 7926 31424 7932 31436
rect 7984 31424 7990 31476
rect 9122 31464 9128 31476
rect 8864 31436 9128 31464
rect 8864 31408 8892 31436
rect 9122 31424 9128 31436
rect 9180 31424 9186 31476
rect 9582 31424 9588 31476
rect 9640 31464 9646 31476
rect 36078 31464 36084 31476
rect 9640 31436 36084 31464
rect 9640 31424 9646 31436
rect 36078 31424 36084 31436
rect 36136 31424 36142 31476
rect 3970 31396 3976 31408
rect 3450 31368 3976 31396
rect 3970 31356 3976 31368
rect 4028 31356 4034 31408
rect 4430 31396 4436 31408
rect 4391 31368 4436 31396
rect 4430 31356 4436 31368
rect 4488 31356 4494 31408
rect 8846 31396 8852 31408
rect 8496 31368 8852 31396
rect 1946 31328 1952 31340
rect 1907 31300 1952 31328
rect 1946 31288 1952 31300
rect 2004 31288 2010 31340
rect 5718 31328 5724 31340
rect 5566 31300 5724 31328
rect 5718 31288 5724 31300
rect 5776 31288 5782 31340
rect 5994 31288 6000 31340
rect 6052 31328 6058 31340
rect 6549 31331 6607 31337
rect 6549 31328 6561 31331
rect 6052 31300 6561 31328
rect 6052 31288 6058 31300
rect 6549 31297 6561 31300
rect 6595 31297 6607 31331
rect 6549 31291 6607 31297
rect 7193 31331 7251 31337
rect 7193 31297 7205 31331
rect 7239 31297 7251 31331
rect 7193 31291 7251 31297
rect 2225 31263 2283 31269
rect 2225 31229 2237 31263
rect 2271 31260 2283 31263
rect 2590 31260 2596 31272
rect 2271 31232 2596 31260
rect 2271 31229 2283 31232
rect 2225 31223 2283 31229
rect 2590 31220 2596 31232
rect 2648 31220 2654 31272
rect 4154 31260 4160 31272
rect 4115 31232 4160 31260
rect 4154 31220 4160 31232
rect 4212 31220 4218 31272
rect 5442 31260 5448 31272
rect 4264 31232 5448 31260
rect 3878 31152 3884 31204
rect 3936 31192 3942 31204
rect 4264 31192 4292 31232
rect 5442 31220 5448 31232
rect 5500 31260 5506 31272
rect 7208 31260 7236 31291
rect 7374 31288 7380 31340
rect 7432 31328 7438 31340
rect 7837 31331 7895 31337
rect 7837 31328 7849 31331
rect 7432 31300 7849 31328
rect 7432 31288 7438 31300
rect 7837 31297 7849 31300
rect 7883 31297 7895 31331
rect 7837 31291 7895 31297
rect 8496 31269 8524 31368
rect 8846 31356 8852 31368
rect 8904 31356 8910 31408
rect 9214 31356 9220 31408
rect 9272 31356 9278 31408
rect 11330 31356 11336 31408
rect 11388 31396 11394 31408
rect 12253 31399 12311 31405
rect 12253 31396 12265 31399
rect 11388 31368 12265 31396
rect 11388 31356 11394 31368
rect 12253 31365 12265 31368
rect 12299 31365 12311 31399
rect 12802 31396 12808 31408
rect 12763 31368 12808 31396
rect 12253 31359 12311 31365
rect 12802 31356 12808 31368
rect 12860 31356 12866 31408
rect 14182 31396 14188 31408
rect 14143 31368 14188 31396
rect 14182 31356 14188 31368
rect 14240 31356 14246 31408
rect 15378 31396 15384 31408
rect 15339 31368 15384 31396
rect 15378 31356 15384 31368
rect 15436 31356 15442 31408
rect 15473 31399 15531 31405
rect 15473 31365 15485 31399
rect 15519 31396 15531 31399
rect 19426 31396 19432 31408
rect 15519 31368 19432 31396
rect 15519 31365 15531 31368
rect 15473 31359 15531 31365
rect 19426 31356 19432 31368
rect 19484 31356 19490 31408
rect 10781 31331 10839 31337
rect 10781 31297 10793 31331
rect 10827 31297 10839 31331
rect 10781 31291 10839 31297
rect 5500 31232 7236 31260
rect 8481 31263 8539 31269
rect 5500 31220 5506 31232
rect 8481 31229 8493 31263
rect 8527 31229 8539 31263
rect 8757 31263 8815 31269
rect 8757 31260 8769 31263
rect 8481 31223 8539 31229
rect 8588 31232 8769 31260
rect 3936 31164 4292 31192
rect 5905 31195 5963 31201
rect 3936 31152 3942 31164
rect 5905 31161 5917 31195
rect 5951 31192 5963 31195
rect 8588 31192 8616 31232
rect 8757 31229 8769 31232
rect 8803 31229 8815 31263
rect 8757 31223 8815 31229
rect 9122 31220 9128 31272
rect 9180 31260 9186 31272
rect 10796 31260 10824 31291
rect 9180 31232 10824 31260
rect 12161 31263 12219 31269
rect 9180 31220 9186 31232
rect 12161 31229 12173 31263
rect 12207 31260 12219 31263
rect 12618 31260 12624 31272
rect 12207 31232 12624 31260
rect 12207 31229 12219 31232
rect 12161 31223 12219 31229
rect 12618 31220 12624 31232
rect 12676 31220 12682 31272
rect 12802 31220 12808 31272
rect 12860 31260 12866 31272
rect 13265 31263 13323 31269
rect 13265 31260 13277 31263
rect 12860 31232 13277 31260
rect 12860 31220 12866 31232
rect 13265 31229 13277 31232
rect 13311 31229 13323 31263
rect 13265 31223 13323 31229
rect 14277 31263 14335 31269
rect 14277 31229 14289 31263
rect 14323 31260 14335 31263
rect 15194 31260 15200 31272
rect 14323 31232 15200 31260
rect 14323 31229 14335 31232
rect 14277 31223 14335 31229
rect 15194 31220 15200 31232
rect 15252 31220 15258 31272
rect 5951 31164 8616 31192
rect 5951 31161 5963 31164
rect 5905 31155 5963 31161
rect 3694 31124 3700 31136
rect 3655 31096 3700 31124
rect 3694 31084 3700 31096
rect 3752 31084 3758 31136
rect 4430 31084 4436 31136
rect 4488 31124 4494 31136
rect 5442 31124 5448 31136
rect 4488 31096 5448 31124
rect 4488 31084 4494 31096
rect 5442 31084 5448 31096
rect 5500 31084 5506 31136
rect 8588 31124 8616 31164
rect 14921 31195 14979 31201
rect 14921 31161 14933 31195
rect 14967 31161 14979 31195
rect 14921 31155 14979 31161
rect 10042 31124 10048 31136
rect 8588 31096 10048 31124
rect 10042 31084 10048 31096
rect 10100 31084 10106 31136
rect 10229 31127 10287 31133
rect 10229 31093 10241 31127
rect 10275 31124 10287 31127
rect 10410 31124 10416 31136
rect 10275 31096 10416 31124
rect 10275 31093 10287 31096
rect 10229 31087 10287 31093
rect 10410 31084 10416 31096
rect 10468 31084 10474 31136
rect 10873 31127 10931 31133
rect 10873 31093 10885 31127
rect 10919 31124 10931 31127
rect 10962 31124 10968 31136
rect 10919 31096 10968 31124
rect 10919 31093 10931 31096
rect 10873 31087 10931 31093
rect 10962 31084 10968 31096
rect 11020 31084 11026 31136
rect 11422 31084 11428 31136
rect 11480 31124 11486 31136
rect 12342 31124 12348 31136
rect 11480 31096 12348 31124
rect 11480 31084 11486 31096
rect 12342 31084 12348 31096
rect 12400 31124 12406 31136
rect 14936 31124 14964 31155
rect 12400 31096 14964 31124
rect 12400 31084 12406 31096
rect 1104 31034 36892 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 36892 31034
rect 1104 30960 36892 30982
rect 4065 30923 4123 30929
rect 4065 30889 4077 30923
rect 4111 30920 4123 30923
rect 6454 30920 6460 30932
rect 4111 30892 6460 30920
rect 4111 30889 4123 30892
rect 4065 30883 4123 30889
rect 6454 30880 6460 30892
rect 6512 30880 6518 30932
rect 8315 30923 8373 30929
rect 8315 30889 8327 30923
rect 8361 30920 8373 30923
rect 9125 30923 9183 30929
rect 9125 30920 9137 30923
rect 8361 30892 9137 30920
rect 8361 30889 8373 30892
rect 8315 30883 8373 30889
rect 9125 30889 9137 30892
rect 9171 30920 9183 30923
rect 10778 30920 10784 30932
rect 9171 30892 10784 30920
rect 9171 30889 9183 30892
rect 9125 30883 9183 30889
rect 10778 30880 10784 30892
rect 10836 30880 10842 30932
rect 1857 30787 1915 30793
rect 1857 30753 1869 30787
rect 1903 30784 1915 30787
rect 3053 30787 3111 30793
rect 1903 30756 2774 30784
rect 1903 30753 1915 30756
rect 1857 30747 1915 30753
rect 2317 30719 2375 30725
rect 2317 30685 2329 30719
rect 2363 30716 2375 30719
rect 2406 30716 2412 30728
rect 2363 30688 2412 30716
rect 2363 30685 2375 30688
rect 2317 30679 2375 30685
rect 2406 30676 2412 30688
rect 2464 30676 2470 30728
rect 1486 30608 1492 30660
rect 1544 30648 1550 30660
rect 1673 30651 1731 30657
rect 1673 30648 1685 30651
rect 1544 30620 1685 30648
rect 1544 30608 1550 30620
rect 1673 30617 1685 30620
rect 1719 30617 1731 30651
rect 2746 30648 2774 30756
rect 3053 30753 3065 30787
rect 3099 30784 3111 30787
rect 8294 30784 8300 30796
rect 3099 30756 8300 30784
rect 3099 30753 3111 30756
rect 3053 30747 3111 30753
rect 8294 30744 8300 30756
rect 8352 30744 8358 30796
rect 8573 30787 8631 30793
rect 8573 30753 8585 30787
rect 8619 30784 8631 30787
rect 8846 30784 8852 30796
rect 8619 30756 8852 30784
rect 8619 30753 8631 30756
rect 8573 30747 8631 30753
rect 8846 30744 8852 30756
rect 8904 30784 8910 30796
rect 10873 30787 10931 30793
rect 10873 30784 10885 30787
rect 8904 30756 10885 30784
rect 8904 30744 8910 30756
rect 10873 30753 10885 30756
rect 10919 30784 10931 30787
rect 11146 30784 11152 30796
rect 10919 30756 11152 30784
rect 10919 30753 10931 30756
rect 10873 30747 10931 30753
rect 11146 30744 11152 30756
rect 11204 30744 11210 30796
rect 14366 30784 14372 30796
rect 14327 30756 14372 30784
rect 14366 30744 14372 30756
rect 14424 30744 14430 30796
rect 2958 30716 2964 30728
rect 2919 30688 2964 30716
rect 2958 30676 2964 30688
rect 3016 30676 3022 30728
rect 5810 30676 5816 30728
rect 5868 30716 5874 30728
rect 5868 30688 5913 30716
rect 5868 30676 5874 30688
rect 7190 30676 7196 30728
rect 7248 30676 7254 30728
rect 13078 30676 13084 30728
rect 13136 30716 13142 30728
rect 13265 30719 13323 30725
rect 13265 30716 13277 30719
rect 13136 30688 13277 30716
rect 13136 30676 13142 30688
rect 13265 30685 13277 30688
rect 13311 30685 13323 30719
rect 13265 30679 13323 30685
rect 15470 30676 15476 30728
rect 15528 30716 15534 30728
rect 15657 30719 15715 30725
rect 15657 30716 15669 30719
rect 15528 30688 15669 30716
rect 15528 30676 15534 30688
rect 15657 30685 15669 30688
rect 15703 30716 15715 30719
rect 15838 30716 15844 30728
rect 15703 30688 15844 30716
rect 15703 30685 15715 30688
rect 15657 30679 15715 30685
rect 15838 30676 15844 30688
rect 15896 30676 15902 30728
rect 2746 30620 4200 30648
rect 1673 30611 1731 30617
rect 2409 30583 2467 30589
rect 2409 30549 2421 30583
rect 2455 30580 2467 30583
rect 3050 30580 3056 30592
rect 2455 30552 3056 30580
rect 2455 30549 2467 30552
rect 2409 30543 2467 30549
rect 3050 30540 3056 30552
rect 3108 30540 3114 30592
rect 4172 30580 4200 30620
rect 4798 30608 4804 30660
rect 4856 30608 4862 30660
rect 5534 30648 5540 30660
rect 5495 30620 5540 30648
rect 5534 30608 5540 30620
rect 5592 30608 5598 30660
rect 5644 30620 6960 30648
rect 5644 30580 5672 30620
rect 4172 30552 5672 30580
rect 6638 30540 6644 30592
rect 6696 30580 6702 30592
rect 6825 30583 6883 30589
rect 6825 30580 6837 30583
rect 6696 30552 6837 30580
rect 6696 30540 6702 30552
rect 6825 30549 6837 30552
rect 6871 30549 6883 30583
rect 6932 30580 6960 30620
rect 8404 30620 9260 30648
rect 8404 30580 8432 30620
rect 6932 30552 8432 30580
rect 9232 30580 9260 30620
rect 9306 30608 9312 30660
rect 9364 30648 9370 30660
rect 10594 30648 10600 30660
rect 9364 30620 9430 30648
rect 10555 30620 10600 30648
rect 9364 30608 9370 30620
rect 10594 30608 10600 30620
rect 10652 30608 10658 30660
rect 11330 30608 11336 30660
rect 11388 30648 11394 30660
rect 11793 30651 11851 30657
rect 11793 30648 11805 30651
rect 11388 30620 11805 30648
rect 11388 30608 11394 30620
rect 11793 30617 11805 30620
rect 11839 30617 11851 30651
rect 11793 30611 11851 30617
rect 11882 30608 11888 30660
rect 11940 30648 11946 30660
rect 12802 30648 12808 30660
rect 11940 30620 11985 30648
rect 12763 30620 12808 30648
rect 11940 30608 11946 30620
rect 12802 30608 12808 30620
rect 12860 30608 12866 30660
rect 14182 30648 14188 30660
rect 13004 30620 14188 30648
rect 13004 30580 13032 30620
rect 14182 30608 14188 30620
rect 14240 30608 14246 30660
rect 14461 30651 14519 30657
rect 14461 30617 14473 30651
rect 14507 30617 14519 30651
rect 14461 30611 14519 30617
rect 15013 30651 15071 30657
rect 15013 30617 15025 30651
rect 15059 30648 15071 30651
rect 15194 30648 15200 30660
rect 15059 30620 15200 30648
rect 15059 30617 15071 30620
rect 15013 30611 15071 30617
rect 9232 30552 13032 30580
rect 6825 30543 6883 30549
rect 13078 30540 13084 30592
rect 13136 30580 13142 30592
rect 13357 30583 13415 30589
rect 13357 30580 13369 30583
rect 13136 30552 13369 30580
rect 13136 30540 13142 30552
rect 13357 30549 13369 30552
rect 13403 30549 13415 30583
rect 13357 30543 13415 30549
rect 13722 30540 13728 30592
rect 13780 30580 13786 30592
rect 14476 30580 14504 30611
rect 15194 30608 15200 30620
rect 15252 30648 15258 30660
rect 16206 30648 16212 30660
rect 15252 30620 16212 30648
rect 15252 30608 15258 30620
rect 16206 30608 16212 30620
rect 16264 30608 16270 30660
rect 15562 30580 15568 30592
rect 13780 30552 14504 30580
rect 15523 30552 15568 30580
rect 13780 30540 13786 30552
rect 15562 30540 15568 30552
rect 15620 30540 15626 30592
rect 15838 30540 15844 30592
rect 15896 30580 15902 30592
rect 16117 30583 16175 30589
rect 16117 30580 16129 30583
rect 15896 30552 16129 30580
rect 15896 30540 15902 30552
rect 16117 30549 16129 30552
rect 16163 30549 16175 30583
rect 16117 30543 16175 30549
rect 1104 30490 36892 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 36892 30490
rect 1104 30416 36892 30438
rect 3329 30379 3387 30385
rect 3329 30345 3341 30379
rect 3375 30376 3387 30379
rect 7926 30376 7932 30388
rect 3375 30348 7932 30376
rect 3375 30345 3387 30348
rect 3329 30339 3387 30345
rect 7926 30336 7932 30348
rect 7984 30336 7990 30388
rect 8294 30336 8300 30388
rect 8352 30336 8358 30388
rect 12802 30336 12808 30388
rect 12860 30376 12866 30388
rect 19334 30376 19340 30388
rect 12860 30348 19340 30376
rect 12860 30336 12866 30348
rect 19334 30336 19340 30348
rect 19392 30336 19398 30388
rect 1946 30308 1952 30320
rect 1596 30280 1952 30308
rect 1596 30249 1624 30280
rect 1946 30268 1952 30280
rect 2004 30268 2010 30320
rect 2314 30268 2320 30320
rect 2372 30268 2378 30320
rect 5534 30268 5540 30320
rect 5592 30268 5598 30320
rect 8018 30308 8024 30320
rect 6748 30280 8024 30308
rect 1581 30243 1639 30249
rect 1581 30209 1593 30243
rect 1627 30209 1639 30243
rect 1581 30203 1639 30209
rect 4154 30200 4160 30252
rect 4212 30240 4218 30252
rect 4249 30243 4307 30249
rect 4249 30240 4261 30243
rect 4212 30212 4261 30240
rect 4212 30200 4218 30212
rect 4249 30209 4261 30212
rect 4295 30209 4307 30243
rect 6546 30240 6552 30252
rect 6507 30212 6552 30240
rect 4249 30203 4307 30209
rect 6546 30200 6552 30212
rect 6604 30200 6610 30252
rect 1857 30175 1915 30181
rect 1857 30141 1869 30175
rect 1903 30172 1915 30175
rect 1903 30144 3096 30172
rect 1903 30141 1915 30144
rect 1857 30135 1915 30141
rect 3068 30104 3096 30144
rect 3142 30132 3148 30184
rect 3200 30172 3206 30184
rect 4525 30175 4583 30181
rect 4525 30172 4537 30175
rect 3200 30144 4537 30172
rect 3200 30132 3206 30144
rect 4525 30141 4537 30144
rect 4571 30172 4583 30175
rect 5902 30172 5908 30184
rect 4571 30144 5908 30172
rect 4571 30141 4583 30144
rect 4525 30135 4583 30141
rect 5902 30132 5908 30144
rect 5960 30132 5966 30184
rect 5997 30175 6055 30181
rect 5997 30141 6009 30175
rect 6043 30172 6055 30175
rect 6748 30172 6776 30280
rect 8018 30268 8024 30280
rect 8076 30268 8082 30320
rect 8312 30308 8340 30336
rect 13449 30311 13507 30317
rect 8312 30280 8418 30308
rect 12820 30280 13400 30308
rect 10134 30200 10140 30252
rect 10192 30240 10198 30252
rect 10321 30243 10379 30249
rect 10321 30240 10333 30243
rect 10192 30212 10333 30240
rect 10192 30200 10198 30212
rect 10321 30209 10333 30212
rect 10367 30209 10379 30243
rect 12158 30240 12164 30252
rect 12119 30212 12164 30240
rect 10321 30203 10379 30209
rect 12158 30200 12164 30212
rect 12216 30240 12222 30252
rect 12820 30249 12848 30280
rect 13372 30249 13400 30280
rect 13449 30277 13461 30311
rect 13495 30308 13507 30311
rect 15473 30311 15531 30317
rect 15473 30308 15485 30311
rect 13495 30280 15485 30308
rect 13495 30277 13507 30280
rect 13449 30271 13507 30277
rect 15473 30277 15485 30280
rect 15519 30277 15531 30311
rect 15473 30271 15531 30277
rect 12805 30243 12863 30249
rect 12805 30240 12817 30243
rect 12216 30212 12817 30240
rect 12216 30200 12222 30212
rect 12805 30209 12817 30212
rect 12851 30209 12863 30243
rect 12805 30203 12863 30209
rect 13357 30243 13415 30249
rect 13357 30209 13369 30243
rect 13403 30209 13415 30243
rect 13357 30203 13415 30209
rect 13906 30200 13912 30252
rect 13964 30240 13970 30252
rect 14090 30240 14096 30252
rect 13964 30212 14096 30240
rect 13964 30200 13970 30212
rect 14090 30200 14096 30212
rect 14148 30240 14154 30252
rect 14185 30243 14243 30249
rect 14185 30240 14197 30243
rect 14148 30212 14197 30240
rect 14148 30200 14154 30212
rect 14185 30209 14197 30212
rect 14231 30209 14243 30243
rect 14185 30203 14243 30209
rect 14274 30200 14280 30252
rect 14332 30240 14338 30252
rect 14829 30243 14887 30249
rect 14829 30240 14841 30243
rect 14332 30212 14841 30240
rect 14332 30200 14338 30212
rect 14829 30209 14841 30212
rect 14875 30240 14887 30243
rect 15102 30240 15108 30252
rect 14875 30212 15108 30240
rect 14875 30209 14887 30212
rect 14829 30203 14887 30209
rect 15102 30200 15108 30212
rect 15160 30200 15166 30252
rect 35894 30200 35900 30252
rect 35952 30240 35958 30252
rect 36081 30243 36139 30249
rect 36081 30240 36093 30243
rect 35952 30212 36093 30240
rect 35952 30200 35958 30212
rect 36081 30209 36093 30212
rect 36127 30209 36139 30243
rect 36081 30203 36139 30209
rect 6043 30144 6776 30172
rect 6043 30141 6055 30144
rect 5997 30135 6055 30141
rect 6822 30132 6828 30184
rect 6880 30172 6886 30184
rect 7653 30175 7711 30181
rect 6880 30144 7604 30172
rect 6880 30132 6886 30144
rect 3694 30104 3700 30116
rect 3068 30076 3700 30104
rect 3694 30064 3700 30076
rect 3752 30064 3758 30116
rect 7374 30104 7380 30116
rect 5552 30076 7380 30104
rect 3234 29996 3240 30048
rect 3292 30036 3298 30048
rect 5552 30036 5580 30076
rect 7374 30064 7380 30076
rect 7432 30064 7438 30116
rect 7576 30104 7604 30144
rect 7653 30141 7665 30175
rect 7699 30141 7711 30175
rect 7926 30172 7932 30184
rect 7887 30144 7932 30172
rect 7653 30135 7711 30141
rect 7668 30104 7696 30135
rect 7926 30132 7932 30144
rect 7984 30132 7990 30184
rect 8018 30132 8024 30184
rect 8076 30172 8082 30184
rect 11054 30172 11060 30184
rect 8076 30144 11060 30172
rect 8076 30132 8082 30144
rect 11054 30132 11060 30144
rect 11112 30132 11118 30184
rect 11149 30175 11207 30181
rect 11149 30141 11161 30175
rect 11195 30172 11207 30175
rect 12986 30172 12992 30184
rect 11195 30144 12992 30172
rect 11195 30141 11207 30144
rect 11149 30135 11207 30141
rect 12986 30132 12992 30144
rect 13044 30132 13050 30184
rect 14366 30132 14372 30184
rect 14424 30172 14430 30184
rect 15381 30175 15439 30181
rect 15381 30172 15393 30175
rect 14424 30144 15393 30172
rect 14424 30132 14430 30144
rect 15381 30141 15393 30144
rect 15427 30141 15439 30175
rect 16022 30172 16028 30184
rect 15983 30144 16028 30172
rect 15381 30135 15439 30141
rect 16022 30132 16028 30144
rect 16080 30132 16086 30184
rect 36354 30172 36360 30184
rect 36315 30144 36360 30172
rect 36354 30132 36360 30144
rect 36412 30132 36418 30184
rect 7576 30076 7696 30104
rect 10413 30107 10471 30113
rect 10413 30073 10425 30107
rect 10459 30104 10471 30107
rect 13170 30104 13176 30116
rect 10459 30076 13176 30104
rect 10459 30073 10471 30076
rect 10413 30067 10471 30073
rect 13170 30064 13176 30076
rect 13228 30064 13234 30116
rect 3292 30008 5580 30036
rect 6641 30039 6699 30045
rect 3292 29996 3298 30008
rect 6641 30005 6653 30039
rect 6687 30036 6699 30039
rect 8570 30036 8576 30048
rect 6687 30008 8576 30036
rect 6687 30005 6699 30008
rect 6641 29999 6699 30005
rect 8570 29996 8576 30008
rect 8628 29996 8634 30048
rect 9401 30039 9459 30045
rect 9401 30005 9413 30039
rect 9447 30036 9459 30039
rect 9766 30036 9772 30048
rect 9447 30008 9772 30036
rect 9447 30005 9459 30008
rect 9401 29999 9459 30005
rect 9766 29996 9772 30008
rect 9824 30036 9830 30048
rect 10502 30036 10508 30048
rect 9824 30008 10508 30036
rect 9824 29996 9830 30008
rect 10502 29996 10508 30008
rect 10560 29996 10566 30048
rect 11974 29996 11980 30048
rect 12032 30036 12038 30048
rect 12069 30039 12127 30045
rect 12069 30036 12081 30039
rect 12032 30008 12081 30036
rect 12032 29996 12038 30008
rect 12069 30005 12081 30008
rect 12115 30005 12127 30039
rect 12069 29999 12127 30005
rect 12434 29996 12440 30048
rect 12492 30036 12498 30048
rect 12713 30039 12771 30045
rect 12713 30036 12725 30039
rect 12492 30008 12725 30036
rect 12492 29996 12498 30008
rect 12713 30005 12725 30008
rect 12759 30005 12771 30039
rect 12713 29999 12771 30005
rect 12894 29996 12900 30048
rect 12952 30036 12958 30048
rect 13722 30036 13728 30048
rect 12952 30008 13728 30036
rect 12952 29996 12958 30008
rect 13722 29996 13728 30008
rect 13780 29996 13786 30048
rect 14090 30036 14096 30048
rect 14051 30008 14096 30036
rect 14090 29996 14096 30008
rect 14148 29996 14154 30048
rect 14737 30039 14795 30045
rect 14737 30005 14749 30039
rect 14783 30036 14795 30039
rect 15010 30036 15016 30048
rect 14783 30008 15016 30036
rect 14783 30005 14795 30008
rect 14737 29999 14795 30005
rect 15010 29996 15016 30008
rect 15068 29996 15074 30048
rect 15102 29996 15108 30048
rect 15160 30036 15166 30048
rect 16945 30039 17003 30045
rect 16945 30036 16957 30039
rect 15160 30008 16957 30036
rect 15160 29996 15166 30008
rect 16945 30005 16957 30008
rect 16991 30036 17003 30039
rect 25866 30036 25872 30048
rect 16991 30008 25872 30036
rect 16991 30005 17003 30008
rect 16945 29999 17003 30005
rect 25866 29996 25872 30008
rect 25924 29996 25930 30048
rect 1104 29946 36892 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 36892 29946
rect 1104 29872 36892 29894
rect 1670 29832 1676 29844
rect 1631 29804 1676 29832
rect 1670 29792 1676 29804
rect 1728 29792 1734 29844
rect 2314 29832 2320 29844
rect 2275 29804 2320 29832
rect 2314 29792 2320 29804
rect 2372 29792 2378 29844
rect 3970 29792 3976 29844
rect 4028 29832 4034 29844
rect 4065 29835 4123 29841
rect 4065 29832 4077 29835
rect 4028 29804 4077 29832
rect 4028 29792 4034 29804
rect 4065 29801 4077 29804
rect 4111 29801 4123 29835
rect 4065 29795 4123 29801
rect 4154 29792 4160 29844
rect 4212 29832 4218 29844
rect 5261 29835 5319 29841
rect 5261 29832 5273 29835
rect 4212 29804 5273 29832
rect 4212 29792 4218 29804
rect 5261 29801 5273 29804
rect 5307 29832 5319 29835
rect 5810 29832 5816 29844
rect 5307 29804 5816 29832
rect 5307 29801 5319 29804
rect 5261 29795 5319 29801
rect 5810 29792 5816 29804
rect 5868 29792 5874 29844
rect 5902 29792 5908 29844
rect 5960 29832 5966 29844
rect 8846 29832 8852 29844
rect 5960 29804 8852 29832
rect 5960 29792 5966 29804
rect 8846 29792 8852 29804
rect 8904 29792 8910 29844
rect 9125 29835 9183 29841
rect 9125 29801 9137 29835
rect 9171 29832 9183 29835
rect 9490 29832 9496 29844
rect 9171 29804 9496 29832
rect 9171 29801 9183 29804
rect 9125 29795 9183 29801
rect 9490 29792 9496 29804
rect 9548 29792 9554 29844
rect 10594 29832 10600 29844
rect 9600 29804 10600 29832
rect 3602 29724 3608 29776
rect 3660 29764 3666 29776
rect 4709 29767 4767 29773
rect 4709 29764 4721 29767
rect 3660 29736 4721 29764
rect 3660 29724 3666 29736
rect 4709 29733 4721 29736
rect 4755 29733 4767 29767
rect 4709 29727 4767 29733
rect 6104 29736 6960 29764
rect 2958 29696 2964 29708
rect 2240 29668 2964 29696
rect 2240 29637 2268 29668
rect 2958 29656 2964 29668
rect 3016 29656 3022 29708
rect 4614 29696 4620 29708
rect 3988 29668 4620 29696
rect 1765 29631 1823 29637
rect 1765 29597 1777 29631
rect 1811 29597 1823 29631
rect 1765 29591 1823 29597
rect 2225 29631 2283 29637
rect 2225 29597 2237 29631
rect 2271 29597 2283 29631
rect 2225 29591 2283 29597
rect 1780 29492 1808 29591
rect 2406 29588 2412 29640
rect 2464 29628 2470 29640
rect 2869 29631 2927 29637
rect 2869 29628 2881 29631
rect 2464 29600 2881 29628
rect 2464 29588 2470 29600
rect 2869 29597 2881 29600
rect 2915 29628 2927 29631
rect 3988 29628 4016 29668
rect 4614 29656 4620 29668
rect 4672 29696 4678 29708
rect 4672 29668 4844 29696
rect 4672 29656 4678 29668
rect 2915 29600 4016 29628
rect 2915 29597 2927 29600
rect 2869 29591 2927 29597
rect 4154 29588 4160 29640
rect 4212 29628 4218 29640
rect 4706 29628 4712 29640
rect 4212 29600 4712 29628
rect 4212 29588 4218 29600
rect 4706 29588 4712 29600
rect 4764 29588 4770 29640
rect 4816 29637 4844 29668
rect 4801 29631 4859 29637
rect 4801 29597 4813 29631
rect 4847 29597 4859 29631
rect 4801 29591 4859 29597
rect 5258 29588 5264 29640
rect 5316 29628 5322 29640
rect 5813 29631 5871 29637
rect 5813 29628 5825 29631
rect 5316 29600 5825 29628
rect 5316 29588 5322 29600
rect 5813 29597 5825 29600
rect 5859 29597 5871 29631
rect 5813 29591 5871 29597
rect 2961 29563 3019 29569
rect 2961 29529 2973 29563
rect 3007 29560 3019 29563
rect 6104 29560 6132 29736
rect 6546 29656 6552 29708
rect 6604 29696 6610 29708
rect 6822 29696 6828 29708
rect 6604 29668 6828 29696
rect 6604 29656 6610 29668
rect 6822 29656 6828 29668
rect 6880 29656 6886 29708
rect 6932 29696 6960 29736
rect 8110 29724 8116 29776
rect 8168 29764 8174 29776
rect 8573 29767 8631 29773
rect 8168 29736 8432 29764
rect 8168 29724 8174 29736
rect 8404 29696 8432 29736
rect 8573 29733 8585 29767
rect 8619 29764 8631 29767
rect 9600 29764 9628 29804
rect 10594 29792 10600 29804
rect 10652 29792 10658 29844
rect 11698 29792 11704 29844
rect 11756 29832 11762 29844
rect 12342 29832 12348 29844
rect 11756 29804 12348 29832
rect 11756 29792 11762 29804
rect 12342 29792 12348 29804
rect 12400 29832 12406 29844
rect 36354 29832 36360 29844
rect 12400 29804 13032 29832
rect 36315 29804 36360 29832
rect 12400 29792 12406 29804
rect 12158 29764 12164 29776
rect 8619 29736 9628 29764
rect 10796 29736 12164 29764
rect 8619 29733 8631 29736
rect 8573 29727 8631 29733
rect 10796 29696 10824 29736
rect 12158 29724 12164 29736
rect 12216 29724 12222 29776
rect 12802 29764 12808 29776
rect 12360 29736 12808 29764
rect 12360 29705 12388 29736
rect 12802 29724 12808 29736
rect 12860 29724 12866 29776
rect 6932 29668 8340 29696
rect 8404 29668 10824 29696
rect 12345 29699 12403 29705
rect 8312 29628 8340 29668
rect 12345 29665 12357 29699
rect 12391 29665 12403 29699
rect 13004 29696 13032 29804
rect 36354 29792 36360 29804
rect 36412 29792 36418 29844
rect 14274 29724 14280 29776
rect 14332 29764 14338 29776
rect 14332 29736 14688 29764
rect 14332 29724 14338 29736
rect 13265 29699 13323 29705
rect 13265 29696 13277 29699
rect 13004 29668 13277 29696
rect 12345 29659 12403 29665
rect 13265 29665 13277 29668
rect 13311 29665 13323 29699
rect 13265 29659 13323 29665
rect 13630 29656 13636 29708
rect 13688 29696 13694 29708
rect 14660 29705 14688 29736
rect 14369 29699 14427 29705
rect 14369 29696 14381 29699
rect 13688 29668 14381 29696
rect 13688 29656 13694 29668
rect 14369 29665 14381 29668
rect 14415 29665 14427 29699
rect 14369 29659 14427 29665
rect 14645 29699 14703 29705
rect 14645 29665 14657 29699
rect 14691 29665 14703 29699
rect 16206 29696 16212 29708
rect 16167 29668 16212 29696
rect 14645 29659 14703 29665
rect 16206 29656 16212 29668
rect 16264 29656 16270 29708
rect 10884 29631 10942 29637
rect 8312 29600 8432 29628
rect 3007 29532 6132 29560
rect 3007 29529 3019 29532
rect 2961 29523 3019 29529
rect 6270 29520 6276 29572
rect 6328 29560 6334 29572
rect 6730 29560 6736 29572
rect 6328 29532 6736 29560
rect 6328 29520 6334 29532
rect 6730 29520 6736 29532
rect 6788 29560 6794 29572
rect 7101 29563 7159 29569
rect 7101 29560 7113 29563
rect 6788 29532 7113 29560
rect 6788 29520 6794 29532
rect 7101 29529 7113 29532
rect 7147 29560 7159 29563
rect 7374 29560 7380 29572
rect 7147 29532 7380 29560
rect 7147 29529 7159 29532
rect 7101 29523 7159 29529
rect 7374 29520 7380 29532
rect 7432 29520 7438 29572
rect 7558 29520 7564 29572
rect 7616 29520 7622 29572
rect 8404 29560 8432 29600
rect 10884 29597 10896 29631
rect 10930 29628 10942 29631
rect 11146 29628 11152 29640
rect 10930 29600 11152 29628
rect 10930 29597 10942 29600
rect 10884 29591 10942 29597
rect 11146 29588 11152 29600
rect 11204 29588 11210 29640
rect 12526 29588 12532 29640
rect 12584 29628 12590 29640
rect 12802 29628 12808 29640
rect 12584 29600 12808 29628
rect 12584 29588 12590 29600
rect 12802 29588 12808 29600
rect 12860 29588 12866 29640
rect 10597 29563 10655 29569
rect 8404 29532 9430 29560
rect 10597 29529 10609 29563
rect 10643 29560 10655 29563
rect 11054 29560 11060 29572
rect 10643 29532 11060 29560
rect 10643 29529 10655 29532
rect 10597 29523 10655 29529
rect 11054 29520 11060 29532
rect 11112 29520 11118 29572
rect 11425 29563 11483 29569
rect 11425 29529 11437 29563
rect 11471 29529 11483 29563
rect 11425 29523 11483 29529
rect 4154 29492 4160 29504
rect 1780 29464 4160 29492
rect 4154 29452 4160 29464
rect 4212 29452 4218 29504
rect 5905 29495 5963 29501
rect 5905 29461 5917 29495
rect 5951 29492 5963 29495
rect 8478 29492 8484 29504
rect 5951 29464 8484 29492
rect 5951 29461 5963 29464
rect 5905 29455 5963 29461
rect 8478 29452 8484 29464
rect 8536 29452 8542 29504
rect 11440 29492 11468 29523
rect 11514 29520 11520 29572
rect 11572 29560 11578 29572
rect 12986 29560 12992 29572
rect 11572 29532 11617 29560
rect 12947 29532 12992 29560
rect 11572 29520 11578 29532
rect 12986 29520 12992 29532
rect 13044 29520 13050 29572
rect 13081 29563 13139 29569
rect 13081 29529 13093 29563
rect 13127 29560 13139 29563
rect 13170 29560 13176 29572
rect 13127 29532 13176 29560
rect 13127 29529 13139 29532
rect 13081 29523 13139 29529
rect 13170 29520 13176 29532
rect 13228 29520 13234 29572
rect 14461 29563 14519 29569
rect 14461 29529 14473 29563
rect 14507 29529 14519 29563
rect 16390 29560 16396 29572
rect 16351 29532 16396 29560
rect 14461 29523 14519 29529
rect 12894 29492 12900 29504
rect 11440 29464 12900 29492
rect 12894 29452 12900 29464
rect 12952 29452 12958 29504
rect 14476 29492 14504 29523
rect 16390 29520 16396 29532
rect 16448 29520 16454 29572
rect 16485 29563 16543 29569
rect 16485 29529 16497 29563
rect 16531 29560 16543 29563
rect 16850 29560 16856 29572
rect 16531 29532 16856 29560
rect 16531 29529 16543 29532
rect 16485 29523 16543 29529
rect 16850 29520 16856 29532
rect 16908 29520 16914 29572
rect 15562 29492 15568 29504
rect 14476 29464 15568 29492
rect 15562 29452 15568 29464
rect 15620 29452 15626 29504
rect 17221 29495 17279 29501
rect 17221 29461 17233 29495
rect 17267 29492 17279 29495
rect 17494 29492 17500 29504
rect 17267 29464 17500 29492
rect 17267 29461 17279 29464
rect 17221 29455 17279 29461
rect 17494 29452 17500 29464
rect 17552 29452 17558 29504
rect 1104 29402 36892 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 36892 29402
rect 1104 29328 36892 29350
rect 2961 29291 3019 29297
rect 1872 29260 2774 29288
rect 1872 29161 1900 29260
rect 1857 29155 1915 29161
rect 1857 29121 1869 29155
rect 1903 29121 1915 29155
rect 1857 29115 1915 29121
rect 1578 29084 1584 29096
rect 1539 29056 1584 29084
rect 1578 29044 1584 29056
rect 1636 29044 1642 29096
rect 2746 29084 2774 29260
rect 2961 29257 2973 29291
rect 3007 29288 3019 29291
rect 3142 29288 3148 29300
rect 3007 29260 3148 29288
rect 3007 29257 3019 29260
rect 2961 29251 3019 29257
rect 3142 29248 3148 29260
rect 3200 29248 3206 29300
rect 5445 29291 5503 29297
rect 5445 29257 5457 29291
rect 5491 29288 5503 29291
rect 5810 29288 5816 29300
rect 5491 29260 5816 29288
rect 5491 29257 5503 29260
rect 5445 29251 5503 29257
rect 3050 29180 3056 29232
rect 3108 29220 3114 29232
rect 3108 29192 3266 29220
rect 3108 29180 3114 29192
rect 4709 29155 4767 29161
rect 4709 29121 4721 29155
rect 4755 29152 4767 29155
rect 5460 29152 5488 29251
rect 5810 29248 5816 29260
rect 5868 29248 5874 29300
rect 5997 29291 6055 29297
rect 5997 29257 6009 29291
rect 6043 29288 6055 29291
rect 6270 29288 6276 29300
rect 6043 29260 6276 29288
rect 6043 29257 6055 29260
rect 5997 29251 6055 29257
rect 6270 29248 6276 29260
rect 6328 29248 6334 29300
rect 8849 29291 8907 29297
rect 6840 29260 8800 29288
rect 6454 29180 6460 29232
rect 6512 29220 6518 29232
rect 6840 29229 6868 29260
rect 6825 29223 6883 29229
rect 6825 29220 6837 29223
rect 6512 29192 6837 29220
rect 6512 29180 6518 29192
rect 6825 29189 6837 29192
rect 6871 29189 6883 29223
rect 6825 29183 6883 29189
rect 7282 29180 7288 29232
rect 7340 29180 7346 29232
rect 6546 29152 6552 29164
rect 4755 29124 6552 29152
rect 4755 29121 4767 29124
rect 4709 29115 4767 29121
rect 6546 29112 6552 29124
rect 6604 29112 6610 29164
rect 8772 29161 8800 29260
rect 8849 29257 8861 29291
rect 8895 29257 8907 29291
rect 8849 29251 8907 29257
rect 9493 29291 9551 29297
rect 9493 29257 9505 29291
rect 9539 29288 9551 29291
rect 11514 29288 11520 29300
rect 9539 29260 11520 29288
rect 9539 29257 9551 29260
rect 9493 29251 9551 29257
rect 8864 29220 8892 29251
rect 11514 29248 11520 29260
rect 11572 29248 11578 29300
rect 12158 29248 12164 29300
rect 12216 29288 12222 29300
rect 13906 29288 13912 29300
rect 12216 29260 13912 29288
rect 12216 29248 12222 29260
rect 13906 29248 13912 29260
rect 13964 29248 13970 29300
rect 14550 29248 14556 29300
rect 14608 29288 14614 29300
rect 17126 29288 17132 29300
rect 14608 29260 17132 29288
rect 14608 29248 14614 29260
rect 9674 29220 9680 29232
rect 8864 29192 9680 29220
rect 9674 29180 9680 29192
rect 9732 29180 9738 29232
rect 9950 29180 9956 29232
rect 10008 29220 10014 29232
rect 10229 29223 10287 29229
rect 10229 29220 10241 29223
rect 10008 29192 10241 29220
rect 10008 29180 10014 29192
rect 10229 29189 10241 29192
rect 10275 29189 10287 29223
rect 10229 29183 10287 29189
rect 10781 29223 10839 29229
rect 10781 29189 10793 29223
rect 10827 29220 10839 29223
rect 11698 29220 11704 29232
rect 10827 29192 11704 29220
rect 10827 29189 10839 29192
rect 10781 29183 10839 29189
rect 11698 29180 11704 29192
rect 11756 29180 11762 29232
rect 12434 29180 12440 29232
rect 12492 29220 12498 29232
rect 12492 29192 12537 29220
rect 12492 29180 12498 29192
rect 12710 29180 12716 29232
rect 12768 29220 12774 29232
rect 13633 29223 13691 29229
rect 13633 29220 13645 29223
rect 12768 29192 13645 29220
rect 12768 29180 12774 29192
rect 13633 29189 13645 29192
rect 13679 29189 13691 29223
rect 13633 29183 13691 29189
rect 13998 29180 14004 29232
rect 14056 29220 14062 29232
rect 16132 29229 16160 29260
rect 17126 29248 17132 29260
rect 17184 29248 17190 29300
rect 18138 29288 18144 29300
rect 17420 29260 18144 29288
rect 15197 29223 15255 29229
rect 15197 29220 15209 29223
rect 14056 29192 15209 29220
rect 14056 29180 14062 29192
rect 15197 29189 15209 29192
rect 15243 29189 15255 29223
rect 15197 29183 15255 29189
rect 16117 29223 16175 29229
rect 16117 29189 16129 29223
rect 16163 29189 16175 29223
rect 16117 29183 16175 29189
rect 16206 29180 16212 29232
rect 16264 29220 16270 29232
rect 17420 29229 17448 29260
rect 18138 29248 18144 29260
rect 18196 29248 18202 29300
rect 16853 29223 16911 29229
rect 16853 29220 16865 29223
rect 16264 29192 16865 29220
rect 16264 29180 16270 29192
rect 16853 29189 16865 29192
rect 16899 29189 16911 29223
rect 16853 29183 16911 29189
rect 17405 29223 17463 29229
rect 17405 29189 17417 29223
rect 17451 29189 17463 29223
rect 17405 29183 17463 29189
rect 17494 29180 17500 29232
rect 17552 29220 17558 29232
rect 17552 29192 17597 29220
rect 17552 29180 17558 29192
rect 8757 29155 8815 29161
rect 8757 29121 8769 29155
rect 8803 29121 8815 29155
rect 8757 29115 8815 29121
rect 8846 29112 8852 29164
rect 8904 29152 8910 29164
rect 9401 29155 9459 29161
rect 9401 29152 9413 29155
rect 8904 29124 9413 29152
rect 8904 29112 8910 29124
rect 9401 29121 9413 29124
rect 9447 29121 9459 29155
rect 18046 29152 18052 29164
rect 18007 29124 18052 29152
rect 9401 29115 9459 29121
rect 18046 29112 18052 29124
rect 18104 29112 18110 29164
rect 2746 29056 8156 29084
rect 5166 29016 5172 29028
rect 4724 28988 5172 29016
rect 4451 28951 4509 28957
rect 4451 28917 4463 28951
rect 4497 28948 4509 28951
rect 4724 28948 4752 28988
rect 5166 28976 5172 28988
rect 5224 28976 5230 29028
rect 4497 28920 4752 28948
rect 4497 28917 4509 28920
rect 4451 28911 4509 28917
rect 4798 28908 4804 28960
rect 4856 28948 4862 28960
rect 5350 28948 5356 28960
rect 4856 28920 5356 28948
rect 4856 28908 4862 28920
rect 5350 28908 5356 28920
rect 5408 28948 5414 28960
rect 7374 28948 7380 28960
rect 5408 28920 7380 28948
rect 5408 28908 5414 28920
rect 7374 28908 7380 28920
rect 7432 28908 7438 28960
rect 8128 28948 8156 29056
rect 8478 29044 8484 29096
rect 8536 29084 8542 29096
rect 10137 29087 10195 29093
rect 10137 29084 10149 29087
rect 8536 29056 10149 29084
rect 8536 29044 8542 29056
rect 10137 29053 10149 29056
rect 10183 29053 10195 29087
rect 10137 29047 10195 29053
rect 10778 29044 10784 29096
rect 10836 29084 10842 29096
rect 12345 29087 12403 29093
rect 12345 29084 12357 29087
rect 10836 29056 12357 29084
rect 10836 29044 10842 29056
rect 12345 29053 12357 29056
rect 12391 29053 12403 29087
rect 12345 29047 12403 29053
rect 12989 29087 13047 29093
rect 12989 29053 13001 29087
rect 13035 29084 13047 29087
rect 13541 29087 13599 29093
rect 13035 29056 13492 29084
rect 13035 29053 13047 29056
rect 12989 29047 13047 29053
rect 8294 29016 8300 29028
rect 8207 28988 8300 29016
rect 8294 28976 8300 28988
rect 8352 29016 8358 29028
rect 9122 29016 9128 29028
rect 8352 28988 9128 29016
rect 8352 28976 8358 28988
rect 9122 28976 9128 28988
rect 9180 28976 9186 29028
rect 10226 29016 10232 29028
rect 9232 28988 10232 29016
rect 9232 28948 9260 28988
rect 10226 28976 10232 28988
rect 10284 28976 10290 29028
rect 10318 28976 10324 29028
rect 10376 29016 10382 29028
rect 13354 29016 13360 29028
rect 10376 28988 13360 29016
rect 10376 28976 10382 28988
rect 13354 28976 13360 28988
rect 13412 28976 13418 29028
rect 13464 29016 13492 29056
rect 13541 29053 13553 29087
rect 13587 29072 13599 29087
rect 13630 29072 13636 29096
rect 13587 29053 13636 29072
rect 13541 29047 13636 29053
rect 13556 29044 13636 29047
rect 13688 29044 13694 29096
rect 14550 29044 14556 29096
rect 14608 29084 14614 29096
rect 15105 29087 15163 29093
rect 14608 29056 14653 29084
rect 14608 29044 14614 29056
rect 15105 29053 15117 29087
rect 15151 29053 15163 29087
rect 15105 29047 15163 29053
rect 15120 29016 15148 29047
rect 16390 29044 16396 29096
rect 16448 29084 16454 29096
rect 18141 29087 18199 29093
rect 18141 29084 18153 29087
rect 16448 29056 18153 29084
rect 16448 29044 16454 29056
rect 18141 29053 18153 29056
rect 18187 29053 18199 29087
rect 18141 29047 18199 29053
rect 16298 29016 16304 29028
rect 13464 28988 16304 29016
rect 16298 28976 16304 28988
rect 16356 28976 16362 29028
rect 8128 28920 9260 28948
rect 12526 28908 12532 28960
rect 12584 28948 12590 28960
rect 13630 28948 13636 28960
rect 12584 28920 13636 28948
rect 12584 28908 12590 28920
rect 13630 28908 13636 28920
rect 13688 28908 13694 28960
rect 18046 28908 18052 28960
rect 18104 28948 18110 28960
rect 18693 28951 18751 28957
rect 18693 28948 18705 28951
rect 18104 28920 18705 28948
rect 18104 28908 18110 28920
rect 18693 28917 18705 28920
rect 18739 28917 18751 28951
rect 18693 28911 18751 28917
rect 1104 28858 36892 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 36892 28858
rect 1104 28784 36892 28806
rect 4062 28744 4068 28756
rect 4023 28716 4068 28744
rect 4062 28704 4068 28716
rect 4120 28744 4126 28756
rect 4709 28747 4767 28753
rect 4709 28744 4721 28747
rect 4120 28716 4721 28744
rect 4120 28704 4126 28716
rect 4709 28713 4721 28716
rect 4755 28713 4767 28747
rect 5810 28744 5816 28756
rect 5771 28716 5816 28744
rect 4709 28707 4767 28713
rect 5810 28704 5816 28716
rect 5868 28704 5874 28756
rect 7282 28744 7288 28756
rect 5920 28716 7288 28744
rect 2317 28679 2375 28685
rect 2317 28645 2329 28679
rect 2363 28676 2375 28679
rect 5920 28676 5948 28716
rect 7282 28704 7288 28716
rect 7340 28704 7346 28756
rect 7374 28704 7380 28756
rect 7432 28744 7438 28756
rect 7432 28716 9352 28744
rect 7432 28704 7438 28716
rect 2363 28648 5948 28676
rect 2363 28645 2375 28648
rect 2317 28639 2375 28645
rect 2498 28568 2504 28620
rect 2556 28608 2562 28620
rect 4982 28608 4988 28620
rect 2556 28580 4988 28608
rect 2556 28568 2562 28580
rect 4982 28568 4988 28580
rect 5040 28568 5046 28620
rect 6546 28568 6552 28620
rect 6604 28608 6610 28620
rect 8113 28611 8171 28617
rect 8113 28608 8125 28611
rect 6604 28580 8125 28608
rect 6604 28568 6610 28580
rect 8113 28577 8125 28580
rect 8159 28577 8171 28611
rect 8113 28571 8171 28577
rect 1765 28543 1823 28549
rect 1765 28509 1777 28543
rect 1811 28509 1823 28543
rect 1765 28503 1823 28509
rect 2225 28543 2283 28549
rect 2225 28509 2237 28543
rect 2271 28540 2283 28543
rect 2866 28540 2872 28552
rect 2271 28512 2872 28540
rect 2271 28509 2283 28512
rect 2225 28503 2283 28509
rect 1780 28472 1808 28503
rect 2866 28500 2872 28512
rect 2924 28500 2930 28552
rect 9324 28549 9352 28716
rect 13354 28704 13360 28756
rect 13412 28744 13418 28756
rect 13814 28744 13820 28756
rect 13412 28716 13820 28744
rect 13412 28704 13418 28716
rect 13814 28704 13820 28716
rect 13872 28704 13878 28756
rect 14826 28704 14832 28756
rect 14884 28744 14890 28756
rect 18138 28744 18144 28756
rect 14884 28716 17080 28744
rect 18099 28716 18144 28744
rect 14884 28704 14890 28716
rect 15010 28676 15016 28688
rect 13740 28648 15016 28676
rect 13644 28623 13702 28629
rect 9401 28611 9459 28617
rect 9401 28577 9413 28611
rect 9447 28608 9459 28611
rect 10689 28611 10747 28617
rect 10689 28608 10701 28611
rect 9447 28580 10701 28608
rect 9447 28577 9459 28580
rect 9401 28571 9459 28577
rect 10689 28577 10701 28580
rect 10735 28608 10747 28611
rect 10778 28608 10784 28620
rect 10735 28580 10784 28608
rect 10735 28577 10747 28580
rect 10689 28571 10747 28577
rect 10778 28568 10784 28580
rect 10836 28568 10842 28620
rect 11606 28568 11612 28620
rect 11664 28608 11670 28620
rect 12342 28608 12348 28620
rect 11664 28580 12348 28608
rect 11664 28568 11670 28580
rect 12342 28568 12348 28580
rect 12400 28608 12406 28620
rect 12989 28611 13047 28617
rect 12989 28608 13001 28611
rect 12400 28580 13001 28608
rect 12400 28568 12406 28580
rect 12989 28577 13001 28580
rect 13035 28577 13047 28611
rect 13644 28589 13656 28623
rect 13690 28620 13702 28623
rect 13740 28620 13768 28648
rect 15010 28636 15016 28648
rect 15068 28636 15074 28688
rect 13690 28592 13768 28620
rect 15286 28608 15292 28620
rect 13690 28589 13702 28592
rect 13644 28583 13702 28589
rect 15247 28580 15292 28608
rect 12989 28571 13047 28577
rect 15286 28568 15292 28580
rect 15344 28568 15350 28620
rect 16022 28568 16028 28620
rect 16080 28608 16086 28620
rect 16209 28611 16267 28617
rect 16209 28608 16221 28611
rect 16080 28580 16221 28608
rect 16080 28568 16086 28580
rect 16209 28577 16221 28580
rect 16255 28608 16267 28611
rect 16482 28608 16488 28620
rect 16255 28580 16488 28608
rect 16255 28577 16267 28580
rect 16209 28571 16267 28577
rect 16482 28568 16488 28580
rect 16540 28568 16546 28620
rect 9309 28543 9367 28549
rect 9309 28509 9321 28543
rect 9355 28509 9367 28543
rect 9309 28503 9367 28509
rect 9953 28543 10011 28549
rect 9953 28509 9965 28543
rect 9999 28509 10011 28543
rect 9953 28503 10011 28509
rect 14277 28543 14335 28549
rect 14277 28509 14289 28543
rect 14323 28540 14335 28543
rect 14642 28540 14648 28552
rect 14323 28512 14648 28540
rect 14323 28509 14335 28512
rect 14277 28503 14335 28509
rect 2961 28475 3019 28481
rect 1780 28444 2774 28472
rect 1670 28404 1676 28416
rect 1631 28376 1676 28404
rect 1670 28364 1676 28376
rect 1728 28364 1734 28416
rect 2746 28404 2774 28444
rect 2961 28441 2973 28475
rect 3007 28472 3019 28475
rect 7837 28475 7895 28481
rect 3007 28444 6670 28472
rect 3007 28441 3019 28444
rect 2961 28435 3019 28441
rect 7837 28441 7849 28475
rect 7883 28472 7895 28475
rect 8294 28472 8300 28484
rect 7883 28444 8300 28472
rect 7883 28441 7895 28444
rect 7837 28435 7895 28441
rect 8294 28432 8300 28444
rect 8352 28432 8358 28484
rect 8386 28432 8392 28484
rect 8444 28472 8450 28484
rect 9968 28472 9996 28503
rect 14642 28500 14648 28512
rect 14700 28500 14706 28552
rect 17052 28540 17080 28716
rect 18138 28704 18144 28716
rect 18196 28704 18202 28756
rect 17405 28543 17463 28549
rect 17405 28540 17417 28543
rect 17052 28512 17417 28540
rect 17405 28509 17417 28512
rect 17451 28509 17463 28543
rect 17405 28503 17463 28509
rect 18046 28500 18052 28552
rect 18104 28540 18110 28552
rect 18233 28543 18291 28549
rect 18233 28540 18245 28543
rect 18104 28512 18245 28540
rect 18104 28500 18110 28512
rect 18233 28509 18245 28512
rect 18279 28509 18291 28543
rect 18233 28503 18291 28509
rect 30469 28543 30527 28549
rect 30469 28509 30481 28543
rect 30515 28540 30527 28543
rect 35986 28540 35992 28552
rect 30515 28512 35992 28540
rect 30515 28509 30527 28512
rect 30469 28503 30527 28509
rect 35986 28500 35992 28512
rect 36044 28500 36050 28552
rect 8444 28444 9996 28472
rect 10781 28475 10839 28481
rect 8444 28432 8450 28444
rect 10781 28441 10793 28475
rect 10827 28472 10839 28475
rect 11054 28472 11060 28484
rect 10827 28444 11060 28472
rect 10827 28441 10839 28444
rect 10781 28435 10839 28441
rect 11054 28432 11060 28444
rect 11112 28432 11118 28484
rect 11330 28472 11336 28484
rect 11291 28444 11336 28472
rect 11330 28432 11336 28444
rect 11388 28432 11394 28484
rect 11885 28475 11943 28481
rect 11885 28441 11897 28475
rect 11931 28441 11943 28475
rect 11885 28435 11943 28441
rect 2866 28404 2872 28416
rect 2746 28376 2872 28404
rect 2866 28364 2872 28376
rect 2924 28404 2930 28416
rect 3878 28404 3884 28416
rect 2924 28376 3884 28404
rect 2924 28364 2930 28376
rect 3878 28364 3884 28376
rect 3936 28364 3942 28416
rect 5258 28404 5264 28416
rect 5219 28376 5264 28404
rect 5258 28364 5264 28376
rect 5316 28364 5322 28416
rect 6365 28407 6423 28413
rect 6365 28373 6377 28407
rect 6411 28404 6423 28407
rect 7006 28404 7012 28416
rect 6411 28376 7012 28404
rect 6411 28373 6423 28376
rect 6365 28367 6423 28373
rect 7006 28364 7012 28376
rect 7064 28404 7070 28416
rect 7926 28404 7932 28416
rect 7064 28376 7932 28404
rect 7064 28364 7070 28376
rect 7926 28364 7932 28376
rect 7984 28364 7990 28416
rect 10045 28407 10103 28413
rect 10045 28373 10057 28407
rect 10091 28404 10103 28407
rect 11422 28404 11428 28416
rect 10091 28376 11428 28404
rect 10091 28373 10103 28376
rect 10045 28367 10103 28373
rect 11422 28364 11428 28376
rect 11480 28404 11486 28416
rect 11900 28404 11928 28435
rect 11974 28432 11980 28484
rect 12032 28472 12038 28484
rect 12526 28472 12532 28484
rect 12032 28444 12077 28472
rect 12487 28444 12532 28472
rect 12032 28432 12038 28444
rect 12526 28432 12532 28444
rect 12584 28432 12590 28484
rect 13541 28475 13599 28481
rect 13541 28441 13553 28475
rect 13587 28441 13599 28475
rect 15470 28472 15476 28484
rect 15431 28444 15476 28472
rect 13541 28435 13599 28441
rect 11480 28376 11928 28404
rect 13556 28404 13584 28435
rect 15470 28432 15476 28444
rect 15528 28432 15534 28484
rect 15562 28432 15568 28484
rect 15620 28472 15626 28484
rect 16761 28475 16819 28481
rect 15620 28444 15665 28472
rect 15620 28432 15626 28444
rect 16761 28441 16773 28475
rect 16807 28441 16819 28475
rect 16761 28435 16819 28441
rect 14090 28404 14096 28416
rect 13556 28376 14096 28404
rect 11480 28364 11486 28376
rect 14090 28364 14096 28376
rect 14148 28364 14154 28416
rect 14366 28404 14372 28416
rect 14327 28376 14372 28404
rect 14366 28364 14372 28376
rect 14424 28364 14430 28416
rect 16776 28404 16804 28435
rect 16850 28432 16856 28484
rect 16908 28472 16914 28484
rect 30377 28475 30435 28481
rect 30377 28472 30389 28475
rect 16908 28444 30389 28472
rect 16908 28432 16914 28444
rect 30377 28441 30389 28444
rect 30423 28441 30435 28475
rect 30377 28435 30435 28441
rect 17497 28407 17555 28413
rect 17497 28404 17509 28407
rect 16776 28376 17509 28404
rect 17497 28373 17509 28376
rect 17543 28373 17555 28407
rect 18690 28404 18696 28416
rect 18651 28376 18696 28404
rect 17497 28367 17555 28373
rect 18690 28364 18696 28376
rect 18748 28364 18754 28416
rect 1104 28314 36892 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 36892 28314
rect 1104 28240 36892 28262
rect 2961 28203 3019 28209
rect 2961 28169 2973 28203
rect 3007 28200 3019 28203
rect 3234 28200 3240 28212
rect 3007 28172 3240 28200
rect 3007 28169 3019 28172
rect 2961 28163 3019 28169
rect 3234 28160 3240 28172
rect 3292 28160 3298 28212
rect 3605 28203 3663 28209
rect 3605 28169 3617 28203
rect 3651 28200 3663 28203
rect 4062 28200 4068 28212
rect 3651 28172 4068 28200
rect 3651 28169 3663 28172
rect 3605 28163 3663 28169
rect 4062 28160 4068 28172
rect 4120 28160 4126 28212
rect 9306 28200 9312 28212
rect 4908 28172 9312 28200
rect 1670 28092 1676 28144
rect 1728 28132 1734 28144
rect 4908 28132 4936 28172
rect 9306 28160 9312 28172
rect 9364 28160 9370 28212
rect 11054 28200 11060 28212
rect 11015 28172 11060 28200
rect 11054 28160 11060 28172
rect 11112 28160 11118 28212
rect 11793 28203 11851 28209
rect 11793 28169 11805 28203
rect 11839 28200 11851 28203
rect 12250 28200 12256 28212
rect 11839 28172 12256 28200
rect 11839 28169 11851 28172
rect 11793 28163 11851 28169
rect 12250 28160 12256 28172
rect 12308 28160 12314 28212
rect 12345 28203 12403 28209
rect 12345 28169 12357 28203
rect 12391 28200 12403 28203
rect 15470 28200 15476 28212
rect 12391 28172 15476 28200
rect 12391 28169 12403 28172
rect 12345 28163 12403 28169
rect 15470 28160 15476 28172
rect 15528 28160 15534 28212
rect 18601 28203 18659 28209
rect 18601 28200 18613 28203
rect 15580 28172 18613 28200
rect 1728 28104 4936 28132
rect 1728 28092 1734 28104
rect 4982 28092 4988 28144
rect 5040 28132 5046 28144
rect 9490 28132 9496 28144
rect 5040 28104 7236 28132
rect 9451 28104 9496 28132
rect 5040 28092 5046 28104
rect 1765 28067 1823 28073
rect 1765 28033 1777 28067
rect 1811 28033 1823 28067
rect 1765 28027 1823 28033
rect 2225 28067 2283 28073
rect 2225 28033 2237 28067
rect 2271 28064 2283 28067
rect 2406 28064 2412 28076
rect 2271 28036 2412 28064
rect 2271 28033 2283 28036
rect 2225 28027 2283 28033
rect 1780 27928 1808 28027
rect 2406 28024 2412 28036
rect 2464 28024 2470 28076
rect 2866 28064 2872 28076
rect 2827 28036 2872 28064
rect 2866 28024 2872 28036
rect 2924 28024 2930 28076
rect 5074 28024 5080 28076
rect 5132 28064 5138 28076
rect 7208 28073 7236 28104
rect 9490 28092 9496 28104
rect 9548 28092 9554 28144
rect 12434 28092 12440 28144
rect 12492 28132 12498 28144
rect 13449 28135 13507 28141
rect 13449 28132 13461 28135
rect 12492 28104 13461 28132
rect 12492 28092 12498 28104
rect 13449 28101 13461 28104
rect 13495 28101 13507 28135
rect 13449 28095 13507 28101
rect 13538 28092 13544 28144
rect 13596 28132 13602 28144
rect 14921 28135 14979 28141
rect 13596 28104 13641 28132
rect 13596 28092 13602 28104
rect 14921 28101 14933 28135
rect 14967 28132 14979 28135
rect 15580 28132 15608 28172
rect 18601 28169 18613 28172
rect 18647 28169 18659 28203
rect 18601 28163 18659 28169
rect 15746 28132 15752 28144
rect 14967 28104 15608 28132
rect 15707 28104 15752 28132
rect 14967 28101 14979 28104
rect 14921 28095 14979 28101
rect 15746 28092 15752 28104
rect 15804 28092 15810 28144
rect 16298 28132 16304 28144
rect 16259 28104 16304 28132
rect 16298 28092 16304 28104
rect 16356 28092 16362 28144
rect 19705 28135 19763 28141
rect 19705 28132 19717 28135
rect 18064 28104 19717 28132
rect 18064 28076 18092 28104
rect 19705 28101 19717 28104
rect 19751 28101 19763 28135
rect 19705 28095 19763 28101
rect 6549 28067 6607 28073
rect 6549 28064 6561 28067
rect 5132 28036 6561 28064
rect 5132 28024 5138 28036
rect 6549 28033 6561 28036
rect 6595 28033 6607 28067
rect 6549 28027 6607 28033
rect 7193 28067 7251 28073
rect 7193 28033 7205 28067
rect 7239 28033 7251 28067
rect 7834 28064 7840 28076
rect 7795 28036 7840 28064
rect 7193 28027 7251 28033
rect 7834 28024 7840 28036
rect 7892 28024 7898 28076
rect 7926 28024 7932 28076
rect 7984 28064 7990 28076
rect 8665 28067 8723 28073
rect 8665 28064 8677 28067
rect 7984 28036 8677 28064
rect 7984 28024 7990 28036
rect 8665 28033 8677 28036
rect 8711 28033 8723 28067
rect 8665 28027 8723 28033
rect 10410 28024 10416 28076
rect 10468 28064 10474 28076
rect 11149 28067 11207 28073
rect 11149 28064 11161 28067
rect 10468 28036 11161 28064
rect 10468 28024 10474 28036
rect 11149 28033 11161 28036
rect 11195 28033 11207 28067
rect 11149 28027 11207 28033
rect 11238 28024 11244 28076
rect 11296 28064 11302 28076
rect 11882 28064 11888 28076
rect 11296 28036 11888 28064
rect 11296 28024 11302 28036
rect 11882 28024 11888 28036
rect 11940 28064 11946 28076
rect 12253 28067 12311 28073
rect 12253 28064 12265 28067
rect 11940 28036 12265 28064
rect 11940 28024 11946 28036
rect 12253 28033 12265 28036
rect 12299 28033 12311 28067
rect 18046 28064 18052 28076
rect 18007 28036 18052 28064
rect 12253 28027 12311 28033
rect 18046 28024 18052 28036
rect 18104 28024 18110 28076
rect 18690 28064 18696 28076
rect 18651 28036 18696 28064
rect 18690 28024 18696 28036
rect 18748 28024 18754 28076
rect 36081 28067 36139 28073
rect 36081 28033 36093 28067
rect 36127 28064 36139 28067
rect 36446 28064 36452 28076
rect 36127 28036 36452 28064
rect 36127 28033 36139 28036
rect 36081 28027 36139 28033
rect 36446 28024 36452 28036
rect 36504 28024 36510 28076
rect 2317 27999 2375 28005
rect 2317 27965 2329 27999
rect 2363 27996 2375 27999
rect 5534 27996 5540 28008
rect 2363 27968 5540 27996
rect 2363 27965 2375 27968
rect 2317 27959 2375 27965
rect 5534 27956 5540 27968
rect 5592 27956 5598 28008
rect 5810 27956 5816 28008
rect 5868 27996 5874 28008
rect 5905 27999 5963 28005
rect 5905 27996 5917 27999
rect 5868 27968 5917 27996
rect 5868 27956 5874 27968
rect 5905 27965 5917 27968
rect 5951 27965 5963 27999
rect 9401 27999 9459 28005
rect 9401 27996 9413 27999
rect 5905 27959 5963 27965
rect 9324 27968 9413 27996
rect 9324 27940 9352 27968
rect 9401 27965 9413 27968
rect 9447 27965 9459 27999
rect 9401 27959 9459 27965
rect 10045 27999 10103 28005
rect 10045 27965 10057 27999
rect 10091 27996 10103 27999
rect 12618 27996 12624 28008
rect 10091 27968 12624 27996
rect 10091 27965 10103 27968
rect 10045 27959 10103 27965
rect 12618 27956 12624 27968
rect 12676 27956 12682 28008
rect 14274 27956 14280 28008
rect 14332 27996 14338 28008
rect 14369 27999 14427 28005
rect 14369 27996 14381 27999
rect 14332 27968 14381 27996
rect 14332 27956 14338 27968
rect 14369 27965 14381 27968
rect 14415 27965 14427 27999
rect 15010 27996 15016 28008
rect 14971 27968 15016 27996
rect 14369 27959 14427 27965
rect 15010 27956 15016 27968
rect 15068 27956 15074 28008
rect 15657 27999 15715 28005
rect 15657 27965 15669 27999
rect 15703 27965 15715 27999
rect 15657 27959 15715 27965
rect 17221 27999 17279 28005
rect 17221 27965 17233 27999
rect 17267 27996 17279 27999
rect 17310 27996 17316 28008
rect 17267 27968 17316 27996
rect 17267 27965 17279 27968
rect 17221 27959 17279 27965
rect 4614 27928 4620 27940
rect 1780 27900 4620 27928
rect 4614 27888 4620 27900
rect 4672 27888 4678 27940
rect 8386 27928 8392 27940
rect 4724 27900 8392 27928
rect 1578 27860 1584 27872
rect 1539 27832 1584 27860
rect 1578 27820 1584 27832
rect 1636 27820 1642 27872
rect 2130 27820 2136 27872
rect 2188 27860 2194 27872
rect 4724 27860 4752 27900
rect 8386 27888 8392 27900
rect 8444 27888 8450 27940
rect 9306 27888 9312 27940
rect 9364 27888 9370 27940
rect 12986 27928 12992 27940
rect 12947 27900 12992 27928
rect 12986 27888 12992 27900
rect 13044 27888 13050 27940
rect 15562 27888 15568 27940
rect 15620 27928 15626 27940
rect 15672 27928 15700 27959
rect 17310 27956 17316 27968
rect 17368 27956 17374 28008
rect 36354 27996 36360 28008
rect 36315 27968 36360 27996
rect 36354 27956 36360 27968
rect 36412 27956 36418 28008
rect 18598 27928 18604 27940
rect 15620 27900 18604 27928
rect 15620 27888 15626 27900
rect 18598 27888 18604 27900
rect 18656 27888 18662 27940
rect 2188 27832 4752 27860
rect 4893 27863 4951 27869
rect 2188 27820 2194 27832
rect 4893 27829 4905 27863
rect 4939 27860 4951 27863
rect 5166 27860 5172 27872
rect 4939 27832 5172 27860
rect 4939 27829 4951 27832
rect 4893 27823 4951 27829
rect 5166 27820 5172 27832
rect 5224 27820 5230 27872
rect 5442 27860 5448 27872
rect 5403 27832 5448 27860
rect 5442 27820 5448 27832
rect 5500 27820 5506 27872
rect 6638 27860 6644 27872
rect 6599 27832 6644 27860
rect 6638 27820 6644 27832
rect 6696 27820 6702 27872
rect 7282 27860 7288 27872
rect 7243 27832 7288 27860
rect 7282 27820 7288 27832
rect 7340 27820 7346 27872
rect 7929 27863 7987 27869
rect 7929 27829 7941 27863
rect 7975 27860 7987 27863
rect 8202 27860 8208 27872
rect 7975 27832 8208 27860
rect 7975 27829 7987 27832
rect 7929 27823 7987 27829
rect 8202 27820 8208 27832
rect 8260 27820 8266 27872
rect 8757 27863 8815 27869
rect 8757 27829 8769 27863
rect 8803 27860 8815 27863
rect 12250 27860 12256 27872
rect 8803 27832 12256 27860
rect 8803 27829 8815 27832
rect 8757 27823 8815 27829
rect 12250 27820 12256 27832
rect 12308 27820 12314 27872
rect 16022 27820 16028 27872
rect 16080 27860 16086 27872
rect 17957 27863 18015 27869
rect 17957 27860 17969 27863
rect 16080 27832 17969 27860
rect 16080 27820 16086 27832
rect 17957 27829 17969 27832
rect 18003 27829 18015 27863
rect 19242 27860 19248 27872
rect 19203 27832 19248 27860
rect 17957 27823 18015 27829
rect 19242 27820 19248 27832
rect 19300 27820 19306 27872
rect 1104 27770 36892 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 36892 27770
rect 1104 27696 36892 27718
rect 4062 27656 4068 27668
rect 4023 27628 4068 27656
rect 4062 27616 4068 27628
rect 4120 27656 4126 27668
rect 4525 27659 4583 27665
rect 4525 27656 4537 27659
rect 4120 27628 4537 27656
rect 4120 27616 4126 27628
rect 4525 27625 4537 27628
rect 4571 27656 4583 27659
rect 5077 27659 5135 27665
rect 5077 27656 5089 27659
rect 4571 27628 5089 27656
rect 4571 27625 4583 27628
rect 4525 27619 4583 27625
rect 5077 27625 5089 27628
rect 5123 27625 5135 27659
rect 5077 27619 5135 27625
rect 5166 27616 5172 27668
rect 5224 27656 5230 27668
rect 8570 27656 8576 27668
rect 5224 27628 8576 27656
rect 5224 27616 5230 27628
rect 8570 27616 8576 27628
rect 8628 27656 8634 27668
rect 8754 27656 8760 27668
rect 8628 27628 8760 27656
rect 8628 27616 8634 27628
rect 8754 27616 8760 27628
rect 8812 27616 8818 27668
rect 12544 27628 13584 27656
rect 1670 27588 1676 27600
rect 1631 27560 1676 27588
rect 1670 27548 1676 27560
rect 1728 27548 1734 27600
rect 3145 27591 3203 27597
rect 3145 27557 3157 27591
rect 3191 27588 3203 27591
rect 7190 27588 7196 27600
rect 3191 27560 7196 27588
rect 3191 27557 3203 27560
rect 3145 27551 3203 27557
rect 7190 27548 7196 27560
rect 7248 27548 7254 27600
rect 11057 27591 11115 27597
rect 11057 27557 11069 27591
rect 11103 27588 11115 27591
rect 12434 27588 12440 27600
rect 11103 27560 12440 27588
rect 11103 27557 11115 27560
rect 11057 27551 11115 27557
rect 12434 27548 12440 27560
rect 12492 27548 12498 27600
rect 2501 27523 2559 27529
rect 2501 27489 2513 27523
rect 2547 27520 2559 27523
rect 2547 27492 4200 27520
rect 2547 27489 2559 27492
rect 2501 27483 2559 27489
rect 2406 27452 2412 27464
rect 2367 27424 2412 27452
rect 2406 27412 2412 27424
rect 2464 27412 2470 27464
rect 2866 27412 2872 27464
rect 2924 27452 2930 27464
rect 3053 27455 3111 27461
rect 3053 27452 3065 27455
rect 2924 27424 3065 27452
rect 2924 27412 2930 27424
rect 3053 27421 3065 27424
rect 3099 27421 3111 27455
rect 4172 27452 4200 27492
rect 4890 27480 4896 27532
rect 4948 27520 4954 27532
rect 4948 27492 6684 27520
rect 4948 27480 4954 27492
rect 5718 27452 5724 27464
rect 4172 27424 5724 27452
rect 3053 27415 3111 27421
rect 5718 27412 5724 27424
rect 5776 27412 5782 27464
rect 6549 27455 6607 27461
rect 6549 27421 6561 27455
rect 6595 27421 6607 27455
rect 6656 27452 6684 27492
rect 6822 27480 6828 27532
rect 6880 27520 6886 27532
rect 7837 27523 7895 27529
rect 7837 27520 7849 27523
rect 6880 27492 7849 27520
rect 6880 27480 6886 27492
rect 7837 27489 7849 27492
rect 7883 27489 7895 27523
rect 7837 27483 7895 27489
rect 8481 27523 8539 27529
rect 8481 27489 8493 27523
rect 8527 27520 8539 27523
rect 8527 27492 10364 27520
rect 8527 27489 8539 27492
rect 8481 27483 8539 27489
rect 7193 27455 7251 27461
rect 7193 27452 7205 27455
rect 6656 27424 7205 27452
rect 6549 27415 6607 27421
rect 7193 27421 7205 27424
rect 7239 27421 7251 27455
rect 7193 27415 7251 27421
rect 3694 27344 3700 27396
rect 3752 27384 3758 27396
rect 6564 27384 6592 27415
rect 3752 27356 6592 27384
rect 6641 27387 6699 27393
rect 3752 27344 3758 27356
rect 6641 27353 6653 27387
rect 6687 27384 6699 27387
rect 7650 27384 7656 27396
rect 6687 27356 7656 27384
rect 6687 27353 6699 27356
rect 6641 27347 6699 27353
rect 7650 27344 7656 27356
rect 7708 27344 7714 27396
rect 8389 27387 8447 27393
rect 8389 27353 8401 27387
rect 8435 27353 8447 27387
rect 8389 27347 8447 27353
rect 5626 27276 5632 27328
rect 5684 27316 5690 27328
rect 5905 27319 5963 27325
rect 5905 27316 5917 27319
rect 5684 27288 5917 27316
rect 5684 27276 5690 27288
rect 5905 27285 5917 27288
rect 5951 27285 5963 27319
rect 5905 27279 5963 27285
rect 7285 27319 7343 27325
rect 7285 27285 7297 27319
rect 7331 27316 7343 27319
rect 8404 27316 8432 27347
rect 9306 27344 9312 27396
rect 9364 27384 9370 27396
rect 9677 27387 9735 27393
rect 9677 27384 9689 27387
rect 9364 27356 9689 27384
rect 9364 27344 9370 27356
rect 9677 27353 9689 27356
rect 9723 27353 9735 27387
rect 9677 27347 9735 27353
rect 9766 27344 9772 27396
rect 9824 27384 9830 27396
rect 10336 27393 10364 27492
rect 10502 27480 10508 27532
rect 10560 27520 10566 27532
rect 12345 27523 12403 27529
rect 10560 27492 12296 27520
rect 10560 27480 10566 27492
rect 10965 27455 11023 27461
rect 10965 27421 10977 27455
rect 11011 27452 11023 27455
rect 11238 27452 11244 27464
rect 11011 27424 11244 27452
rect 11011 27421 11023 27424
rect 10965 27415 11023 27421
rect 11238 27412 11244 27424
rect 11296 27412 11302 27464
rect 11609 27455 11667 27461
rect 11609 27421 11621 27455
rect 11655 27452 11667 27455
rect 12158 27452 12164 27464
rect 11655 27424 12164 27452
rect 11655 27421 11667 27424
rect 11609 27415 11667 27421
rect 12158 27412 12164 27424
rect 12216 27412 12222 27464
rect 12268 27461 12296 27492
rect 12345 27489 12357 27523
rect 12391 27520 12403 27523
rect 12544 27520 12572 27628
rect 13556 27588 13584 27628
rect 13722 27616 13728 27668
rect 13780 27656 13786 27668
rect 18598 27656 18604 27668
rect 13780 27628 18460 27656
rect 18559 27628 18604 27656
rect 13780 27616 13786 27628
rect 14921 27591 14979 27597
rect 13556 27560 13860 27588
rect 12391 27492 12572 27520
rect 12391 27489 12403 27492
rect 12345 27483 12403 27489
rect 12618 27480 12624 27532
rect 12676 27520 12682 27532
rect 13265 27523 13323 27529
rect 13265 27520 13277 27523
rect 12676 27492 13277 27520
rect 12676 27480 12682 27492
rect 13265 27489 13277 27492
rect 13311 27520 13323 27523
rect 13722 27520 13728 27532
rect 13311 27492 13728 27520
rect 13311 27489 13323 27492
rect 13265 27483 13323 27489
rect 13722 27480 13728 27492
rect 13780 27480 13786 27532
rect 13832 27520 13860 27560
rect 14921 27557 14933 27591
rect 14967 27588 14979 27591
rect 15746 27588 15752 27600
rect 14967 27560 15752 27588
rect 14967 27557 14979 27560
rect 14921 27551 14979 27557
rect 15746 27548 15752 27560
rect 15804 27548 15810 27600
rect 18046 27588 18052 27600
rect 16040 27560 18052 27588
rect 15102 27520 15108 27532
rect 13832 27492 15108 27520
rect 15102 27480 15108 27492
rect 15160 27480 15166 27532
rect 15286 27480 15292 27532
rect 15344 27520 15350 27532
rect 15473 27523 15531 27529
rect 15473 27520 15485 27523
rect 15344 27492 15485 27520
rect 15344 27480 15350 27492
rect 15473 27489 15485 27492
rect 15519 27489 15531 27523
rect 15473 27483 15531 27489
rect 15654 27480 15660 27532
rect 15712 27520 15718 27532
rect 16040 27520 16068 27560
rect 18046 27548 18052 27560
rect 18104 27548 18110 27600
rect 15712 27492 16068 27520
rect 16117 27523 16175 27529
rect 15712 27480 15718 27492
rect 16117 27489 16129 27523
rect 16163 27520 16175 27523
rect 16298 27520 16304 27532
rect 16163 27492 16304 27520
rect 16163 27489 16175 27492
rect 16117 27483 16175 27489
rect 16298 27480 16304 27492
rect 16356 27520 16362 27532
rect 17957 27523 18015 27529
rect 17957 27520 17969 27523
rect 16356 27492 17969 27520
rect 16356 27480 16362 27492
rect 17957 27489 17969 27492
rect 18003 27489 18015 27523
rect 18432 27520 18460 27628
rect 18598 27616 18604 27628
rect 18656 27616 18662 27668
rect 36354 27656 36360 27668
rect 36315 27628 36360 27656
rect 36354 27616 36360 27628
rect 36412 27616 36418 27668
rect 19150 27520 19156 27532
rect 18432 27492 19156 27520
rect 17957 27483 18015 27489
rect 12253 27455 12311 27461
rect 12253 27421 12265 27455
rect 12299 27421 12311 27455
rect 14826 27452 14832 27464
rect 14787 27424 14832 27452
rect 12253 27415 12311 27421
rect 14826 27412 14832 27424
rect 14884 27412 14890 27464
rect 18049 27455 18107 27461
rect 18049 27421 18061 27455
rect 18095 27452 18107 27455
rect 18598 27452 18604 27464
rect 18095 27424 18604 27452
rect 18095 27421 18107 27424
rect 18049 27415 18107 27421
rect 18598 27412 18604 27424
rect 18656 27412 18662 27464
rect 18708 27461 18736 27492
rect 19150 27480 19156 27492
rect 19208 27520 19214 27532
rect 19429 27523 19487 27529
rect 19429 27520 19441 27523
rect 19208 27492 19441 27520
rect 19208 27480 19214 27492
rect 19429 27489 19441 27492
rect 19475 27489 19487 27523
rect 19429 27483 19487 27489
rect 18693 27455 18751 27461
rect 18693 27421 18705 27455
rect 18739 27421 18751 27455
rect 27249 27455 27307 27461
rect 18693 27415 18751 27421
rect 19352 27424 22094 27452
rect 10321 27387 10379 27393
rect 9824 27356 9869 27384
rect 9824 27344 9830 27356
rect 10321 27353 10333 27387
rect 10367 27384 10379 27387
rect 10502 27384 10508 27396
rect 10367 27356 10508 27384
rect 10367 27353 10379 27356
rect 10321 27347 10379 27353
rect 10502 27344 10508 27356
rect 10560 27344 10566 27396
rect 11701 27387 11759 27393
rect 11701 27353 11713 27387
rect 11747 27384 11759 27387
rect 12618 27384 12624 27396
rect 11747 27356 12624 27384
rect 11747 27353 11759 27356
rect 11701 27347 11759 27353
rect 12618 27344 12624 27356
rect 12676 27344 12682 27396
rect 12710 27344 12716 27396
rect 12768 27384 12774 27396
rect 12989 27387 13047 27393
rect 12989 27384 13001 27387
rect 12768 27356 13001 27384
rect 12768 27344 12774 27356
rect 12989 27353 13001 27356
rect 13035 27353 13047 27387
rect 12989 27347 13047 27353
rect 13078 27344 13084 27396
rect 13136 27384 13142 27396
rect 15654 27384 15660 27396
rect 13136 27356 13181 27384
rect 14292 27356 15660 27384
rect 13136 27344 13142 27356
rect 7331 27288 8432 27316
rect 7331 27285 7343 27288
rect 7285 27279 7343 27285
rect 12434 27276 12440 27328
rect 12492 27316 12498 27328
rect 14292 27316 14320 27356
rect 15654 27344 15660 27356
rect 15712 27344 15718 27396
rect 16022 27384 16028 27396
rect 15983 27356 16028 27384
rect 16022 27344 16028 27356
rect 16080 27344 16086 27396
rect 16669 27387 16727 27393
rect 16669 27353 16681 27387
rect 16715 27353 16727 27387
rect 17218 27384 17224 27396
rect 17179 27356 17224 27384
rect 16669 27347 16727 27353
rect 12492 27288 14320 27316
rect 14369 27319 14427 27325
rect 12492 27276 12498 27288
rect 14369 27285 14381 27319
rect 14415 27316 14427 27319
rect 14550 27316 14556 27328
rect 14415 27288 14556 27316
rect 14415 27285 14427 27288
rect 14369 27279 14427 27285
rect 14550 27276 14556 27288
rect 14608 27276 14614 27328
rect 15194 27276 15200 27328
rect 15252 27316 15258 27328
rect 16684 27316 16712 27347
rect 17218 27344 17224 27356
rect 17276 27344 17282 27396
rect 17313 27387 17371 27393
rect 17313 27353 17325 27387
rect 17359 27384 17371 27387
rect 19352 27384 19380 27424
rect 17359 27356 19380 27384
rect 22066 27384 22094 27424
rect 27249 27421 27261 27455
rect 27295 27452 27307 27455
rect 36446 27452 36452 27464
rect 27295 27424 36452 27452
rect 27295 27421 27307 27424
rect 27249 27415 27307 27421
rect 36446 27412 36452 27424
rect 36504 27412 36510 27464
rect 27157 27387 27215 27393
rect 27157 27384 27169 27387
rect 22066 27356 27169 27384
rect 17359 27353 17371 27356
rect 17313 27347 17371 27353
rect 27157 27353 27169 27356
rect 27203 27353 27215 27387
rect 27157 27347 27215 27353
rect 15252 27288 16712 27316
rect 15252 27276 15258 27288
rect 19150 27276 19156 27328
rect 19208 27316 19214 27328
rect 24854 27316 24860 27328
rect 19208 27288 24860 27316
rect 19208 27276 19214 27288
rect 24854 27276 24860 27288
rect 24912 27276 24918 27328
rect 1104 27226 36892 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 36892 27226
rect 1104 27152 36892 27174
rect 2501 27115 2559 27121
rect 2501 27081 2513 27115
rect 2547 27112 2559 27115
rect 3326 27112 3332 27124
rect 2547 27084 3332 27112
rect 2547 27081 2559 27084
rect 2501 27075 2559 27081
rect 3326 27072 3332 27084
rect 3384 27072 3390 27124
rect 3881 27115 3939 27121
rect 3881 27081 3893 27115
rect 3927 27112 3939 27115
rect 4062 27112 4068 27124
rect 3927 27084 4068 27112
rect 3927 27081 3939 27084
rect 3881 27075 3939 27081
rect 4062 27072 4068 27084
rect 4120 27112 4126 27124
rect 4341 27115 4399 27121
rect 4341 27112 4353 27115
rect 4120 27084 4353 27112
rect 4120 27072 4126 27084
rect 4341 27081 4353 27084
rect 4387 27081 4399 27115
rect 4341 27075 4399 27081
rect 9125 27115 9183 27121
rect 9125 27081 9137 27115
rect 9171 27112 9183 27115
rect 9490 27112 9496 27124
rect 9171 27084 9496 27112
rect 9171 27081 9183 27084
rect 9125 27075 9183 27081
rect 9490 27072 9496 27084
rect 9548 27072 9554 27124
rect 9766 27072 9772 27124
rect 9824 27112 9830 27124
rect 10413 27115 10471 27121
rect 10413 27112 10425 27115
rect 9824 27084 10425 27112
rect 9824 27072 9830 27084
rect 10413 27081 10425 27084
rect 10459 27081 10471 27115
rect 10413 27075 10471 27081
rect 10502 27072 10508 27124
rect 10560 27112 10566 27124
rect 14274 27112 14280 27124
rect 10560 27084 14280 27112
rect 10560 27072 10566 27084
rect 14274 27072 14280 27084
rect 14332 27072 14338 27124
rect 14550 27072 14556 27124
rect 14608 27112 14614 27124
rect 15838 27112 15844 27124
rect 14608 27084 15844 27112
rect 14608 27072 14614 27084
rect 15838 27072 15844 27084
rect 15896 27072 15902 27124
rect 16298 27072 16304 27124
rect 16356 27072 16362 27124
rect 18782 27112 18788 27124
rect 18743 27084 18788 27112
rect 18782 27072 18788 27084
rect 18840 27072 18846 27124
rect 35986 27072 35992 27124
rect 36044 27112 36050 27124
rect 36173 27115 36231 27121
rect 36173 27112 36185 27115
rect 36044 27084 36185 27112
rect 36044 27072 36050 27084
rect 36173 27081 36185 27084
rect 36219 27081 36231 27115
rect 36173 27075 36231 27081
rect 6270 27004 6276 27056
rect 6328 27044 6334 27056
rect 7745 27047 7803 27053
rect 7745 27044 7757 27047
rect 6328 27016 7757 27044
rect 6328 27004 6334 27016
rect 7745 27013 7757 27016
rect 7791 27013 7803 27047
rect 7745 27007 7803 27013
rect 7837 27047 7895 27053
rect 7837 27013 7849 27047
rect 7883 27044 7895 27047
rect 12710 27044 12716 27056
rect 7883 27016 12572 27044
rect 12671 27016 12716 27044
rect 7883 27013 7895 27016
rect 7837 27007 7895 27013
rect 1578 26976 1584 26988
rect 1539 26948 1584 26976
rect 1578 26936 1584 26948
rect 1636 26936 1642 26988
rect 2130 26936 2136 26988
rect 2188 26976 2194 26988
rect 2317 26979 2375 26985
rect 2317 26976 2329 26979
rect 2188 26948 2329 26976
rect 2188 26936 2194 26948
rect 2317 26945 2329 26948
rect 2363 26945 2375 26979
rect 9030 26976 9036 26988
rect 8991 26948 9036 26976
rect 2317 26939 2375 26945
rect 9030 26936 9036 26948
rect 9088 26976 9094 26988
rect 9677 26979 9735 26985
rect 9677 26976 9689 26979
rect 9088 26948 9689 26976
rect 9088 26936 9094 26948
rect 9677 26945 9689 26948
rect 9723 26945 9735 26979
rect 10502 26976 10508 26988
rect 10463 26948 10508 26976
rect 9677 26939 9735 26945
rect 10502 26936 10508 26948
rect 10560 26936 10566 26988
rect 11977 26979 12035 26985
rect 11977 26945 11989 26979
rect 12023 26976 12035 26979
rect 12434 26976 12440 26988
rect 12023 26948 12440 26976
rect 12023 26945 12035 26948
rect 11977 26939 12035 26945
rect 6822 26868 6828 26920
rect 6880 26908 6886 26920
rect 7193 26911 7251 26917
rect 7193 26908 7205 26911
rect 6880 26880 7205 26908
rect 6880 26868 6886 26880
rect 7193 26877 7205 26880
rect 7239 26877 7251 26911
rect 8570 26908 8576 26920
rect 8483 26880 8576 26908
rect 7193 26871 7251 26877
rect 8570 26868 8576 26880
rect 8628 26908 8634 26920
rect 11992 26908 12020 26939
rect 12434 26936 12440 26948
rect 12492 26936 12498 26988
rect 8628 26880 12020 26908
rect 12544 26908 12572 27016
rect 12710 27004 12716 27016
rect 12768 27004 12774 27056
rect 12805 27047 12863 27053
rect 12805 27013 12817 27047
rect 12851 27044 12863 27047
rect 13078 27044 13084 27056
rect 12851 27016 13084 27044
rect 12851 27013 12863 27016
rect 12805 27007 12863 27013
rect 13078 27004 13084 27016
rect 13136 27004 13142 27056
rect 13722 27004 13728 27056
rect 13780 27044 13786 27056
rect 13817 27047 13875 27053
rect 13817 27044 13829 27047
rect 13780 27016 13829 27044
rect 13780 27004 13786 27016
rect 13817 27013 13829 27016
rect 13863 27013 13875 27047
rect 14366 27044 14372 27056
rect 14327 27016 14372 27044
rect 13817 27007 13875 27013
rect 14366 27004 14372 27016
rect 14424 27004 14430 27056
rect 16114 27044 16120 27056
rect 16075 27016 16120 27044
rect 16114 27004 16120 27016
rect 16172 27004 16178 27056
rect 16209 27047 16267 27053
rect 16209 27013 16221 27047
rect 16255 27044 16267 27047
rect 16316 27044 16344 27072
rect 16255 27016 16344 27044
rect 17037 27047 17095 27053
rect 16255 27013 16267 27016
rect 16209 27007 16267 27013
rect 17037 27013 17049 27047
rect 17083 27044 17095 27047
rect 17126 27044 17132 27056
rect 17083 27016 17132 27044
rect 17083 27013 17095 27016
rect 17037 27007 17095 27013
rect 17126 27004 17132 27016
rect 17184 27004 17190 27056
rect 17957 27047 18015 27053
rect 17957 27013 17969 27047
rect 18003 27044 18015 27047
rect 18414 27044 18420 27056
rect 18003 27016 18420 27044
rect 18003 27013 18015 27016
rect 17957 27007 18015 27013
rect 18414 27004 18420 27016
rect 18472 27004 18478 27056
rect 26142 27044 26148 27056
rect 22066 27016 26148 27044
rect 14734 26936 14740 26988
rect 14792 26976 14798 26988
rect 15010 26976 15016 26988
rect 14792 26948 15016 26976
rect 14792 26936 14798 26948
rect 15010 26936 15016 26948
rect 15068 26936 15074 26988
rect 16482 26936 16488 26988
rect 16540 26976 16546 26988
rect 18598 26976 18604 26988
rect 16540 26948 17172 26976
rect 18511 26948 18604 26976
rect 16540 26936 16546 26948
rect 14461 26911 14519 26917
rect 12544 26880 14412 26908
rect 8628 26868 8634 26880
rect 6730 26800 6736 26852
rect 6788 26840 6794 26852
rect 9582 26840 9588 26852
rect 6788 26812 9588 26840
rect 6788 26800 6794 26812
rect 9582 26800 9588 26812
rect 9640 26800 9646 26852
rect 10870 26840 10876 26852
rect 9692 26812 10876 26840
rect 1762 26772 1768 26784
rect 1723 26744 1768 26772
rect 1762 26732 1768 26744
rect 1820 26732 1826 26784
rect 5626 26732 5632 26784
rect 5684 26772 5690 26784
rect 9692 26772 9720 26812
rect 10870 26800 10876 26812
rect 10928 26840 10934 26852
rect 11057 26843 11115 26849
rect 11057 26840 11069 26843
rect 10928 26812 11069 26840
rect 10928 26800 10934 26812
rect 11057 26809 11069 26812
rect 11103 26809 11115 26843
rect 11057 26803 11115 26809
rect 12158 26800 12164 26852
rect 12216 26840 12222 26852
rect 13262 26840 13268 26852
rect 12216 26812 13268 26840
rect 12216 26800 12222 26812
rect 13262 26800 13268 26812
rect 13320 26800 13326 26852
rect 14384 26840 14412 26880
rect 14461 26877 14473 26911
rect 14507 26908 14519 26911
rect 15933 26911 15991 26917
rect 14507 26880 15608 26908
rect 14507 26877 14519 26880
rect 14461 26871 14519 26877
rect 15194 26840 15200 26852
rect 14384 26812 15200 26840
rect 15194 26800 15200 26812
rect 15252 26800 15258 26852
rect 15580 26784 15608 26880
rect 15933 26877 15945 26911
rect 15979 26908 15991 26911
rect 16206 26908 16212 26920
rect 15979 26880 16212 26908
rect 15979 26877 15991 26880
rect 15933 26871 15991 26877
rect 16206 26868 16212 26880
rect 16264 26868 16270 26920
rect 17144 26908 17172 26948
rect 18598 26936 18604 26948
rect 18656 26976 18662 26988
rect 19242 26976 19248 26988
rect 18656 26948 19248 26976
rect 18656 26936 18662 26948
rect 19242 26936 19248 26948
rect 19300 26936 19306 26988
rect 17494 26908 17500 26920
rect 17144 26880 17500 26908
rect 17494 26868 17500 26880
rect 17552 26908 17558 26920
rect 18049 26911 18107 26917
rect 18049 26908 18061 26911
rect 17552 26880 18061 26908
rect 17552 26868 17558 26880
rect 18049 26877 18061 26880
rect 18095 26877 18107 26911
rect 18049 26871 18107 26877
rect 16114 26800 16120 26852
rect 16172 26840 16178 26852
rect 17862 26840 17868 26852
rect 16172 26812 17868 26840
rect 16172 26800 16178 26812
rect 17862 26800 17868 26812
rect 17920 26800 17926 26852
rect 22066 26840 22094 27016
rect 26142 27004 26148 27016
rect 26200 27004 26206 27056
rect 35713 26979 35771 26985
rect 35713 26945 35725 26979
rect 35759 26976 35771 26979
rect 36354 26976 36360 26988
rect 35759 26948 36360 26976
rect 35759 26945 35771 26948
rect 35713 26939 35771 26945
rect 36354 26936 36360 26948
rect 36412 26936 36418 26988
rect 17972 26812 22094 26840
rect 5684 26744 9720 26772
rect 9769 26775 9827 26781
rect 5684 26732 5690 26744
rect 9769 26741 9781 26775
rect 9815 26772 9827 26775
rect 10594 26772 10600 26784
rect 9815 26744 10600 26772
rect 9815 26741 9827 26744
rect 9769 26735 9827 26741
rect 10594 26732 10600 26744
rect 10652 26732 10658 26784
rect 12069 26775 12127 26781
rect 12069 26741 12081 26775
rect 12115 26772 12127 26775
rect 13538 26772 13544 26784
rect 12115 26744 13544 26772
rect 12115 26741 12127 26744
rect 12069 26735 12127 26741
rect 13538 26732 13544 26744
rect 13596 26732 13602 26784
rect 13814 26732 13820 26784
rect 13872 26772 13878 26784
rect 15470 26772 15476 26784
rect 13872 26744 15476 26772
rect 13872 26732 13878 26744
rect 15470 26732 15476 26744
rect 15528 26732 15534 26784
rect 15562 26732 15568 26784
rect 15620 26772 15626 26784
rect 17972 26772 18000 26812
rect 19242 26772 19248 26784
rect 15620 26744 18000 26772
rect 19203 26744 19248 26772
rect 15620 26732 15626 26744
rect 19242 26732 19248 26744
rect 19300 26732 19306 26784
rect 1104 26682 36892 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 36892 26682
rect 1104 26608 36892 26630
rect 1486 26528 1492 26580
rect 1544 26568 1550 26580
rect 1581 26571 1639 26577
rect 1581 26568 1593 26571
rect 1544 26540 1593 26568
rect 1544 26528 1550 26540
rect 1581 26537 1593 26540
rect 1627 26537 1639 26571
rect 2222 26568 2228 26580
rect 2183 26540 2228 26568
rect 1581 26531 1639 26537
rect 2222 26528 2228 26540
rect 2280 26528 2286 26580
rect 6270 26568 6276 26580
rect 6231 26540 6276 26568
rect 6270 26528 6276 26540
rect 6328 26528 6334 26580
rect 6362 26528 6368 26580
rect 6420 26568 6426 26580
rect 8294 26568 8300 26580
rect 6420 26540 8300 26568
rect 6420 26528 6426 26540
rect 8294 26528 8300 26540
rect 8352 26528 8358 26580
rect 8389 26571 8447 26577
rect 8389 26537 8401 26571
rect 8435 26568 8447 26571
rect 9306 26568 9312 26580
rect 8435 26540 9312 26568
rect 8435 26537 8447 26540
rect 8389 26531 8447 26537
rect 9306 26528 9312 26540
rect 9364 26528 9370 26580
rect 12526 26568 12532 26580
rect 9416 26540 12532 26568
rect 1762 26460 1768 26512
rect 1820 26500 1826 26512
rect 1820 26472 8340 26500
rect 1820 26460 1826 26472
rect 2590 26324 2596 26376
rect 2648 26364 2654 26376
rect 8312 26373 8340 26472
rect 6181 26367 6239 26373
rect 6181 26364 6193 26367
rect 2648 26336 6193 26364
rect 2648 26324 2654 26336
rect 6181 26333 6193 26336
rect 6227 26333 6239 26367
rect 6181 26327 6239 26333
rect 8297 26367 8355 26373
rect 8297 26333 8309 26367
rect 8343 26333 8355 26367
rect 8297 26327 8355 26333
rect 6086 26256 6092 26308
rect 6144 26296 6150 26308
rect 6822 26296 6828 26308
rect 6144 26268 6828 26296
rect 6144 26256 6150 26268
rect 6822 26256 6828 26268
rect 6880 26296 6886 26308
rect 7101 26299 7159 26305
rect 7101 26296 7113 26299
rect 6880 26268 7113 26296
rect 6880 26256 6886 26268
rect 7101 26265 7113 26268
rect 7147 26265 7159 26299
rect 7650 26296 7656 26308
rect 7611 26268 7656 26296
rect 7101 26259 7159 26265
rect 7650 26256 7656 26268
rect 7708 26256 7714 26308
rect 7745 26299 7803 26305
rect 7745 26265 7757 26299
rect 7791 26296 7803 26299
rect 9416 26296 9444 26540
rect 12526 26528 12532 26540
rect 12584 26528 12590 26580
rect 12820 26540 18368 26568
rect 9582 26460 9588 26512
rect 9640 26500 9646 26512
rect 12820 26500 12848 26540
rect 9640 26472 12848 26500
rect 9640 26460 9646 26472
rect 13262 26460 13268 26512
rect 13320 26500 13326 26512
rect 15013 26503 15071 26509
rect 15013 26500 15025 26503
rect 13320 26472 15025 26500
rect 13320 26460 13326 26472
rect 15013 26469 15025 26472
rect 15059 26469 15071 26503
rect 15013 26463 15071 26469
rect 15470 26460 15476 26512
rect 15528 26500 15534 26512
rect 15528 26472 16436 26500
rect 15528 26460 15534 26472
rect 11422 26432 11428 26444
rect 11383 26404 11428 26432
rect 11422 26392 11428 26404
rect 11480 26392 11486 26444
rect 12069 26435 12127 26441
rect 12069 26401 12081 26435
rect 12115 26432 12127 26435
rect 12158 26432 12164 26444
rect 12115 26404 12164 26432
rect 12115 26401 12127 26404
rect 12069 26395 12127 26401
rect 12158 26392 12164 26404
rect 12216 26392 12222 26444
rect 14369 26435 14427 26441
rect 14369 26401 14381 26435
rect 14415 26432 14427 26435
rect 15286 26432 15292 26444
rect 14415 26404 15292 26432
rect 14415 26401 14427 26404
rect 14369 26395 14427 26401
rect 15286 26392 15292 26404
rect 15344 26392 15350 26444
rect 15562 26432 15568 26444
rect 15523 26404 15568 26432
rect 15562 26392 15568 26404
rect 15620 26392 15626 26444
rect 9769 26367 9827 26373
rect 9769 26333 9781 26367
rect 9815 26364 9827 26367
rect 10410 26364 10416 26376
rect 9815 26336 10416 26364
rect 9815 26333 9827 26336
rect 9769 26327 9827 26333
rect 10410 26324 10416 26336
rect 10468 26324 10474 26376
rect 10686 26364 10692 26376
rect 10647 26336 10692 26364
rect 10686 26324 10692 26336
rect 10744 26324 10750 26376
rect 12710 26324 12716 26376
rect 12768 26364 12774 26376
rect 12894 26364 12900 26376
rect 12768 26336 12900 26364
rect 12768 26324 12774 26336
rect 12894 26324 12900 26336
rect 12952 26324 12958 26376
rect 14277 26367 14335 26373
rect 14277 26333 14289 26367
rect 14323 26364 14335 26367
rect 14826 26364 14832 26376
rect 14323 26336 14832 26364
rect 14323 26333 14335 26336
rect 14277 26327 14335 26333
rect 14826 26324 14832 26336
rect 14884 26324 14890 26376
rect 16408 26374 16436 26472
rect 16850 26460 16856 26512
rect 16908 26500 16914 26512
rect 18230 26500 18236 26512
rect 16908 26472 18236 26500
rect 16908 26460 16914 26472
rect 18230 26460 18236 26472
rect 18288 26460 18294 26512
rect 16577 26435 16635 26441
rect 16577 26401 16589 26435
rect 16623 26432 16635 26435
rect 17221 26435 17279 26441
rect 16623 26404 17080 26432
rect 16623 26401 16635 26404
rect 16577 26395 16635 26401
rect 16408 26373 16528 26374
rect 16408 26367 16543 26373
rect 16408 26346 16497 26367
rect 16485 26333 16497 26346
rect 16531 26364 16543 26367
rect 16531 26336 16988 26364
rect 16531 26333 16543 26336
rect 16485 26327 16543 26333
rect 7791 26268 9444 26296
rect 7791 26265 7803 26268
rect 7745 26259 7803 26265
rect 9490 26256 9496 26308
rect 9548 26296 9554 26308
rect 9677 26299 9735 26305
rect 9677 26296 9689 26299
rect 9548 26268 9689 26296
rect 9548 26256 9554 26268
rect 9677 26265 9689 26268
rect 9723 26265 9735 26299
rect 9677 26259 9735 26265
rect 10781 26299 10839 26305
rect 10781 26265 10793 26299
rect 10827 26296 10839 26299
rect 11517 26299 11575 26305
rect 10827 26268 11376 26296
rect 10827 26265 10839 26268
rect 10781 26259 10839 26265
rect 11348 26228 11376 26268
rect 11517 26265 11529 26299
rect 11563 26265 11575 26299
rect 12986 26296 12992 26308
rect 12947 26268 12992 26296
rect 11517 26259 11575 26265
rect 11532 26228 11560 26259
rect 12986 26256 12992 26268
rect 13044 26256 13050 26308
rect 13538 26296 13544 26308
rect 13499 26268 13544 26296
rect 13538 26256 13544 26268
rect 13596 26256 13602 26308
rect 13633 26299 13691 26305
rect 13633 26265 13645 26299
rect 13679 26296 13691 26299
rect 13998 26296 14004 26308
rect 13679 26268 14004 26296
rect 13679 26265 13691 26268
rect 13633 26259 13691 26265
rect 13998 26256 14004 26268
rect 14056 26256 14062 26308
rect 15473 26299 15531 26305
rect 15473 26265 15485 26299
rect 15519 26296 15531 26299
rect 16850 26296 16856 26308
rect 15519 26268 16856 26296
rect 15519 26265 15531 26268
rect 15473 26259 15531 26265
rect 16850 26256 16856 26268
rect 16908 26256 16914 26308
rect 11348 26200 11560 26228
rect 12526 26188 12532 26240
rect 12584 26228 12590 26240
rect 15378 26228 15384 26240
rect 12584 26200 15384 26228
rect 12584 26188 12590 26200
rect 15378 26188 15384 26200
rect 15436 26188 15442 26240
rect 16960 26228 16988 26336
rect 17052 26296 17080 26404
rect 17221 26401 17233 26435
rect 17267 26432 17279 26435
rect 17310 26432 17316 26444
rect 17267 26404 17316 26432
rect 17267 26401 17279 26404
rect 17221 26395 17279 26401
rect 17310 26392 17316 26404
rect 17368 26392 17374 26444
rect 17494 26432 17500 26444
rect 17455 26404 17500 26432
rect 17494 26392 17500 26404
rect 17552 26392 17558 26444
rect 18340 26432 18368 26540
rect 19429 26435 19487 26441
rect 19429 26432 19441 26435
rect 18340 26404 19441 26432
rect 18340 26364 18368 26404
rect 18509 26367 18567 26373
rect 18509 26364 18521 26367
rect 18340 26336 18521 26364
rect 18509 26333 18521 26336
rect 18555 26333 18567 26367
rect 18509 26327 18567 26333
rect 17313 26299 17371 26305
rect 17313 26296 17325 26299
rect 17052 26268 17325 26296
rect 17313 26265 17325 26268
rect 17359 26265 17371 26299
rect 17954 26296 17960 26308
rect 17313 26259 17371 26265
rect 17420 26268 17960 26296
rect 17420 26228 17448 26268
rect 17954 26256 17960 26268
rect 18012 26256 18018 26308
rect 18414 26296 18420 26308
rect 18375 26268 18420 26296
rect 18414 26256 18420 26268
rect 18472 26256 18478 26308
rect 19168 26296 19196 26404
rect 19429 26401 19441 26404
rect 19475 26401 19487 26435
rect 19429 26395 19487 26401
rect 19242 26324 19248 26376
rect 19300 26364 19306 26376
rect 32398 26364 32404 26376
rect 19300 26336 32404 26364
rect 19300 26324 19306 26336
rect 32398 26324 32404 26336
rect 32456 26324 32462 26376
rect 35526 26296 35532 26308
rect 19168 26268 35532 26296
rect 35526 26256 35532 26268
rect 35584 26256 35590 26308
rect 19978 26228 19984 26240
rect 16960 26200 17448 26228
rect 19939 26200 19984 26228
rect 19978 26188 19984 26200
rect 20036 26188 20042 26240
rect 1104 26138 36892 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 36892 26138
rect 1104 26064 36892 26086
rect 8294 25984 8300 26036
rect 8352 26024 8358 26036
rect 9125 26027 9183 26033
rect 9125 26024 9137 26027
rect 8352 25996 9137 26024
rect 8352 25984 8358 25996
rect 9125 25993 9137 25996
rect 9171 26024 9183 26027
rect 10502 26024 10508 26036
rect 9171 25996 10508 26024
rect 9171 25993 9183 25996
rect 9125 25987 9183 25993
rect 10502 25984 10508 25996
rect 10560 25984 10566 26036
rect 10962 25984 10968 26036
rect 11020 26024 11026 26036
rect 17218 26024 17224 26036
rect 11020 25996 12296 26024
rect 11020 25984 11026 25996
rect 12158 25956 12164 25968
rect 12119 25928 12164 25956
rect 12158 25916 12164 25928
rect 12216 25916 12222 25968
rect 12268 25965 12296 25996
rect 14108 25996 15424 26024
rect 17179 25996 17224 26024
rect 14108 25965 14136 25996
rect 12253 25959 12311 25965
rect 12253 25925 12265 25959
rect 12299 25925 12311 25959
rect 12253 25919 12311 25925
rect 14093 25959 14151 25965
rect 14093 25925 14105 25959
rect 14139 25925 14151 25959
rect 15286 25956 15292 25968
rect 15247 25928 15292 25956
rect 14093 25919 14151 25925
rect 15286 25916 15292 25928
rect 15344 25916 15350 25968
rect 15396 25956 15424 25996
rect 17218 25984 17224 25996
rect 17276 25984 17282 26036
rect 17862 26024 17868 26036
rect 17823 25996 17868 26024
rect 17862 25984 17868 25996
rect 17920 25984 17926 26036
rect 18509 25959 18567 25965
rect 18509 25956 18521 25959
rect 15396 25928 18521 25956
rect 18509 25925 18521 25928
rect 18555 25925 18567 25959
rect 18509 25919 18567 25925
rect 10226 25888 10232 25900
rect 10187 25860 10232 25888
rect 10226 25848 10232 25860
rect 10284 25888 10290 25900
rect 10965 25891 11023 25897
rect 10965 25888 10977 25891
rect 10284 25860 10977 25888
rect 10284 25848 10290 25860
rect 10965 25857 10977 25860
rect 11011 25857 11023 25891
rect 10965 25851 11023 25857
rect 17129 25891 17187 25897
rect 17129 25857 17141 25891
rect 17175 25857 17187 25891
rect 17954 25888 17960 25900
rect 17915 25860 17960 25888
rect 17129 25851 17187 25857
rect 10502 25780 10508 25832
rect 10560 25820 10566 25832
rect 13170 25820 13176 25832
rect 10560 25792 12434 25820
rect 13131 25792 13176 25820
rect 10560 25780 10566 25792
rect 10321 25755 10379 25761
rect 10321 25721 10333 25755
rect 10367 25752 10379 25755
rect 12066 25752 12072 25764
rect 10367 25724 12072 25752
rect 10367 25721 10379 25724
rect 10321 25715 10379 25721
rect 12066 25712 12072 25724
rect 12124 25712 12130 25764
rect 9766 25684 9772 25696
rect 9727 25656 9772 25684
rect 9766 25644 9772 25656
rect 9824 25644 9830 25696
rect 11054 25684 11060 25696
rect 11015 25656 11060 25684
rect 11054 25644 11060 25656
rect 11112 25644 11118 25696
rect 12406 25684 12434 25792
rect 13170 25780 13176 25792
rect 13228 25780 13234 25832
rect 13998 25820 14004 25832
rect 13959 25792 14004 25820
rect 13998 25780 14004 25792
rect 14056 25780 14062 25832
rect 14918 25780 14924 25832
rect 14976 25820 14982 25832
rect 15197 25823 15255 25829
rect 15197 25820 15209 25823
rect 14976 25792 15209 25820
rect 14976 25780 14982 25792
rect 15197 25789 15209 25792
rect 15243 25789 15255 25823
rect 15197 25783 15255 25789
rect 15473 25823 15531 25829
rect 15473 25789 15485 25823
rect 15519 25789 15531 25823
rect 15473 25783 15531 25789
rect 13630 25712 13636 25764
rect 13688 25752 13694 25764
rect 14553 25755 14611 25761
rect 14553 25752 14565 25755
rect 13688 25724 14565 25752
rect 13688 25712 13694 25724
rect 14553 25721 14565 25724
rect 14599 25752 14611 25755
rect 15488 25752 15516 25783
rect 14599 25724 15516 25752
rect 17144 25752 17172 25851
rect 17954 25848 17960 25860
rect 18012 25888 18018 25900
rect 18601 25891 18659 25897
rect 18601 25888 18613 25891
rect 18012 25860 18613 25888
rect 18012 25848 18018 25860
rect 18601 25857 18613 25860
rect 18647 25888 18659 25891
rect 19061 25891 19119 25897
rect 19061 25888 19073 25891
rect 18647 25860 19073 25888
rect 18647 25857 18659 25860
rect 18601 25851 18659 25857
rect 19061 25857 19073 25860
rect 19107 25888 19119 25891
rect 19613 25891 19671 25897
rect 19613 25888 19625 25891
rect 19107 25860 19625 25888
rect 19107 25857 19119 25860
rect 19061 25851 19119 25857
rect 19613 25857 19625 25860
rect 19659 25888 19671 25891
rect 19978 25888 19984 25900
rect 19659 25860 19984 25888
rect 19659 25857 19671 25860
rect 19613 25851 19671 25857
rect 19978 25848 19984 25860
rect 20036 25848 20042 25900
rect 20165 25755 20223 25761
rect 20165 25752 20177 25755
rect 17144 25724 20177 25752
rect 14599 25721 14611 25724
rect 14553 25715 14611 25721
rect 16942 25684 16948 25696
rect 12406 25656 16948 25684
rect 16942 25644 16948 25656
rect 17000 25684 17006 25696
rect 17144 25684 17172 25724
rect 20165 25721 20177 25724
rect 20211 25721 20223 25755
rect 20165 25715 20223 25721
rect 17000 25656 17172 25684
rect 17000 25644 17006 25656
rect 1104 25594 36892 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 36892 25594
rect 1104 25520 36892 25542
rect 11057 25483 11115 25489
rect 11057 25449 11069 25483
rect 11103 25480 11115 25483
rect 13078 25480 13084 25492
rect 11103 25452 13084 25480
rect 11103 25449 11115 25452
rect 11057 25443 11115 25449
rect 13078 25440 13084 25452
rect 13136 25440 13142 25492
rect 14642 25440 14648 25492
rect 14700 25480 14706 25492
rect 18230 25480 18236 25492
rect 14700 25452 18000 25480
rect 18191 25452 18236 25480
rect 14700 25440 14706 25452
rect 9769 25415 9827 25421
rect 9769 25381 9781 25415
rect 9815 25412 9827 25415
rect 11790 25412 11796 25424
rect 9815 25384 11796 25412
rect 9815 25381 9827 25384
rect 9769 25375 9827 25381
rect 11790 25372 11796 25384
rect 11848 25412 11854 25424
rect 12897 25415 12955 25421
rect 12897 25412 12909 25415
rect 11848 25384 12909 25412
rect 11848 25372 11854 25384
rect 12897 25381 12909 25384
rect 12943 25381 12955 25415
rect 15194 25412 15200 25424
rect 15155 25384 15200 25412
rect 12897 25375 12955 25381
rect 15194 25372 15200 25384
rect 15252 25412 15258 25424
rect 16393 25415 16451 25421
rect 16393 25412 16405 25415
rect 15252 25384 16405 25412
rect 15252 25372 15258 25384
rect 16393 25381 16405 25384
rect 16439 25381 16451 25415
rect 16393 25375 16451 25381
rect 12253 25347 12311 25353
rect 12253 25313 12265 25347
rect 12299 25344 12311 25347
rect 13446 25344 13452 25356
rect 12299 25316 13452 25344
rect 12299 25313 12311 25316
rect 12253 25307 12311 25313
rect 13446 25304 13452 25316
rect 13504 25304 13510 25356
rect 15749 25347 15807 25353
rect 15749 25313 15761 25347
rect 15795 25344 15807 25347
rect 17862 25344 17868 25356
rect 15795 25316 17868 25344
rect 15795 25313 15807 25316
rect 15749 25307 15807 25313
rect 17862 25304 17868 25316
rect 17920 25304 17926 25356
rect 17972 25344 18000 25452
rect 18230 25440 18236 25452
rect 18288 25440 18294 25492
rect 19429 25415 19487 25421
rect 19429 25412 19441 25415
rect 19306 25384 19441 25412
rect 19306 25344 19334 25384
rect 19429 25381 19441 25384
rect 19475 25381 19487 25415
rect 19429 25375 19487 25381
rect 17972 25316 19334 25344
rect 1578 25276 1584 25288
rect 1539 25248 1584 25276
rect 1578 25236 1584 25248
rect 1636 25276 1642 25288
rect 2225 25279 2283 25285
rect 2225 25276 2237 25279
rect 1636 25248 2237 25276
rect 1636 25236 1642 25248
rect 2225 25245 2237 25248
rect 2271 25245 2283 25279
rect 2225 25239 2283 25245
rect 10134 25236 10140 25288
rect 10192 25276 10198 25288
rect 10321 25279 10379 25285
rect 10321 25276 10333 25279
rect 10192 25248 10333 25276
rect 10192 25236 10198 25248
rect 10321 25245 10333 25248
rect 10367 25245 10379 25279
rect 10321 25239 10379 25245
rect 10870 25236 10876 25288
rect 10928 25276 10934 25288
rect 10965 25279 11023 25285
rect 10965 25276 10977 25279
rect 10928 25248 10977 25276
rect 10928 25236 10934 25248
rect 10965 25245 10977 25248
rect 11011 25245 11023 25279
rect 14461 25279 14519 25285
rect 14461 25276 14473 25279
rect 10965 25239 11023 25245
rect 14384 25248 14473 25276
rect 7926 25168 7932 25220
rect 7984 25208 7990 25220
rect 9217 25211 9275 25217
rect 9217 25208 9229 25211
rect 7984 25180 9229 25208
rect 7984 25168 7990 25180
rect 9217 25177 9229 25180
rect 9263 25177 9275 25211
rect 9217 25171 9275 25177
rect 9306 25168 9312 25220
rect 9364 25208 9370 25220
rect 10413 25211 10471 25217
rect 9364 25180 9409 25208
rect 9364 25168 9370 25180
rect 10413 25177 10425 25211
rect 10459 25208 10471 25211
rect 11238 25208 11244 25220
rect 10459 25180 11244 25208
rect 10459 25177 10471 25180
rect 10413 25171 10471 25177
rect 11238 25168 11244 25180
rect 11296 25168 11302 25220
rect 11606 25208 11612 25220
rect 11567 25180 11612 25208
rect 11606 25168 11612 25180
rect 11664 25168 11670 25220
rect 12158 25208 12164 25220
rect 12119 25180 12164 25208
rect 12158 25168 12164 25180
rect 12216 25168 12222 25220
rect 12618 25168 12624 25220
rect 12676 25208 12682 25220
rect 13357 25211 13415 25217
rect 13357 25208 13369 25211
rect 12676 25180 13369 25208
rect 12676 25168 12682 25180
rect 13357 25177 13369 25180
rect 13403 25177 13415 25211
rect 13357 25171 13415 25177
rect 13449 25211 13507 25217
rect 13449 25177 13461 25211
rect 13495 25208 13507 25211
rect 13722 25208 13728 25220
rect 13495 25180 13728 25208
rect 13495 25177 13507 25180
rect 13449 25171 13507 25177
rect 13722 25168 13728 25180
rect 13780 25168 13786 25220
rect 14384 25152 14412 25248
rect 14461 25245 14473 25248
rect 14507 25276 14519 25279
rect 15010 25276 15016 25288
rect 14507 25248 15016 25276
rect 14507 25245 14519 25248
rect 14461 25239 14519 25245
rect 15010 25236 15016 25248
rect 15068 25236 15074 25288
rect 17681 25279 17739 25285
rect 17681 25245 17693 25279
rect 17727 25276 17739 25279
rect 17972 25276 18000 25316
rect 18322 25276 18328 25288
rect 17727 25248 18000 25276
rect 18283 25248 18328 25276
rect 17727 25245 17739 25248
rect 17681 25239 17739 25245
rect 18322 25236 18328 25248
rect 18380 25276 18386 25288
rect 18785 25279 18843 25285
rect 18785 25276 18797 25279
rect 18380 25248 18797 25276
rect 18380 25236 18386 25248
rect 18785 25245 18797 25248
rect 18831 25245 18843 25279
rect 18785 25239 18843 25245
rect 15657 25211 15715 25217
rect 15657 25177 15669 25211
rect 15703 25177 15715 25211
rect 16850 25208 16856 25220
rect 16811 25180 16856 25208
rect 15657 25171 15715 25177
rect 1762 25140 1768 25152
rect 1675 25112 1768 25140
rect 1762 25100 1768 25112
rect 1820 25140 1826 25152
rect 2498 25140 2504 25152
rect 1820 25112 2504 25140
rect 1820 25100 1826 25112
rect 2498 25100 2504 25112
rect 2556 25100 2562 25152
rect 9766 25100 9772 25152
rect 9824 25140 9830 25152
rect 14366 25140 14372 25152
rect 9824 25112 14372 25140
rect 9824 25100 9830 25112
rect 14366 25100 14372 25112
rect 14424 25100 14430 25152
rect 14553 25143 14611 25149
rect 14553 25109 14565 25143
rect 14599 25140 14611 25143
rect 15672 25140 15700 25171
rect 16850 25168 16856 25180
rect 16908 25168 16914 25220
rect 16945 25211 17003 25217
rect 16945 25177 16957 25211
rect 16991 25208 17003 25211
rect 17494 25208 17500 25220
rect 16991 25180 17500 25208
rect 16991 25177 17003 25180
rect 16945 25171 17003 25177
rect 17494 25168 17500 25180
rect 17552 25168 17558 25220
rect 14599 25112 15700 25140
rect 14599 25109 14611 25112
rect 14553 25103 14611 25109
rect 16574 25100 16580 25152
rect 16632 25140 16638 25152
rect 17589 25143 17647 25149
rect 17589 25140 17601 25143
rect 16632 25112 17601 25140
rect 16632 25100 16638 25112
rect 17589 25109 17601 25112
rect 17635 25109 17647 25143
rect 17589 25103 17647 25109
rect 1104 25050 36892 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 36892 25050
rect 1104 24976 36892 24998
rect 9033 24939 9091 24945
rect 9033 24905 9045 24939
rect 9079 24936 9091 24939
rect 9306 24936 9312 24948
rect 9079 24908 9312 24936
rect 9079 24905 9091 24908
rect 9033 24899 9091 24905
rect 9306 24896 9312 24908
rect 9364 24896 9370 24948
rect 11793 24939 11851 24945
rect 11793 24905 11805 24939
rect 11839 24936 11851 24939
rect 12526 24936 12532 24948
rect 11839 24908 12532 24936
rect 11839 24905 11851 24908
rect 11793 24899 11851 24905
rect 12526 24896 12532 24908
rect 12584 24896 12590 24948
rect 15102 24896 15108 24948
rect 15160 24936 15166 24948
rect 15160 24908 17448 24936
rect 15160 24896 15166 24908
rect 10134 24868 10140 24880
rect 9692 24840 10140 24868
rect 8386 24760 8392 24812
rect 8444 24800 8450 24812
rect 8481 24803 8539 24809
rect 8481 24800 8493 24803
rect 8444 24772 8493 24800
rect 8444 24760 8450 24772
rect 8481 24769 8493 24772
rect 8527 24800 8539 24803
rect 8662 24800 8668 24812
rect 8527 24772 8668 24800
rect 8527 24769 8539 24772
rect 8481 24763 8539 24769
rect 8662 24760 8668 24772
rect 8720 24760 8726 24812
rect 9125 24803 9183 24809
rect 9125 24769 9137 24803
rect 9171 24800 9183 24803
rect 9692 24800 9720 24840
rect 10134 24828 10140 24840
rect 10192 24828 10198 24880
rect 10594 24868 10600 24880
rect 10555 24840 10600 24868
rect 10594 24828 10600 24840
rect 10652 24828 10658 24880
rect 12437 24871 12495 24877
rect 12437 24868 12449 24871
rect 11716 24840 12449 24868
rect 9171 24772 9720 24800
rect 9769 24803 9827 24809
rect 9171 24769 9183 24772
rect 9125 24763 9183 24769
rect 9769 24769 9781 24803
rect 9815 24769 9827 24803
rect 11716 24800 11744 24840
rect 12437 24837 12449 24840
rect 12483 24837 12495 24871
rect 12437 24831 12495 24837
rect 16117 24871 16175 24877
rect 16117 24837 16129 24871
rect 16163 24868 16175 24871
rect 16574 24868 16580 24880
rect 16163 24840 16580 24868
rect 16163 24837 16175 24840
rect 16117 24831 16175 24837
rect 16574 24828 16580 24840
rect 16632 24828 16638 24880
rect 17420 24877 17448 24908
rect 17405 24871 17463 24877
rect 17405 24837 17417 24871
rect 17451 24837 17463 24871
rect 17405 24831 17463 24837
rect 9769 24763 9827 24769
rect 11624 24772 11744 24800
rect 14277 24803 14335 24809
rect 8680 24732 8708 24760
rect 9784 24732 9812 24763
rect 10502 24732 10508 24744
rect 8680 24704 9812 24732
rect 10463 24704 10508 24732
rect 10502 24692 10508 24704
rect 10560 24692 10566 24744
rect 11624 24732 11652 24772
rect 14277 24769 14289 24803
rect 14323 24769 14335 24803
rect 14277 24763 14335 24769
rect 10980 24704 11652 24732
rect 9674 24624 9680 24676
rect 9732 24664 9738 24676
rect 10980 24664 11008 24704
rect 11698 24692 11704 24744
rect 11756 24732 11762 24744
rect 12345 24735 12403 24741
rect 12345 24732 12357 24735
rect 11756 24704 12357 24732
rect 11756 24692 11762 24704
rect 12345 24701 12357 24704
rect 12391 24701 12403 24735
rect 13170 24732 13176 24744
rect 13131 24704 13176 24732
rect 12345 24695 12403 24701
rect 13170 24692 13176 24704
rect 13228 24692 13234 24744
rect 14292 24732 14320 24763
rect 14366 24760 14372 24812
rect 14424 24800 14430 24812
rect 14921 24803 14979 24809
rect 14921 24800 14933 24803
rect 14424 24772 14933 24800
rect 14424 24760 14430 24772
rect 14921 24769 14933 24772
rect 14967 24769 14979 24803
rect 14921 24763 14979 24769
rect 17862 24760 17868 24812
rect 17920 24800 17926 24812
rect 18325 24803 18383 24809
rect 18325 24800 18337 24803
rect 17920 24772 18337 24800
rect 17920 24760 17926 24772
rect 18325 24769 18337 24772
rect 18371 24769 18383 24803
rect 18325 24763 18383 24769
rect 18417 24803 18475 24809
rect 18417 24769 18429 24803
rect 18463 24800 18475 24803
rect 25866 24800 25872 24812
rect 18463 24772 19012 24800
rect 25827 24772 25872 24800
rect 18463 24769 18475 24772
rect 18417 24763 18475 24769
rect 15838 24732 15844 24744
rect 14292 24704 15844 24732
rect 15838 24692 15844 24704
rect 15896 24692 15902 24744
rect 16209 24735 16267 24741
rect 16209 24701 16221 24735
rect 16255 24732 16267 24735
rect 16482 24732 16488 24744
rect 16255 24704 16488 24732
rect 16255 24701 16267 24704
rect 16209 24695 16267 24701
rect 16482 24692 16488 24704
rect 16540 24692 16546 24744
rect 17494 24732 17500 24744
rect 17407 24704 17500 24732
rect 17494 24692 17500 24704
rect 17552 24732 17558 24744
rect 17552 24704 17908 24732
rect 17552 24692 17558 24704
rect 9732 24636 11008 24664
rect 11057 24667 11115 24673
rect 9732 24624 9738 24636
rect 11057 24633 11069 24667
rect 11103 24664 11115 24667
rect 15657 24667 15715 24673
rect 15657 24664 15669 24667
rect 11103 24636 12434 24664
rect 11103 24633 11115 24636
rect 11057 24627 11115 24633
rect 9861 24599 9919 24605
rect 9861 24565 9873 24599
rect 9907 24596 9919 24599
rect 12158 24596 12164 24608
rect 9907 24568 12164 24596
rect 9907 24565 9919 24568
rect 9861 24559 9919 24565
rect 12158 24556 12164 24568
rect 12216 24556 12222 24608
rect 12406 24596 12434 24636
rect 13372 24636 15669 24664
rect 13372 24608 13400 24636
rect 15657 24633 15669 24636
rect 15703 24633 15715 24667
rect 15657 24627 15715 24633
rect 15746 24624 15752 24676
rect 15804 24664 15810 24676
rect 16945 24667 17003 24673
rect 16945 24664 16957 24667
rect 15804 24636 16957 24664
rect 15804 24624 15810 24636
rect 16945 24633 16957 24636
rect 16991 24633 17003 24667
rect 16945 24627 17003 24633
rect 17880 24608 17908 24704
rect 18984 24673 19012 24772
rect 25866 24760 25872 24772
rect 25924 24800 25930 24812
rect 26513 24803 26571 24809
rect 26513 24800 26525 24803
rect 25924 24772 26525 24800
rect 25924 24760 25930 24772
rect 26513 24769 26525 24772
rect 26559 24769 26571 24803
rect 33410 24800 33416 24812
rect 33371 24772 33416 24800
rect 26513 24763 26571 24769
rect 33410 24760 33416 24772
rect 33468 24760 33474 24812
rect 35526 24800 35532 24812
rect 35487 24772 35532 24800
rect 35526 24760 35532 24772
rect 35584 24800 35590 24812
rect 36081 24803 36139 24809
rect 36081 24800 36093 24803
rect 35584 24772 36093 24800
rect 35584 24760 35590 24772
rect 36081 24769 36093 24772
rect 36127 24769 36139 24803
rect 36081 24763 36139 24769
rect 33428 24732 33456 24760
rect 33428 24704 35894 24732
rect 18969 24667 19027 24673
rect 18969 24633 18981 24667
rect 19015 24664 19027 24667
rect 22186 24664 22192 24676
rect 19015 24636 22192 24664
rect 19015 24633 19027 24636
rect 18969 24627 19027 24633
rect 22186 24624 22192 24636
rect 22244 24624 22250 24676
rect 26053 24667 26111 24673
rect 26053 24633 26065 24667
rect 26099 24664 26111 24667
rect 33594 24664 33600 24676
rect 26099 24636 26234 24664
rect 33555 24636 33600 24664
rect 26099 24633 26111 24636
rect 26053 24627 26111 24633
rect 13354 24596 13360 24608
rect 12406 24568 13360 24596
rect 13354 24556 13360 24568
rect 13412 24556 13418 24608
rect 14369 24599 14427 24605
rect 14369 24565 14381 24599
rect 14415 24596 14427 24599
rect 14826 24596 14832 24608
rect 14415 24568 14832 24596
rect 14415 24565 14427 24568
rect 14369 24559 14427 24565
rect 14826 24556 14832 24568
rect 14884 24556 14890 24608
rect 15013 24599 15071 24605
rect 15013 24565 15025 24599
rect 15059 24596 15071 24599
rect 16022 24596 16028 24608
rect 15059 24568 16028 24596
rect 15059 24565 15071 24568
rect 15013 24559 15071 24565
rect 16022 24556 16028 24568
rect 16080 24556 16086 24608
rect 17862 24556 17868 24608
rect 17920 24596 17926 24608
rect 19521 24599 19579 24605
rect 19521 24596 19533 24599
rect 17920 24568 19533 24596
rect 17920 24556 17926 24568
rect 19521 24565 19533 24568
rect 19567 24596 19579 24599
rect 24486 24596 24492 24608
rect 19567 24568 24492 24596
rect 19567 24565 19579 24568
rect 19521 24559 19579 24565
rect 24486 24556 24492 24568
rect 24544 24556 24550 24608
rect 26206 24596 26234 24636
rect 33594 24624 33600 24636
rect 33652 24624 33658 24676
rect 35866 24664 35894 24704
rect 36078 24664 36084 24676
rect 35866 24636 36084 24664
rect 36078 24624 36084 24636
rect 36136 24624 36142 24676
rect 35986 24596 35992 24608
rect 26206 24568 35992 24596
rect 35986 24556 35992 24568
rect 36044 24556 36050 24608
rect 36262 24596 36268 24608
rect 36223 24568 36268 24596
rect 36262 24556 36268 24568
rect 36320 24556 36326 24608
rect 1104 24506 36892 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 36892 24506
rect 1104 24432 36892 24454
rect 11790 24352 11796 24404
rect 11848 24392 11854 24404
rect 12342 24392 12348 24404
rect 11848 24364 12348 24392
rect 11848 24352 11854 24364
rect 12342 24352 12348 24364
rect 12400 24392 12406 24404
rect 15746 24392 15752 24404
rect 12400 24364 15752 24392
rect 12400 24352 12406 24364
rect 15746 24352 15752 24364
rect 15804 24352 15810 24404
rect 16850 24352 16856 24404
rect 16908 24392 16914 24404
rect 17405 24395 17463 24401
rect 17405 24392 17417 24395
rect 16908 24364 17417 24392
rect 16908 24352 16914 24364
rect 17405 24361 17417 24364
rect 17451 24361 17463 24395
rect 17405 24355 17463 24361
rect 17862 24352 17868 24404
rect 17920 24392 17926 24404
rect 17957 24395 18015 24401
rect 17957 24392 17969 24395
rect 17920 24364 17969 24392
rect 17920 24352 17926 24364
rect 17957 24361 17969 24364
rect 18003 24361 18015 24395
rect 17957 24355 18015 24361
rect 26142 24352 26148 24404
rect 26200 24392 26206 24404
rect 28813 24395 28871 24401
rect 28813 24392 28825 24395
rect 26200 24364 28825 24392
rect 26200 24352 26206 24364
rect 28813 24361 28825 24364
rect 28859 24361 28871 24395
rect 28813 24355 28871 24361
rect 9953 24327 10011 24333
rect 9953 24293 9965 24327
rect 9999 24324 10011 24327
rect 12986 24324 12992 24336
rect 9999 24296 12992 24324
rect 9999 24293 10011 24296
rect 9953 24287 10011 24293
rect 12986 24284 12992 24296
rect 13044 24284 13050 24336
rect 13556 24296 22094 24324
rect 11057 24259 11115 24265
rect 11057 24225 11069 24259
rect 11103 24256 11115 24259
rect 11146 24256 11152 24268
rect 11103 24228 11152 24256
rect 11103 24225 11115 24228
rect 11057 24219 11115 24225
rect 11146 24216 11152 24228
rect 11204 24216 11210 24268
rect 11701 24259 11759 24265
rect 11701 24225 11713 24259
rect 11747 24256 11759 24259
rect 11790 24256 11796 24268
rect 11747 24228 11796 24256
rect 11747 24225 11759 24228
rect 11701 24219 11759 24225
rect 11790 24216 11796 24228
rect 11848 24216 11854 24268
rect 12066 24216 12072 24268
rect 12124 24256 12130 24268
rect 12161 24259 12219 24265
rect 12161 24256 12173 24259
rect 12124 24228 12173 24256
rect 12124 24216 12130 24228
rect 12161 24225 12173 24228
rect 12207 24225 12219 24259
rect 12161 24219 12219 24225
rect 12526 24216 12532 24268
rect 12584 24256 12590 24268
rect 13446 24256 13452 24268
rect 12584 24228 13452 24256
rect 12584 24216 12590 24228
rect 13446 24216 13452 24228
rect 13504 24256 13510 24268
rect 13556 24256 13584 24296
rect 13504 24228 13584 24256
rect 13504 24216 13510 24228
rect 12342 24188 12348 24200
rect 12303 24160 12348 24188
rect 12342 24148 12348 24160
rect 12400 24148 12406 24200
rect 13556 24197 13584 24228
rect 13633 24259 13691 24265
rect 13633 24225 13645 24259
rect 13679 24256 13691 24259
rect 14918 24256 14924 24268
rect 13679 24228 14924 24256
rect 13679 24225 13691 24228
rect 13633 24219 13691 24225
rect 14918 24216 14924 24228
rect 14976 24216 14982 24268
rect 15378 24216 15384 24268
rect 15436 24256 15442 24268
rect 15473 24259 15531 24265
rect 15473 24256 15485 24259
rect 15436 24228 15485 24256
rect 15436 24216 15442 24228
rect 15473 24225 15485 24228
rect 15519 24225 15531 24259
rect 15473 24219 15531 24225
rect 15838 24216 15844 24268
rect 15896 24256 15902 24268
rect 18509 24259 18567 24265
rect 18509 24256 18521 24259
rect 15896 24228 16344 24256
rect 15896 24216 15902 24228
rect 13541 24191 13599 24197
rect 13541 24157 13553 24191
rect 13587 24157 13599 24191
rect 13541 24151 13599 24157
rect 7834 24120 7840 24132
rect 7795 24092 7840 24120
rect 7834 24080 7840 24092
rect 7892 24080 7898 24132
rect 8389 24123 8447 24129
rect 8389 24089 8401 24123
rect 8435 24089 8447 24123
rect 8389 24083 8447 24089
rect 6638 24012 6644 24064
rect 6696 24052 6702 24064
rect 8404 24052 8432 24083
rect 8478 24080 8484 24132
rect 8536 24120 8542 24132
rect 8536 24092 8581 24120
rect 8536 24080 8542 24092
rect 8938 24080 8944 24132
rect 8996 24120 9002 24132
rect 9401 24123 9459 24129
rect 9401 24120 9413 24123
rect 8996 24092 9413 24120
rect 8996 24080 9002 24092
rect 9401 24089 9413 24092
rect 9447 24089 9459 24123
rect 9401 24083 9459 24089
rect 9490 24080 9496 24132
rect 9548 24120 9554 24132
rect 11149 24123 11207 24129
rect 9548 24092 9593 24120
rect 9548 24080 9554 24092
rect 11149 24089 11161 24123
rect 11195 24120 11207 24123
rect 11238 24120 11244 24132
rect 11195 24092 11244 24120
rect 11195 24089 11207 24092
rect 11149 24083 11207 24089
rect 11238 24080 11244 24092
rect 11296 24080 11302 24132
rect 11790 24080 11796 24132
rect 11848 24120 11854 24132
rect 11848 24092 13768 24120
rect 11848 24080 11854 24092
rect 12802 24052 12808 24064
rect 6696 24024 8432 24052
rect 12763 24024 12808 24052
rect 6696 24012 6702 24024
rect 12802 24012 12808 24024
rect 12860 24012 12866 24064
rect 13740 24052 13768 24092
rect 14182 24080 14188 24132
rect 14240 24120 14246 24132
rect 14277 24123 14335 24129
rect 14277 24120 14289 24123
rect 14240 24092 14289 24120
rect 14240 24080 14246 24092
rect 14277 24089 14289 24092
rect 14323 24089 14335 24123
rect 14277 24083 14335 24089
rect 14829 24123 14887 24129
rect 14829 24089 14841 24123
rect 14875 24089 14887 24123
rect 16022 24120 16028 24132
rect 15983 24092 16028 24120
rect 14829 24083 14887 24089
rect 14844 24052 14872 24083
rect 16022 24080 16028 24092
rect 16080 24080 16086 24132
rect 16114 24080 16120 24132
rect 16172 24120 16178 24132
rect 16316 24120 16344 24228
rect 16960 24228 18521 24256
rect 16960 24200 16988 24228
rect 18509 24225 18521 24228
rect 18555 24225 18567 24259
rect 22066 24256 22094 24296
rect 25314 24256 25320 24268
rect 22066 24228 25320 24256
rect 18509 24219 18567 24225
rect 25314 24216 25320 24228
rect 25372 24216 25378 24268
rect 16853 24191 16911 24197
rect 16853 24157 16865 24191
rect 16899 24188 16911 24191
rect 16942 24188 16948 24200
rect 16899 24160 16948 24188
rect 16899 24157 16911 24160
rect 16853 24151 16911 24157
rect 16942 24148 16948 24160
rect 17000 24148 17006 24200
rect 17494 24188 17500 24200
rect 17455 24160 17500 24188
rect 17494 24148 17500 24160
rect 17552 24148 17558 24200
rect 28905 24191 28963 24197
rect 28905 24157 28917 24191
rect 28951 24188 28963 24191
rect 33410 24188 33416 24200
rect 28951 24160 33416 24188
rect 28951 24157 28963 24160
rect 28905 24151 28963 24157
rect 33410 24148 33416 24160
rect 33468 24148 33474 24200
rect 17512 24120 17540 24148
rect 16172 24092 16217 24120
rect 16316 24092 17540 24120
rect 16172 24080 16178 24092
rect 13740 24024 14872 24052
rect 15378 24012 15384 24064
rect 15436 24052 15442 24064
rect 16761 24055 16819 24061
rect 16761 24052 16773 24055
rect 15436 24024 16773 24052
rect 15436 24012 15442 24024
rect 16761 24021 16773 24024
rect 16807 24021 16819 24055
rect 16761 24015 16819 24021
rect 1104 23962 36892 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 36892 23962
rect 1104 23888 36892 23910
rect 6641 23851 6699 23857
rect 6641 23817 6653 23851
rect 6687 23848 6699 23851
rect 7926 23848 7932 23860
rect 6687 23820 7932 23848
rect 6687 23817 6699 23820
rect 6641 23811 6699 23817
rect 7926 23808 7932 23820
rect 7984 23808 7990 23860
rect 9861 23851 9919 23857
rect 9861 23817 9873 23851
rect 9907 23848 9919 23851
rect 10870 23848 10876 23860
rect 9907 23820 10876 23848
rect 9907 23817 9919 23820
rect 9861 23811 9919 23817
rect 10870 23808 10876 23820
rect 10928 23808 10934 23860
rect 11057 23851 11115 23857
rect 11057 23817 11069 23851
rect 11103 23848 11115 23851
rect 11790 23848 11796 23860
rect 11103 23820 11796 23848
rect 11103 23817 11115 23820
rect 11057 23811 11115 23817
rect 11790 23808 11796 23820
rect 11848 23808 11854 23860
rect 12342 23848 12348 23860
rect 11900 23820 12348 23848
rect 10413 23783 10471 23789
rect 10413 23749 10425 23783
rect 10459 23780 10471 23783
rect 11900 23780 11928 23820
rect 12342 23808 12348 23820
rect 12400 23808 12406 23860
rect 16114 23808 16120 23860
rect 16172 23848 16178 23860
rect 16853 23851 16911 23857
rect 16853 23848 16865 23851
rect 16172 23820 16865 23848
rect 16172 23808 16178 23820
rect 16853 23817 16865 23820
rect 16899 23817 16911 23851
rect 17494 23848 17500 23860
rect 17455 23820 17500 23848
rect 16853 23811 16911 23817
rect 17494 23808 17500 23820
rect 17552 23808 17558 23860
rect 36081 23851 36139 23857
rect 36081 23817 36093 23851
rect 36127 23848 36139 23851
rect 36170 23848 36176 23860
rect 36127 23820 36176 23848
rect 36127 23817 36139 23820
rect 36081 23811 36139 23817
rect 36170 23808 36176 23820
rect 36228 23808 36234 23860
rect 12250 23780 12256 23792
rect 10459 23752 11928 23780
rect 12211 23752 12256 23780
rect 10459 23749 10471 23752
rect 10413 23743 10471 23749
rect 12250 23740 12256 23752
rect 12308 23740 12314 23792
rect 13170 23780 13176 23792
rect 13131 23752 13176 23780
rect 13170 23740 13176 23752
rect 13228 23740 13234 23792
rect 13814 23780 13820 23792
rect 13775 23752 13820 23780
rect 13814 23740 13820 23752
rect 13872 23740 13878 23792
rect 15378 23780 15384 23792
rect 15339 23752 15384 23780
rect 15378 23740 15384 23752
rect 15436 23740 15442 23792
rect 1854 23712 1860 23724
rect 1815 23684 1860 23712
rect 1854 23672 1860 23684
rect 1912 23672 1918 23724
rect 2498 23712 2504 23724
rect 2459 23684 2504 23712
rect 2498 23672 2504 23684
rect 2556 23672 2562 23724
rect 6546 23712 6552 23724
rect 6459 23684 6552 23712
rect 6546 23672 6552 23684
rect 6604 23712 6610 23724
rect 7193 23715 7251 23721
rect 7193 23712 7205 23715
rect 6604 23684 7205 23712
rect 6604 23672 6610 23684
rect 7193 23681 7205 23684
rect 7239 23681 7251 23715
rect 10318 23712 10324 23724
rect 10231 23684 10324 23712
rect 7193 23675 7251 23681
rect 10318 23672 10324 23684
rect 10376 23712 10382 23724
rect 10686 23712 10692 23724
rect 10376 23684 10692 23712
rect 10376 23672 10382 23684
rect 10686 23672 10692 23684
rect 10744 23672 10750 23724
rect 10870 23672 10876 23724
rect 10928 23712 10934 23724
rect 10965 23715 11023 23721
rect 10965 23712 10977 23715
rect 10928 23684 10977 23712
rect 10928 23672 10934 23684
rect 10965 23681 10977 23684
rect 11011 23712 11023 23715
rect 11974 23712 11980 23724
rect 11011 23684 11980 23712
rect 11011 23681 11023 23684
rect 10965 23675 11023 23681
rect 11974 23672 11980 23684
rect 12032 23672 12038 23724
rect 22186 23672 22192 23724
rect 22244 23712 22250 23724
rect 22373 23715 22431 23721
rect 22373 23712 22385 23715
rect 22244 23684 22385 23712
rect 22244 23672 22250 23684
rect 22373 23681 22385 23684
rect 22419 23681 22431 23715
rect 22373 23675 22431 23681
rect 35894 23672 35900 23724
rect 35952 23712 35958 23724
rect 35952 23684 35997 23712
rect 35952 23672 35958 23684
rect 12161 23647 12219 23653
rect 12161 23613 12173 23647
rect 12207 23644 12219 23647
rect 12802 23644 12808 23656
rect 12207 23616 12808 23644
rect 12207 23613 12219 23616
rect 12161 23607 12219 23613
rect 12802 23604 12808 23616
rect 12860 23604 12866 23656
rect 13722 23644 13728 23656
rect 13683 23616 13728 23644
rect 13722 23604 13728 23616
rect 13780 23604 13786 23656
rect 14001 23647 14059 23653
rect 14001 23613 14013 23647
rect 14047 23644 14059 23647
rect 14182 23644 14188 23656
rect 14047 23616 14188 23644
rect 14047 23613 14059 23616
rect 14001 23607 14059 23613
rect 11698 23536 11704 23588
rect 11756 23576 11762 23588
rect 14016 23576 14044 23607
rect 14182 23604 14188 23616
rect 14240 23604 14246 23656
rect 15289 23647 15347 23653
rect 15289 23613 15301 23647
rect 15335 23644 15347 23647
rect 15378 23644 15384 23656
rect 15335 23616 15384 23644
rect 15335 23613 15347 23616
rect 15289 23607 15347 23613
rect 15378 23604 15384 23616
rect 15436 23604 15442 23656
rect 15470 23604 15476 23656
rect 15528 23644 15534 23656
rect 15565 23647 15623 23653
rect 15565 23644 15577 23647
rect 15528 23616 15577 23644
rect 15528 23604 15534 23616
rect 15565 23613 15577 23616
rect 15611 23613 15623 23647
rect 15565 23607 15623 23613
rect 11756 23548 14044 23576
rect 11756 23536 11762 23548
rect 1670 23508 1676 23520
rect 1631 23480 1676 23508
rect 1670 23468 1676 23480
rect 1728 23468 1734 23520
rect 2314 23508 2320 23520
rect 2275 23480 2320 23508
rect 2314 23468 2320 23480
rect 2372 23468 2378 23520
rect 22465 23511 22523 23517
rect 22465 23477 22477 23511
rect 22511 23508 22523 23511
rect 35434 23508 35440 23520
rect 22511 23480 35440 23508
rect 22511 23477 22523 23480
rect 22465 23471 22523 23477
rect 35434 23468 35440 23480
rect 35492 23468 35498 23520
rect 1104 23418 36892 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 36892 23418
rect 1104 23344 36892 23366
rect 13449 23307 13507 23313
rect 13449 23273 13461 23307
rect 13495 23304 13507 23307
rect 13814 23304 13820 23316
rect 13495 23276 13820 23304
rect 13495 23273 13507 23276
rect 13449 23267 13507 23273
rect 13814 23264 13820 23276
rect 13872 23264 13878 23316
rect 11698 23236 11704 23248
rect 11659 23208 11704 23236
rect 11698 23196 11704 23208
rect 11756 23196 11762 23248
rect 15194 23236 15200 23248
rect 15155 23208 15200 23236
rect 15194 23196 15200 23208
rect 15252 23196 15258 23248
rect 10597 23171 10655 23177
rect 10597 23137 10609 23171
rect 10643 23168 10655 23171
rect 12253 23171 12311 23177
rect 12253 23168 12265 23171
rect 10643 23140 12265 23168
rect 10643 23137 10655 23140
rect 10597 23131 10655 23137
rect 12253 23137 12265 23140
rect 12299 23137 12311 23171
rect 12253 23131 12311 23137
rect 14384 23140 16436 23168
rect 6086 23100 6092 23112
rect 6047 23072 6092 23100
rect 6086 23060 6092 23072
rect 6144 23060 6150 23112
rect 12342 23060 12348 23112
rect 12400 23100 12406 23112
rect 12437 23103 12495 23109
rect 12437 23100 12449 23103
rect 12400 23072 12449 23100
rect 12400 23060 12406 23072
rect 12437 23069 12449 23072
rect 12483 23069 12495 23103
rect 12437 23063 12495 23069
rect 12618 23060 12624 23112
rect 12676 23100 12682 23112
rect 13357 23103 13415 23109
rect 13357 23100 13369 23103
rect 12676 23072 13369 23100
rect 12676 23060 12682 23072
rect 13357 23069 13369 23072
rect 13403 23069 13415 23103
rect 13357 23063 13415 23069
rect 14182 23060 14188 23112
rect 14240 23100 14246 23112
rect 14384 23109 14412 23140
rect 16408 23109 16436 23140
rect 16482 23128 16488 23180
rect 16540 23168 16546 23180
rect 31113 23171 31171 23177
rect 31113 23168 31125 23171
rect 16540 23140 31125 23168
rect 16540 23128 16546 23140
rect 31113 23137 31125 23140
rect 31159 23137 31171 23171
rect 31113 23131 31171 23137
rect 14369 23103 14427 23109
rect 14369 23100 14381 23103
rect 14240 23072 14381 23100
rect 14240 23060 14246 23072
rect 14369 23069 14381 23072
rect 14415 23069 14427 23103
rect 14369 23063 14427 23069
rect 16393 23103 16451 23109
rect 16393 23069 16405 23103
rect 16439 23100 16451 23103
rect 17037 23103 17095 23109
rect 17037 23100 17049 23103
rect 16439 23072 17049 23100
rect 16439 23069 16451 23072
rect 16393 23063 16451 23069
rect 17037 23069 17049 23072
rect 17083 23100 17095 23103
rect 17589 23103 17647 23109
rect 17589 23100 17601 23103
rect 17083 23072 17601 23100
rect 17083 23069 17095 23072
rect 17037 23063 17095 23069
rect 17589 23069 17601 23072
rect 17635 23069 17647 23103
rect 22186 23100 22192 23112
rect 22147 23072 22192 23100
rect 17589 23063 17647 23069
rect 22186 23060 22192 23072
rect 22244 23060 22250 23112
rect 31205 23103 31263 23109
rect 31205 23069 31217 23103
rect 31251 23100 31263 23103
rect 35894 23100 35900 23112
rect 31251 23072 35900 23100
rect 31251 23069 31263 23072
rect 31205 23063 31263 23069
rect 35894 23060 35900 23072
rect 35952 23100 35958 23112
rect 36446 23100 36452 23112
rect 35952 23072 36452 23100
rect 35952 23060 35958 23072
rect 36446 23060 36452 23072
rect 36504 23060 36510 23112
rect 11146 23032 11152 23044
rect 11107 23004 11152 23032
rect 11146 22992 11152 23004
rect 11204 22992 11210 23044
rect 11241 23035 11299 23041
rect 11241 23001 11253 23035
rect 11287 23032 11299 23035
rect 11514 23032 11520 23044
rect 11287 23004 11520 23032
rect 11287 23001 11299 23004
rect 11241 22995 11299 23001
rect 11514 22992 11520 23004
rect 11572 22992 11578 23044
rect 15654 23032 15660 23044
rect 15615 23004 15660 23032
rect 15654 22992 15660 23004
rect 15712 22992 15718 23044
rect 15749 23035 15807 23041
rect 15749 23001 15761 23035
rect 15795 23032 15807 23035
rect 16482 23032 16488 23044
rect 15795 23004 16488 23032
rect 15795 23001 15807 23004
rect 15749 22995 15807 23001
rect 16482 22992 16488 23004
rect 16540 22992 16546 23044
rect 16577 23035 16635 23041
rect 16577 23001 16589 23035
rect 16623 23032 16635 23035
rect 16623 23004 22232 23032
rect 16623 23001 16635 23004
rect 16577 22995 16635 23001
rect 5994 22964 6000 22976
rect 5955 22936 6000 22964
rect 5994 22924 6000 22936
rect 6052 22924 6058 22976
rect 12802 22924 12808 22976
rect 12860 22964 12866 22976
rect 12897 22967 12955 22973
rect 12897 22964 12909 22967
rect 12860 22936 12909 22964
rect 12860 22924 12866 22936
rect 12897 22933 12909 22936
rect 12943 22964 12955 22967
rect 13538 22964 13544 22976
rect 12943 22936 13544 22964
rect 12943 22933 12955 22936
rect 12897 22927 12955 22933
rect 13538 22924 13544 22936
rect 13596 22924 13602 22976
rect 14553 22967 14611 22973
rect 14553 22933 14565 22967
rect 14599 22964 14611 22967
rect 14734 22964 14740 22976
rect 14599 22936 14740 22964
rect 14599 22933 14611 22936
rect 14553 22927 14611 22933
rect 14734 22924 14740 22936
rect 14792 22924 14798 22976
rect 22204 22964 22232 23004
rect 35342 22964 35348 22976
rect 22204 22936 35348 22964
rect 35342 22924 35348 22936
rect 35400 22924 35406 22976
rect 1104 22874 36892 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 36892 22874
rect 1104 22800 36892 22822
rect 1854 22720 1860 22772
rect 1912 22760 1918 22772
rect 1949 22763 2007 22769
rect 1949 22760 1961 22763
rect 1912 22732 1961 22760
rect 1912 22720 1918 22732
rect 1949 22729 1961 22732
rect 1995 22729 2007 22763
rect 1949 22723 2007 22729
rect 8478 22720 8484 22772
rect 8536 22760 8542 22772
rect 12342 22760 12348 22772
rect 8536 22732 11192 22760
rect 12303 22732 12348 22760
rect 8536 22720 8542 22732
rect 8202 22692 8208 22704
rect 8163 22664 8208 22692
rect 8202 22652 8208 22664
rect 8260 22652 8266 22704
rect 9030 22692 9036 22704
rect 8991 22664 9036 22692
rect 9030 22652 9036 22664
rect 9088 22652 9094 22704
rect 9600 22701 9628 22732
rect 9585 22695 9643 22701
rect 9585 22661 9597 22695
rect 9631 22661 9643 22695
rect 10594 22692 10600 22704
rect 10555 22664 10600 22692
rect 9585 22655 9643 22661
rect 10594 22652 10600 22664
rect 10652 22652 10658 22704
rect 11164 22701 11192 22732
rect 12342 22720 12348 22732
rect 12400 22720 12406 22772
rect 12989 22763 13047 22769
rect 12989 22729 13001 22763
rect 13035 22760 13047 22763
rect 15654 22760 15660 22772
rect 13035 22732 15660 22760
rect 13035 22729 13047 22732
rect 12989 22723 13047 22729
rect 15654 22720 15660 22732
rect 15712 22720 15718 22772
rect 11149 22695 11207 22701
rect 11149 22661 11161 22695
rect 11195 22692 11207 22695
rect 11606 22692 11612 22704
rect 11195 22664 11612 22692
rect 11195 22661 11207 22664
rect 11149 22655 11207 22661
rect 11606 22652 11612 22664
rect 11664 22652 11670 22704
rect 13538 22692 13544 22704
rect 13499 22664 13544 22692
rect 13538 22652 13544 22664
rect 13596 22652 13602 22704
rect 14734 22692 14740 22704
rect 14695 22664 14740 22692
rect 14734 22652 14740 22664
rect 14792 22652 14798 22704
rect 14826 22652 14832 22704
rect 14884 22692 14890 22704
rect 15381 22695 15439 22701
rect 14884 22664 14929 22692
rect 14884 22652 14890 22664
rect 15381 22661 15393 22695
rect 15427 22692 15439 22695
rect 15470 22692 15476 22704
rect 15427 22664 15476 22692
rect 15427 22661 15439 22664
rect 15381 22655 15439 22661
rect 15470 22652 15476 22664
rect 15528 22652 15534 22704
rect 2133 22627 2191 22633
rect 2133 22593 2145 22627
rect 2179 22624 2191 22627
rect 2179 22596 2728 22624
rect 2179 22593 2191 22596
rect 2133 22587 2191 22593
rect 2700 22429 2728 22596
rect 11974 22584 11980 22636
rect 12032 22624 12038 22636
rect 12250 22624 12256 22636
rect 12032 22596 12256 22624
rect 12032 22584 12038 22596
rect 12250 22584 12256 22596
rect 12308 22584 12314 22636
rect 12897 22627 12955 22633
rect 12897 22624 12909 22627
rect 12406 22596 12909 22624
rect 7466 22516 7472 22568
rect 7524 22556 7530 22568
rect 7834 22556 7840 22568
rect 7524 22528 7840 22556
rect 7524 22516 7530 22528
rect 7834 22516 7840 22528
rect 7892 22516 7898 22568
rect 8294 22556 8300 22568
rect 8255 22528 8300 22556
rect 8294 22516 8300 22528
rect 8352 22516 8358 22568
rect 8938 22556 8944 22568
rect 8899 22528 8944 22556
rect 8938 22516 8944 22528
rect 8996 22516 9002 22568
rect 10502 22556 10508 22568
rect 10463 22528 10508 22556
rect 10502 22516 10508 22528
rect 10560 22556 10566 22568
rect 10870 22556 10876 22568
rect 10560 22528 10876 22556
rect 10560 22516 10566 22528
rect 10870 22516 10876 22528
rect 10928 22516 10934 22568
rect 8386 22448 8392 22500
rect 8444 22488 8450 22500
rect 11701 22491 11759 22497
rect 11701 22488 11713 22491
rect 8444 22460 11713 22488
rect 8444 22448 8450 22460
rect 11701 22457 11713 22460
rect 11747 22488 11759 22491
rect 12406 22488 12434 22596
rect 12897 22593 12909 22596
rect 12943 22593 12955 22627
rect 12897 22587 12955 22593
rect 14001 22627 14059 22633
rect 14001 22593 14013 22627
rect 14047 22624 14059 22627
rect 16025 22627 16083 22633
rect 14047 22596 14596 22624
rect 14047 22593 14059 22596
rect 14001 22587 14059 22593
rect 14185 22559 14243 22565
rect 14185 22525 14197 22559
rect 14231 22525 14243 22559
rect 14568 22556 14596 22596
rect 16025 22593 16037 22627
rect 16071 22624 16083 22627
rect 16853 22627 16911 22633
rect 16853 22624 16865 22627
rect 16071 22596 16865 22624
rect 16071 22593 16083 22596
rect 16025 22587 16083 22593
rect 16853 22593 16865 22596
rect 16899 22624 16911 22627
rect 18322 22624 18328 22636
rect 16899 22596 18328 22624
rect 16899 22593 16911 22596
rect 16853 22587 16911 22593
rect 15933 22559 15991 22565
rect 15933 22556 15945 22559
rect 14568 22528 15945 22556
rect 14185 22519 14243 22525
rect 15933 22525 15945 22528
rect 15979 22525 15991 22559
rect 15933 22519 15991 22525
rect 11747 22460 12434 22488
rect 14200 22488 14228 22519
rect 15010 22488 15016 22500
rect 14200 22460 15016 22488
rect 11747 22457 11759 22460
rect 11701 22451 11759 22457
rect 15010 22448 15016 22460
rect 15068 22448 15074 22500
rect 2685 22423 2743 22429
rect 2685 22389 2697 22423
rect 2731 22420 2743 22423
rect 3234 22420 3240 22432
rect 2731 22392 3240 22420
rect 2731 22389 2743 22392
rect 2685 22383 2743 22389
rect 3234 22380 3240 22392
rect 3292 22420 3298 22432
rect 6546 22420 6552 22432
rect 3292 22392 6552 22420
rect 3292 22380 3298 22392
rect 6546 22380 6552 22392
rect 6604 22380 6610 22432
rect 12618 22380 12624 22432
rect 12676 22420 12682 22432
rect 16040 22420 16068 22587
rect 18322 22584 18328 22596
rect 18380 22584 18386 22636
rect 36078 22624 36084 22636
rect 36039 22596 36084 22624
rect 36078 22584 36084 22596
rect 36136 22584 36142 22636
rect 36262 22488 36268 22500
rect 36223 22460 36268 22488
rect 36262 22448 36268 22460
rect 36320 22448 36326 22500
rect 12676 22392 16068 22420
rect 12676 22380 12682 22392
rect 1104 22330 36892 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 36892 22330
rect 1104 22256 36892 22278
rect 9030 22176 9036 22228
rect 9088 22216 9094 22228
rect 9217 22219 9275 22225
rect 9217 22216 9229 22219
rect 9088 22188 9229 22216
rect 9088 22176 9094 22188
rect 9217 22185 9229 22188
rect 9263 22185 9275 22219
rect 9217 22179 9275 22185
rect 10594 22176 10600 22228
rect 10652 22216 10658 22228
rect 10873 22219 10931 22225
rect 10873 22216 10885 22219
rect 10652 22188 10885 22216
rect 10652 22176 10658 22188
rect 10873 22185 10885 22188
rect 10919 22185 10931 22219
rect 11514 22216 11520 22228
rect 11475 22188 11520 22216
rect 10873 22179 10931 22185
rect 11514 22176 11520 22188
rect 11572 22176 11578 22228
rect 8294 22108 8300 22160
rect 8352 22148 8358 22160
rect 15194 22148 15200 22160
rect 8352 22120 15200 22148
rect 8352 22108 8358 22120
rect 7009 22083 7067 22089
rect 7009 22049 7021 22083
rect 7055 22080 7067 22083
rect 8938 22080 8944 22092
rect 7055 22052 8944 22080
rect 7055 22049 7067 22052
rect 7009 22043 7067 22049
rect 8938 22040 8944 22052
rect 8996 22040 9002 22092
rect 10318 22040 10324 22092
rect 10376 22080 10382 22092
rect 12621 22083 12679 22089
rect 10376 22052 11468 22080
rect 10376 22040 10382 22052
rect 5721 22015 5779 22021
rect 5721 21981 5733 22015
rect 5767 22012 5779 22015
rect 6917 22015 6975 22021
rect 6917 22012 6929 22015
rect 5767 21984 6929 22012
rect 5767 21981 5779 21984
rect 5721 21975 5779 21981
rect 6288 21888 6316 21984
rect 6917 21981 6929 21984
rect 6963 22012 6975 22015
rect 7561 22015 7619 22021
rect 7561 22012 7573 22015
rect 6963 21984 7573 22012
rect 6963 21981 6975 21984
rect 6917 21975 6975 21981
rect 7561 21981 7573 21984
rect 7607 21981 7619 22015
rect 7561 21975 7619 21981
rect 9309 22015 9367 22021
rect 9309 21981 9321 22015
rect 9355 22012 9367 22015
rect 9398 22012 9404 22024
rect 9355 21984 9404 22012
rect 9355 21981 9367 21984
rect 9309 21975 9367 21981
rect 8573 21947 8631 21953
rect 8573 21913 8585 21947
rect 8619 21944 8631 21947
rect 9324 21944 9352 21975
rect 9398 21972 9404 21984
rect 9456 21972 9462 22024
rect 11440 22021 11468 22052
rect 12621 22049 12633 22083
rect 12667 22080 12679 22083
rect 12710 22080 12716 22092
rect 12667 22052 12716 22080
rect 12667 22049 12679 22052
rect 12621 22043 12679 22049
rect 12710 22040 12716 22052
rect 12768 22040 12774 22092
rect 13633 22083 13691 22089
rect 13633 22049 13645 22083
rect 13679 22080 13691 22083
rect 13998 22080 14004 22092
rect 13679 22052 14004 22080
rect 13679 22049 13691 22052
rect 13633 22043 13691 22049
rect 13998 22040 14004 22052
rect 14056 22040 14062 22092
rect 14844 22089 14872 22120
rect 15194 22108 15200 22120
rect 15252 22108 15258 22160
rect 14829 22083 14887 22089
rect 14829 22049 14841 22083
rect 14875 22049 14887 22083
rect 14829 22043 14887 22049
rect 15286 22040 15292 22092
rect 15344 22080 15350 22092
rect 15344 22052 16252 22080
rect 15344 22040 15350 22052
rect 16224 22024 16252 22052
rect 10965 22015 11023 22021
rect 10965 21981 10977 22015
rect 11011 21981 11023 22015
rect 10965 21975 11023 21981
rect 11425 22015 11483 22021
rect 11425 21981 11437 22015
rect 11471 21981 11483 22015
rect 11425 21975 11483 21981
rect 8619 21916 9352 21944
rect 8619 21913 8631 21916
rect 8573 21907 8631 21913
rect 5902 21876 5908 21888
rect 5863 21848 5908 21876
rect 5902 21836 5908 21848
rect 5960 21836 5966 21888
rect 6270 21836 6276 21888
rect 6328 21876 6334 21888
rect 6365 21879 6423 21885
rect 6365 21876 6377 21879
rect 6328 21848 6377 21876
rect 6328 21836 6334 21848
rect 6365 21845 6377 21848
rect 6411 21845 6423 21879
rect 9324 21876 9352 21916
rect 10321 21947 10379 21953
rect 10321 21913 10333 21947
rect 10367 21944 10379 21947
rect 10980 21944 11008 21975
rect 11974 21972 11980 22024
rect 12032 22012 12038 22024
rect 12529 22015 12587 22021
rect 12529 22012 12541 22015
rect 12032 21984 12541 22012
rect 12032 21972 12038 21984
rect 12529 21981 12541 21984
rect 12575 21981 12587 22015
rect 12529 21975 12587 21981
rect 13725 22015 13783 22021
rect 13725 21981 13737 22015
rect 13771 22012 13783 22015
rect 14090 22012 14096 22024
rect 13771 21984 14096 22012
rect 13771 21981 13783 21984
rect 13725 21975 13783 21981
rect 14090 21972 14096 21984
rect 14148 21972 14154 22024
rect 16206 22012 16212 22024
rect 16119 21984 16212 22012
rect 16206 21972 16212 21984
rect 16264 22012 16270 22024
rect 16669 22015 16727 22021
rect 16669 22012 16681 22015
rect 16264 21984 16681 22012
rect 16264 21972 16270 21984
rect 16669 21981 16681 21984
rect 16715 21981 16727 22015
rect 16669 21975 16727 21981
rect 31941 22015 31999 22021
rect 31941 21981 31953 22015
rect 31987 22012 31999 22015
rect 31987 21984 32536 22012
rect 31987 21981 31999 21984
rect 31941 21975 31999 21981
rect 13906 21944 13912 21956
rect 10367 21916 13912 21944
rect 10367 21913 10379 21916
rect 10321 21907 10379 21913
rect 13906 21904 13912 21916
rect 13964 21904 13970 21956
rect 15286 21944 15292 21956
rect 14016 21916 15292 21944
rect 14016 21876 14044 21916
rect 15286 21904 15292 21916
rect 15344 21904 15350 21956
rect 15381 21947 15439 21953
rect 15381 21913 15393 21947
rect 15427 21913 15439 21947
rect 15381 21907 15439 21913
rect 15473 21947 15531 21953
rect 15473 21913 15485 21947
rect 15519 21944 15531 21947
rect 30558 21944 30564 21956
rect 15519 21916 30564 21944
rect 15519 21913 15531 21916
rect 15473 21907 15531 21913
rect 9324 21848 14044 21876
rect 6365 21839 6423 21845
rect 14090 21836 14096 21888
rect 14148 21876 14154 21888
rect 14277 21879 14335 21885
rect 14277 21876 14289 21879
rect 14148 21848 14289 21876
rect 14148 21836 14154 21848
rect 14277 21845 14289 21848
rect 14323 21845 14335 21879
rect 15396 21876 15424 21907
rect 30558 21904 30564 21916
rect 30616 21904 30622 21956
rect 16117 21879 16175 21885
rect 16117 21876 16129 21879
rect 15396 21848 16129 21876
rect 14277 21839 14335 21845
rect 16117 21845 16129 21848
rect 16163 21845 16175 21879
rect 31754 21876 31760 21888
rect 31715 21848 31760 21876
rect 16117 21839 16175 21845
rect 31754 21836 31760 21848
rect 31812 21836 31818 21888
rect 32508 21885 32536 21984
rect 32493 21879 32551 21885
rect 32493 21845 32505 21879
rect 32539 21876 32551 21879
rect 35894 21876 35900 21888
rect 32539 21848 35900 21876
rect 32539 21845 32551 21848
rect 32493 21839 32551 21845
rect 35894 21836 35900 21848
rect 35952 21836 35958 21888
rect 1104 21786 36892 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 36892 21786
rect 1104 21712 36892 21734
rect 12618 21672 12624 21684
rect 12579 21644 12624 21672
rect 12618 21632 12624 21644
rect 12676 21632 12682 21684
rect 13265 21675 13323 21681
rect 13265 21641 13277 21675
rect 13311 21672 13323 21675
rect 13722 21672 13728 21684
rect 13311 21644 13728 21672
rect 13311 21641 13323 21644
rect 13265 21635 13323 21641
rect 13722 21632 13728 21644
rect 13780 21632 13786 21684
rect 27154 21672 27160 21684
rect 13832 21644 27160 21672
rect 7282 21564 7288 21616
rect 7340 21604 7346 21616
rect 7929 21607 7987 21613
rect 7929 21604 7941 21607
rect 7340 21576 7941 21604
rect 7340 21564 7346 21576
rect 7929 21573 7941 21576
rect 7975 21573 7987 21607
rect 7929 21567 7987 21573
rect 11974 21564 11980 21616
rect 12032 21604 12038 21616
rect 13832 21604 13860 21644
rect 27154 21632 27160 21644
rect 27212 21632 27218 21684
rect 12032 21576 13860 21604
rect 13909 21607 13967 21613
rect 12032 21564 12038 21576
rect 13909 21573 13921 21607
rect 13955 21604 13967 21607
rect 15657 21607 15715 21613
rect 15657 21604 15669 21607
rect 13955 21576 15669 21604
rect 13955 21573 13967 21576
rect 13909 21567 13967 21573
rect 15657 21573 15669 21576
rect 15703 21573 15715 21607
rect 15657 21567 15715 21573
rect 1857 21539 1915 21545
rect 1857 21505 1869 21539
rect 1903 21536 1915 21539
rect 2314 21536 2320 21548
rect 1903 21508 2320 21536
rect 1903 21505 1915 21508
rect 1857 21499 1915 21505
rect 2314 21496 2320 21508
rect 2372 21496 2378 21548
rect 12986 21496 12992 21548
rect 13044 21536 13050 21548
rect 13357 21539 13415 21545
rect 13357 21536 13369 21539
rect 13044 21508 13369 21536
rect 13044 21496 13050 21508
rect 13357 21505 13369 21508
rect 13403 21505 13415 21539
rect 13814 21536 13820 21548
rect 13775 21508 13820 21536
rect 13357 21499 13415 21505
rect 13814 21496 13820 21508
rect 13872 21496 13878 21548
rect 35986 21496 35992 21548
rect 36044 21536 36050 21548
rect 36081 21539 36139 21545
rect 36081 21536 36093 21539
rect 36044 21508 36093 21536
rect 36044 21496 36050 21508
rect 36081 21505 36093 21508
rect 36127 21505 36139 21539
rect 36081 21499 36139 21505
rect 7282 21428 7288 21480
rect 7340 21468 7346 21480
rect 7377 21471 7435 21477
rect 7377 21468 7389 21471
rect 7340 21440 7389 21468
rect 7340 21428 7346 21440
rect 7377 21437 7389 21440
rect 7423 21437 7435 21471
rect 7377 21431 7435 21437
rect 8021 21471 8079 21477
rect 8021 21437 8033 21471
rect 8067 21468 8079 21471
rect 8202 21468 8208 21480
rect 8067 21440 8208 21468
rect 8067 21437 8079 21440
rect 8021 21431 8079 21437
rect 8202 21428 8208 21440
rect 8260 21428 8266 21480
rect 14645 21471 14703 21477
rect 14645 21437 14657 21471
rect 14691 21468 14703 21471
rect 14734 21468 14740 21480
rect 14691 21440 14740 21468
rect 14691 21437 14703 21440
rect 14645 21431 14703 21437
rect 14734 21428 14740 21440
rect 14792 21428 14798 21480
rect 15746 21468 15752 21480
rect 15707 21440 15752 21468
rect 15746 21428 15752 21440
rect 15804 21428 15810 21480
rect 15194 21400 15200 21412
rect 15155 21372 15200 21400
rect 15194 21360 15200 21372
rect 15252 21360 15258 21412
rect 1670 21332 1676 21344
rect 1631 21304 1676 21332
rect 1670 21292 1676 21304
rect 1728 21292 1734 21344
rect 11974 21292 11980 21344
rect 12032 21332 12038 21344
rect 12069 21335 12127 21341
rect 12069 21332 12081 21335
rect 12032 21304 12081 21332
rect 12032 21292 12038 21304
rect 12069 21301 12081 21304
rect 12115 21301 12127 21335
rect 36262 21332 36268 21344
rect 36223 21304 36268 21332
rect 12069 21295 12127 21301
rect 36262 21292 36268 21304
rect 36320 21292 36326 21344
rect 1104 21242 36892 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 36892 21242
rect 1104 21168 36892 21190
rect 12161 21131 12219 21137
rect 12161 21097 12173 21131
rect 12207 21128 12219 21131
rect 12250 21128 12256 21140
rect 12207 21100 12256 21128
rect 12207 21097 12219 21100
rect 12161 21091 12219 21097
rect 12250 21088 12256 21100
rect 12308 21088 12314 21140
rect 12986 21088 12992 21140
rect 13044 21128 13050 21140
rect 25406 21128 25412 21140
rect 13044 21100 25412 21128
rect 13044 21088 13050 21100
rect 25406 21088 25412 21100
rect 25464 21088 25470 21140
rect 30558 21128 30564 21140
rect 30519 21100 30564 21128
rect 30558 21088 30564 21100
rect 30616 21088 30622 21140
rect 36078 21128 36084 21140
rect 36039 21100 36084 21128
rect 36078 21088 36084 21100
rect 36136 21088 36142 21140
rect 13725 21063 13783 21069
rect 13725 21029 13737 21063
rect 13771 21060 13783 21063
rect 13814 21060 13820 21072
rect 13771 21032 13820 21060
rect 13771 21029 13783 21032
rect 13725 21023 13783 21029
rect 13814 21020 13820 21032
rect 13872 21020 13878 21072
rect 14734 20992 14740 21004
rect 14695 20964 14740 20992
rect 14734 20952 14740 20964
rect 14792 20952 14798 21004
rect 30653 20927 30711 20933
rect 30653 20893 30665 20927
rect 30699 20924 30711 20927
rect 31205 20927 31263 20933
rect 31205 20924 31217 20927
rect 30699 20896 31217 20924
rect 30699 20893 30711 20896
rect 30653 20887 30711 20893
rect 31205 20893 31217 20896
rect 31251 20924 31263 20927
rect 35437 20927 35495 20933
rect 35437 20924 35449 20927
rect 31251 20896 35449 20924
rect 31251 20893 31263 20896
rect 31205 20887 31263 20893
rect 35437 20893 35449 20896
rect 35483 20924 35495 20927
rect 35710 20924 35716 20936
rect 35483 20896 35716 20924
rect 35483 20893 35495 20896
rect 35437 20887 35495 20893
rect 35710 20884 35716 20896
rect 35768 20924 35774 20936
rect 35897 20927 35955 20933
rect 35897 20924 35909 20927
rect 35768 20896 35909 20924
rect 35768 20884 35774 20896
rect 35897 20893 35909 20896
rect 35943 20893 35955 20927
rect 35897 20887 35955 20893
rect 14826 20856 14832 20868
rect 14787 20828 14832 20856
rect 14826 20816 14832 20828
rect 14884 20816 14890 20868
rect 15381 20859 15439 20865
rect 15381 20825 15393 20859
rect 15427 20856 15439 20859
rect 16390 20856 16396 20868
rect 15427 20828 16396 20856
rect 15427 20825 15439 20828
rect 15381 20819 15439 20825
rect 16390 20816 16396 20828
rect 16448 20816 16454 20868
rect 12986 20788 12992 20800
rect 12947 20760 12992 20788
rect 12986 20748 12992 20760
rect 13044 20748 13050 20800
rect 1104 20698 36892 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 36892 20698
rect 1104 20624 36892 20646
rect 14369 20587 14427 20593
rect 14369 20553 14381 20587
rect 14415 20584 14427 20587
rect 14826 20584 14832 20596
rect 14415 20556 14832 20584
rect 14415 20553 14427 20556
rect 14369 20547 14427 20553
rect 14826 20544 14832 20556
rect 14884 20544 14890 20596
rect 16206 20584 16212 20596
rect 16167 20556 16212 20584
rect 16206 20544 16212 20556
rect 16264 20544 16270 20596
rect 13814 20408 13820 20460
rect 13872 20448 13878 20460
rect 14277 20451 14335 20457
rect 14277 20448 14289 20451
rect 13872 20420 14289 20448
rect 13872 20408 13878 20420
rect 14277 20417 14289 20420
rect 14323 20448 14335 20451
rect 14921 20451 14979 20457
rect 14921 20448 14933 20451
rect 14323 20420 14933 20448
rect 14323 20417 14335 20420
rect 14277 20411 14335 20417
rect 14921 20417 14933 20420
rect 14967 20417 14979 20451
rect 14921 20411 14979 20417
rect 15565 20451 15623 20457
rect 15565 20417 15577 20451
rect 15611 20448 15623 20451
rect 16224 20448 16252 20544
rect 15611 20420 16252 20448
rect 15611 20417 15623 20420
rect 15565 20411 15623 20417
rect 15657 20315 15715 20321
rect 15657 20281 15669 20315
rect 15703 20312 15715 20315
rect 16942 20312 16948 20324
rect 15703 20284 16948 20312
rect 15703 20281 15715 20284
rect 15657 20275 15715 20281
rect 16942 20272 16948 20284
rect 17000 20272 17006 20324
rect 1104 20154 36892 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 36892 20154
rect 1104 20080 36892 20102
rect 3053 20043 3111 20049
rect 3053 20040 3065 20043
rect 2746 20012 3065 20040
rect 1857 19839 1915 19845
rect 1857 19805 1869 19839
rect 1903 19805 1915 19839
rect 1857 19799 1915 19805
rect 2501 19839 2559 19845
rect 2501 19805 2513 19839
rect 2547 19836 2559 19839
rect 2746 19836 2774 20012
rect 3053 20009 3065 20012
rect 3099 20040 3111 20043
rect 5258 20040 5264 20052
rect 3099 20012 5264 20040
rect 3099 20009 3111 20012
rect 3053 20003 3111 20009
rect 5258 20000 5264 20012
rect 5316 20000 5322 20052
rect 8205 20043 8263 20049
rect 8205 20009 8217 20043
rect 8251 20040 8263 20043
rect 8386 20040 8392 20052
rect 8251 20012 8392 20040
rect 8251 20009 8263 20012
rect 8205 20003 8263 20009
rect 2547 19808 2774 19836
rect 7653 19839 7711 19845
rect 2547 19805 2559 19808
rect 2501 19799 2559 19805
rect 7653 19805 7665 19839
rect 7699 19836 7711 19839
rect 8220 19836 8248 20003
rect 8386 20000 8392 20012
rect 8444 20000 8450 20052
rect 9217 20043 9275 20049
rect 9217 20009 9229 20043
rect 9263 20040 9275 20043
rect 11146 20040 11152 20052
rect 9263 20012 11152 20040
rect 9263 20009 9275 20012
rect 9217 20003 9275 20009
rect 11146 20000 11152 20012
rect 11204 20000 11210 20052
rect 21818 20040 21824 20052
rect 21779 20012 21824 20040
rect 21818 20000 21824 20012
rect 21876 20000 21882 20052
rect 7699 19808 8248 19836
rect 9125 19839 9183 19845
rect 7699 19805 7711 19808
rect 7653 19799 7711 19805
rect 9125 19805 9137 19839
rect 9171 19836 9183 19839
rect 9769 19839 9827 19845
rect 9769 19836 9781 19839
rect 9171 19808 9781 19836
rect 9171 19805 9183 19808
rect 9125 19799 9183 19805
rect 9769 19805 9781 19808
rect 9815 19805 9827 19839
rect 9769 19799 9827 19805
rect 21361 19839 21419 19845
rect 21361 19805 21373 19839
rect 21407 19836 21419 19839
rect 21818 19836 21824 19848
rect 21407 19808 21824 19836
rect 21407 19805 21419 19808
rect 21361 19799 21419 19805
rect 1872 19768 1900 19799
rect 5994 19768 6000 19780
rect 1872 19740 6000 19768
rect 5994 19728 6000 19740
rect 6052 19728 6058 19780
rect 6178 19728 6184 19780
rect 6236 19768 6242 19780
rect 9140 19768 9168 19799
rect 21818 19796 21824 19808
rect 21876 19796 21882 19848
rect 6236 19740 9168 19768
rect 6236 19728 6242 19740
rect 1670 19700 1676 19712
rect 1631 19672 1676 19700
rect 1670 19660 1676 19672
rect 1728 19660 1734 19712
rect 1946 19660 1952 19712
rect 2004 19700 2010 19712
rect 2317 19703 2375 19709
rect 2317 19700 2329 19703
rect 2004 19672 2329 19700
rect 2004 19660 2010 19672
rect 2317 19669 2329 19672
rect 2363 19669 2375 19703
rect 7558 19700 7564 19712
rect 7519 19672 7564 19700
rect 2317 19663 2375 19669
rect 7558 19660 7564 19672
rect 7616 19660 7622 19712
rect 20806 19660 20812 19712
rect 20864 19700 20870 19712
rect 21177 19703 21235 19709
rect 21177 19700 21189 19703
rect 20864 19672 21189 19700
rect 20864 19660 20870 19672
rect 21177 19669 21189 19672
rect 21223 19669 21235 19703
rect 21177 19663 21235 19669
rect 1104 19610 36892 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 36892 19610
rect 1104 19536 36892 19558
rect 1104 19066 36892 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 36892 19066
rect 1104 18992 36892 19014
rect 2498 18816 2504 18828
rect 2459 18788 2504 18816
rect 2498 18776 2504 18788
rect 2556 18776 2562 18828
rect 8113 18819 8171 18825
rect 8113 18785 8125 18819
rect 8159 18816 8171 18819
rect 8202 18816 8208 18828
rect 8159 18788 8208 18816
rect 8159 18785 8171 18788
rect 8113 18779 8171 18785
rect 8202 18776 8208 18788
rect 8260 18816 8266 18828
rect 16390 18816 16396 18828
rect 8260 18788 16396 18816
rect 8260 18776 8266 18788
rect 16390 18776 16396 18788
rect 16448 18776 16454 18828
rect 1949 18751 2007 18757
rect 1949 18717 1961 18751
rect 1995 18748 2007 18751
rect 2516 18748 2544 18776
rect 1995 18720 2544 18748
rect 1995 18717 2007 18720
rect 1949 18711 2007 18717
rect 7469 18683 7527 18689
rect 7469 18680 7481 18683
rect 7392 18652 7481 18680
rect 7392 18624 7420 18652
rect 7469 18649 7481 18652
rect 7515 18649 7527 18683
rect 7469 18643 7527 18649
rect 7558 18640 7564 18692
rect 7616 18680 7622 18692
rect 16942 18680 16948 18692
rect 7616 18652 7661 18680
rect 16903 18652 16948 18680
rect 7616 18640 7622 18652
rect 16942 18640 16948 18652
rect 17000 18640 17006 18692
rect 17037 18683 17095 18689
rect 17037 18649 17049 18683
rect 17083 18680 17095 18683
rect 17083 18652 17724 18680
rect 17083 18649 17095 18652
rect 17037 18643 17095 18649
rect 17696 18624 17724 18652
rect 1762 18612 1768 18624
rect 1723 18584 1768 18612
rect 1762 18572 1768 18584
rect 1820 18572 1826 18624
rect 7374 18572 7380 18624
rect 7432 18572 7438 18624
rect 17678 18612 17684 18624
rect 17639 18584 17684 18612
rect 17678 18572 17684 18584
rect 17736 18572 17742 18624
rect 1104 18522 36892 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 36892 18522
rect 1104 18448 36892 18470
rect 1578 18232 1584 18284
rect 1636 18272 1642 18284
rect 1673 18275 1731 18281
rect 1673 18272 1685 18275
rect 1636 18244 1685 18272
rect 1636 18232 1642 18244
rect 1673 18241 1685 18244
rect 1719 18241 1731 18275
rect 1673 18235 1731 18241
rect 1765 18071 1823 18077
rect 1765 18037 1777 18071
rect 1811 18068 1823 18071
rect 12986 18068 12992 18080
rect 1811 18040 12992 18068
rect 1811 18037 1823 18040
rect 1765 18031 1823 18037
rect 12986 18028 12992 18040
rect 13044 18028 13050 18080
rect 1104 17978 36892 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 36892 17978
rect 1104 17904 36892 17926
rect 1578 17796 1584 17808
rect 1539 17768 1584 17796
rect 1578 17756 1584 17768
rect 1636 17756 1642 17808
rect 1104 17434 36892 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 36892 17434
rect 1104 17360 36892 17382
rect 27341 17323 27399 17329
rect 27341 17289 27353 17323
rect 27387 17320 27399 17323
rect 27387 17292 35894 17320
rect 27387 17289 27399 17292
rect 27341 17283 27399 17289
rect 27154 17184 27160 17196
rect 27115 17156 27160 17184
rect 27154 17144 27160 17156
rect 27212 17184 27218 17196
rect 27801 17187 27859 17193
rect 27801 17184 27813 17187
rect 27212 17156 27813 17184
rect 27212 17144 27218 17156
rect 27801 17153 27813 17156
rect 27847 17153 27859 17187
rect 35866 17184 35894 17292
rect 36081 17187 36139 17193
rect 36081 17184 36093 17187
rect 35866 17156 36093 17184
rect 27801 17147 27859 17153
rect 36081 17153 36093 17156
rect 36127 17153 36139 17187
rect 36081 17147 36139 17153
rect 36262 17048 36268 17060
rect 36223 17020 36268 17048
rect 36262 17008 36268 17020
rect 36320 17008 36326 17060
rect 1104 16890 36892 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 36892 16890
rect 1104 16816 36892 16838
rect 1104 16346 36892 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 36892 16346
rect 1104 16272 36892 16294
rect 1857 16099 1915 16105
rect 1857 16065 1869 16099
rect 1903 16096 1915 16099
rect 13817 16099 13875 16105
rect 1903 16068 2774 16096
rect 1903 16065 1915 16068
rect 1857 16059 1915 16065
rect 2746 15960 2774 16068
rect 13817 16065 13829 16099
rect 13863 16096 13875 16099
rect 14090 16096 14096 16108
rect 13863 16068 14096 16096
rect 13863 16065 13875 16068
rect 13817 16059 13875 16065
rect 14090 16056 14096 16068
rect 14148 16096 14154 16108
rect 25406 16096 25412 16108
rect 14148 16068 14412 16096
rect 25319 16068 25412 16096
rect 14148 16056 14154 16068
rect 14384 15969 14412 16068
rect 25406 16056 25412 16068
rect 25464 16096 25470 16108
rect 26053 16099 26111 16105
rect 26053 16096 26065 16099
rect 25464 16068 26065 16096
rect 25464 16056 25470 16068
rect 26053 16065 26065 16068
rect 26099 16065 26111 16099
rect 26053 16059 26111 16065
rect 36081 16099 36139 16105
rect 36081 16065 36093 16099
rect 36127 16096 36139 16099
rect 36170 16096 36176 16108
rect 36127 16068 36176 16096
rect 36127 16065 36139 16068
rect 36081 16059 36139 16065
rect 36170 16056 36176 16068
rect 36228 16056 36234 16108
rect 36354 16028 36360 16040
rect 36315 16000 36360 16028
rect 36354 15988 36360 16000
rect 36412 15988 36418 16040
rect 13633 15963 13691 15969
rect 13633 15960 13645 15963
rect 2746 15932 13645 15960
rect 13633 15929 13645 15932
rect 13679 15929 13691 15963
rect 13633 15923 13691 15929
rect 14369 15963 14427 15969
rect 14369 15929 14381 15963
rect 14415 15960 14427 15963
rect 34146 15960 34152 15972
rect 14415 15932 34152 15960
rect 14415 15929 14427 15932
rect 14369 15923 14427 15929
rect 34146 15920 34152 15932
rect 34204 15920 34210 15972
rect 1670 15892 1676 15904
rect 1631 15864 1676 15892
rect 1670 15852 1676 15864
rect 1728 15852 1734 15904
rect 25590 15892 25596 15904
rect 25551 15864 25596 15892
rect 25590 15852 25596 15864
rect 25648 15852 25654 15904
rect 1104 15802 36892 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 36892 15802
rect 1104 15728 36892 15750
rect 25590 15648 25596 15700
rect 25648 15688 25654 15700
rect 34514 15688 34520 15700
rect 25648 15660 34520 15688
rect 25648 15648 25654 15660
rect 34514 15648 34520 15660
rect 34572 15648 34578 15700
rect 36354 15688 36360 15700
rect 36315 15660 36360 15688
rect 36354 15648 36360 15660
rect 36412 15648 36418 15700
rect 1104 15258 36892 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 36892 15258
rect 1104 15184 36892 15206
rect 1104 14714 36892 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 36892 14714
rect 1104 14640 36892 14662
rect 24854 14396 24860 14408
rect 24815 14368 24860 14396
rect 24854 14356 24860 14368
rect 24912 14396 24918 14408
rect 25501 14399 25559 14405
rect 25501 14396 25513 14399
rect 24912 14368 25513 14396
rect 24912 14356 24918 14368
rect 25501 14365 25513 14368
rect 25547 14365 25559 14399
rect 25501 14359 25559 14365
rect 31389 14399 31447 14405
rect 31389 14365 31401 14399
rect 31435 14396 31447 14399
rect 36170 14396 36176 14408
rect 31435 14368 36176 14396
rect 31435 14365 31447 14368
rect 31389 14359 31447 14365
rect 36170 14356 36176 14368
rect 36228 14356 36234 14408
rect 1670 14328 1676 14340
rect 1631 14300 1676 14328
rect 1670 14288 1676 14300
rect 1728 14288 1734 14340
rect 1857 14331 1915 14337
rect 1857 14297 1869 14331
rect 1903 14328 1915 14331
rect 6178 14328 6184 14340
rect 1903 14300 6184 14328
rect 1903 14297 1915 14300
rect 1857 14291 1915 14297
rect 6178 14288 6184 14300
rect 6236 14288 6242 14340
rect 17678 14288 17684 14340
rect 17736 14328 17742 14340
rect 31297 14331 31355 14337
rect 31297 14328 31309 14331
rect 17736 14300 31309 14328
rect 17736 14288 17742 14300
rect 31297 14297 31309 14300
rect 31343 14297 31355 14331
rect 31297 14291 31355 14297
rect 25038 14260 25044 14272
rect 24999 14232 25044 14260
rect 25038 14220 25044 14232
rect 25096 14220 25102 14272
rect 1104 14170 36892 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 36892 14170
rect 1104 14096 36892 14118
rect 1670 14056 1676 14068
rect 1631 14028 1676 14056
rect 1670 14016 1676 14028
rect 1728 14016 1734 14068
rect 13078 14016 13084 14068
rect 13136 14056 13142 14068
rect 13173 14059 13231 14065
rect 13173 14056 13185 14059
rect 13136 14028 13185 14056
rect 13136 14016 13142 14028
rect 13173 14025 13185 14028
rect 13219 14025 13231 14059
rect 13173 14019 13231 14025
rect 13357 13923 13415 13929
rect 13357 13889 13369 13923
rect 13403 13920 13415 13923
rect 13446 13920 13452 13932
rect 13403 13892 13452 13920
rect 13403 13889 13415 13892
rect 13357 13883 13415 13889
rect 13446 13880 13452 13892
rect 13504 13920 13510 13932
rect 13817 13923 13875 13929
rect 13817 13920 13829 13923
rect 13504 13892 13829 13920
rect 13504 13880 13510 13892
rect 13817 13889 13829 13892
rect 13863 13889 13875 13923
rect 13817 13883 13875 13889
rect 34514 13880 34520 13932
rect 34572 13920 34578 13932
rect 36081 13923 36139 13929
rect 36081 13920 36093 13923
rect 34572 13892 36093 13920
rect 34572 13880 34578 13892
rect 36081 13889 36093 13892
rect 36127 13889 36139 13923
rect 36081 13883 36139 13889
rect 36262 13716 36268 13728
rect 36223 13688 36268 13716
rect 36262 13676 36268 13688
rect 36320 13676 36326 13728
rect 1104 13626 36892 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 36892 13626
rect 1104 13552 36892 13574
rect 1949 13311 2007 13317
rect 1949 13277 1961 13311
rect 1995 13308 2007 13311
rect 7282 13308 7288 13320
rect 1995 13280 7288 13308
rect 1995 13277 2007 13280
rect 1949 13271 2007 13277
rect 7282 13268 7288 13280
rect 7340 13268 7346 13320
rect 1854 13172 1860 13184
rect 1815 13144 1860 13172
rect 1854 13132 1860 13144
rect 1912 13132 1918 13184
rect 1104 13082 36892 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 36892 13082
rect 1104 13008 36892 13030
rect 1854 12832 1860 12844
rect 1815 12804 1860 12832
rect 1854 12792 1860 12804
rect 1912 12792 1918 12844
rect 1670 12628 1676 12640
rect 1631 12600 1676 12628
rect 1670 12588 1676 12600
rect 1728 12588 1734 12640
rect 1104 12538 36892 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 36892 12538
rect 1104 12464 36892 12486
rect 1104 11994 36892 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 36892 11994
rect 1104 11920 36892 11942
rect 35713 11747 35771 11753
rect 35713 11713 35725 11747
rect 35759 11744 35771 11747
rect 36354 11744 36360 11756
rect 35759 11716 36360 11744
rect 35759 11713 35771 11716
rect 35713 11707 35771 11713
rect 36354 11704 36360 11716
rect 36412 11704 36418 11756
rect 36170 11540 36176 11552
rect 36131 11512 36176 11540
rect 36170 11500 36176 11512
rect 36228 11500 36234 11552
rect 1104 11450 36892 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 36892 11450
rect 1104 11376 36892 11398
rect 1104 10906 36892 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 36892 10906
rect 1104 10832 36892 10854
rect 1857 10659 1915 10665
rect 1857 10625 1869 10659
rect 1903 10656 1915 10659
rect 1946 10656 1952 10668
rect 1903 10628 1952 10656
rect 1903 10625 1915 10628
rect 1857 10619 1915 10625
rect 1946 10616 1952 10628
rect 2004 10616 2010 10668
rect 36081 10659 36139 10665
rect 36081 10625 36093 10659
rect 36127 10656 36139 10659
rect 36446 10656 36452 10668
rect 36127 10628 36452 10656
rect 36127 10625 36139 10628
rect 36081 10619 36139 10625
rect 36446 10616 36452 10628
rect 36504 10616 36510 10668
rect 36354 10588 36360 10600
rect 36315 10560 36360 10588
rect 36354 10548 36360 10560
rect 36412 10548 36418 10600
rect 1670 10452 1676 10464
rect 1631 10424 1676 10452
rect 1670 10412 1676 10424
rect 1728 10412 1734 10464
rect 1104 10362 36892 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 36892 10362
rect 1104 10288 36892 10310
rect 36354 10248 36360 10260
rect 36315 10220 36360 10248
rect 36354 10208 36360 10220
rect 36412 10208 36418 10260
rect 1104 9818 36892 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 36892 9818
rect 1104 9744 36892 9766
rect 5353 9639 5411 9645
rect 5353 9605 5365 9639
rect 5399 9636 5411 9639
rect 7374 9636 7380 9648
rect 5399 9608 7380 9636
rect 5399 9605 5411 9608
rect 5353 9599 5411 9605
rect 7374 9596 7380 9608
rect 7432 9596 7438 9648
rect 2774 9528 2780 9580
rect 2832 9568 2838 9580
rect 5261 9571 5319 9577
rect 5261 9568 5273 9571
rect 2832 9540 5273 9568
rect 2832 9528 2838 9540
rect 5261 9537 5273 9540
rect 5307 9537 5319 9571
rect 35989 9571 36047 9577
rect 35989 9568 36001 9571
rect 5261 9531 5319 9537
rect 35866 9540 36001 9568
rect 13170 9324 13176 9376
rect 13228 9364 13234 9376
rect 35437 9367 35495 9373
rect 35437 9364 35449 9367
rect 13228 9336 35449 9364
rect 13228 9324 13234 9336
rect 35437 9333 35449 9336
rect 35483 9364 35495 9367
rect 35866 9364 35894 9540
rect 35989 9537 36001 9540
rect 36035 9537 36047 9571
rect 35989 9531 36047 9537
rect 36078 9364 36084 9376
rect 35483 9336 35894 9364
rect 36039 9336 36084 9364
rect 35483 9333 35495 9336
rect 35437 9327 35495 9333
rect 36078 9324 36084 9336
rect 36136 9324 36142 9376
rect 1104 9274 36892 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 36892 9274
rect 1104 9200 36892 9222
rect 1857 9027 1915 9033
rect 1857 8993 1869 9027
rect 1903 9024 1915 9027
rect 6270 9024 6276 9036
rect 1903 8996 6276 9024
rect 1903 8993 1915 8996
rect 1857 8987 1915 8993
rect 6270 8984 6276 8996
rect 6328 8984 6334 9036
rect 1578 8956 1584 8968
rect 1539 8928 1584 8956
rect 1578 8916 1584 8928
rect 1636 8916 1642 8968
rect 1104 8730 36892 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 36892 8730
rect 1104 8656 36892 8678
rect 1578 8616 1584 8628
rect 1539 8588 1584 8616
rect 1578 8576 1584 8588
rect 1636 8576 1642 8628
rect 10870 8616 10876 8628
rect 10831 8588 10876 8616
rect 10870 8576 10876 8588
rect 10928 8576 10934 8628
rect 15197 8619 15255 8625
rect 15197 8585 15209 8619
rect 15243 8616 15255 8619
rect 15378 8616 15384 8628
rect 15243 8588 15384 8616
rect 15243 8585 15255 8588
rect 15197 8579 15255 8585
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 24486 8616 24492 8628
rect 24447 8588 24492 8616
rect 24486 8576 24492 8588
rect 24544 8576 24550 8628
rect 36170 8548 36176 8560
rect 35866 8520 36176 8548
rect 10962 8480 10968 8492
rect 10923 8452 10968 8480
rect 10962 8440 10968 8452
rect 11020 8440 11026 8492
rect 15102 8480 15108 8492
rect 15063 8452 15108 8480
rect 15102 8440 15108 8452
rect 15160 8480 15166 8492
rect 15749 8483 15807 8489
rect 15749 8480 15761 8483
rect 15160 8452 15761 8480
rect 15160 8440 15166 8452
rect 15749 8449 15761 8452
rect 15795 8449 15807 8483
rect 15749 8443 15807 8449
rect 24581 8483 24639 8489
rect 24581 8449 24593 8483
rect 24627 8480 24639 8483
rect 30006 8480 30012 8492
rect 24627 8452 30012 8480
rect 24627 8449 24639 8452
rect 24581 8443 24639 8449
rect 30006 8440 30012 8452
rect 30064 8440 30070 8492
rect 35437 8483 35495 8489
rect 35437 8449 35449 8483
rect 35483 8480 35495 8483
rect 35866 8480 35894 8520
rect 36170 8508 36176 8520
rect 36228 8508 36234 8560
rect 36078 8480 36084 8492
rect 35483 8452 35894 8480
rect 36039 8452 36084 8480
rect 35483 8449 35495 8452
rect 35437 8443 35495 8449
rect 36078 8440 36084 8452
rect 36136 8440 36142 8492
rect 35621 8347 35679 8353
rect 35621 8313 35633 8347
rect 35667 8344 35679 8347
rect 36078 8344 36084 8356
rect 35667 8316 36084 8344
rect 35667 8313 35679 8316
rect 35621 8307 35679 8313
rect 36078 8304 36084 8316
rect 36136 8304 36142 8356
rect 36262 8344 36268 8356
rect 36223 8316 36268 8344
rect 36262 8304 36268 8316
rect 36320 8304 36326 8356
rect 1104 8186 36892 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 36892 8186
rect 1104 8112 36892 8134
rect 15746 8072 15752 8084
rect 15707 8044 15752 8072
rect 15746 8032 15752 8044
rect 15804 8032 15810 8084
rect 15838 7868 15844 7880
rect 15799 7840 15844 7868
rect 15838 7828 15844 7840
rect 15896 7828 15902 7880
rect 1104 7642 36892 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 36892 7642
rect 1104 7568 36892 7590
rect 1854 7392 1860 7404
rect 1815 7364 1860 7392
rect 1854 7352 1860 7364
rect 1912 7352 1918 7404
rect 1670 7188 1676 7200
rect 1631 7160 1676 7188
rect 1670 7148 1676 7160
rect 1728 7148 1734 7200
rect 1104 7098 36892 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 36892 7098
rect 1104 7024 36892 7046
rect 6362 6780 6368 6792
rect 6323 6752 6368 6780
rect 6362 6740 6368 6752
rect 6420 6780 6426 6792
rect 7009 6783 7067 6789
rect 7009 6780 7021 6783
rect 6420 6752 7021 6780
rect 6420 6740 6426 6752
rect 7009 6749 7021 6752
rect 7055 6749 7067 6783
rect 7009 6743 7067 6749
rect 6546 6644 6552 6656
rect 6507 6616 6552 6644
rect 6546 6604 6552 6616
rect 6604 6604 6610 6656
rect 1104 6554 36892 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 36892 6554
rect 1104 6480 36892 6502
rect 15010 6440 15016 6452
rect 14971 6412 15016 6440
rect 15010 6400 15016 6412
rect 15068 6400 15074 6452
rect 35894 6400 35900 6452
rect 35952 6440 35958 6452
rect 36173 6443 36231 6449
rect 36173 6440 36185 6443
rect 35952 6412 36185 6440
rect 35952 6400 35958 6412
rect 36173 6409 36185 6412
rect 36219 6409 36231 6443
rect 36173 6403 36231 6409
rect 15105 6307 15163 6313
rect 15105 6273 15117 6307
rect 15151 6304 15163 6307
rect 15562 6304 15568 6316
rect 15151 6276 15568 6304
rect 15151 6273 15163 6276
rect 15105 6267 15163 6273
rect 15562 6264 15568 6276
rect 15620 6264 15626 6316
rect 35713 6307 35771 6313
rect 35713 6273 35725 6307
rect 35759 6304 35771 6307
rect 36354 6304 36360 6316
rect 35759 6276 36360 6304
rect 35759 6273 35771 6276
rect 35713 6267 35771 6273
rect 36354 6264 36360 6276
rect 36412 6264 36418 6316
rect 1104 6010 36892 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 36892 6010
rect 1104 5936 36892 5958
rect 1104 5466 36892 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 36892 5466
rect 1104 5392 36892 5414
rect 1578 5216 1584 5228
rect 1539 5188 1584 5216
rect 1578 5176 1584 5188
rect 1636 5216 1642 5228
rect 2225 5219 2283 5225
rect 2225 5216 2237 5219
rect 1636 5188 2237 5216
rect 1636 5176 1642 5188
rect 2225 5185 2237 5188
rect 2271 5185 2283 5219
rect 36078 5216 36084 5228
rect 36039 5188 36084 5216
rect 2225 5179 2283 5185
rect 36078 5176 36084 5188
rect 36136 5176 36142 5228
rect 1765 5015 1823 5021
rect 1765 4981 1777 5015
rect 1811 5012 1823 5015
rect 2774 5012 2780 5024
rect 1811 4984 2780 5012
rect 1811 4981 1823 4984
rect 1765 4975 1823 4981
rect 2774 4972 2780 4984
rect 2832 5012 2838 5024
rect 3970 5012 3976 5024
rect 2832 4984 3976 5012
rect 2832 4972 2838 4984
rect 3970 4972 3976 4984
rect 4028 4972 4034 5024
rect 36262 5012 36268 5024
rect 36223 4984 36268 5012
rect 36262 4972 36268 4984
rect 36320 4972 36326 5024
rect 1104 4922 36892 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 36892 4922
rect 1104 4848 36892 4870
rect 1104 4378 36892 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 36892 4378
rect 1104 4304 36892 4326
rect 36354 3924 36360 3936
rect 36315 3896 36360 3924
rect 36354 3884 36360 3896
rect 36412 3884 36418 3936
rect 1104 3834 36892 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 36892 3834
rect 1104 3760 36892 3782
rect 1854 3680 1860 3732
rect 1912 3720 1918 3732
rect 2317 3723 2375 3729
rect 2317 3720 2329 3723
rect 1912 3692 2329 3720
rect 1912 3680 1918 3692
rect 2317 3689 2329 3692
rect 2363 3689 2375 3723
rect 15562 3720 15568 3732
rect 15523 3692 15568 3720
rect 2317 3683 2375 3689
rect 15562 3680 15568 3692
rect 15620 3680 15626 3732
rect 1857 3519 1915 3525
rect 1857 3485 1869 3519
rect 1903 3485 1915 3519
rect 2498 3516 2504 3528
rect 2459 3488 2504 3516
rect 1857 3479 1915 3485
rect 1872 3448 1900 3479
rect 2498 3476 2504 3488
rect 2556 3476 2562 3528
rect 15105 3519 15163 3525
rect 15105 3485 15117 3519
rect 15151 3516 15163 3519
rect 15562 3516 15568 3528
rect 15151 3488 15568 3516
rect 15151 3485 15163 3488
rect 15105 3479 15163 3485
rect 15562 3476 15568 3488
rect 15620 3516 15626 3528
rect 36081 3519 36139 3525
rect 36081 3516 36093 3519
rect 15620 3488 16574 3516
rect 15620 3476 15626 3488
rect 11698 3448 11704 3460
rect 1872 3420 11704 3448
rect 11698 3408 11704 3420
rect 11756 3408 11762 3460
rect 16546 3448 16574 3488
rect 35866 3488 36093 3516
rect 34882 3448 34888 3460
rect 16546 3420 34888 3448
rect 34882 3408 34888 3420
rect 34940 3408 34946 3460
rect 1670 3380 1676 3392
rect 1631 3352 1676 3380
rect 1670 3340 1676 3352
rect 1728 3340 1734 3392
rect 14918 3380 14924 3392
rect 14879 3352 14924 3380
rect 14918 3340 14924 3352
rect 14976 3340 14982 3392
rect 33134 3340 33140 3392
rect 33192 3380 33198 3392
rect 35529 3383 35587 3389
rect 35529 3380 35541 3383
rect 33192 3352 35541 3380
rect 33192 3340 33198 3352
rect 35529 3349 35541 3352
rect 35575 3380 35587 3383
rect 35866 3380 35894 3488
rect 36081 3485 36093 3488
rect 36127 3485 36139 3519
rect 36081 3479 36139 3485
rect 36262 3380 36268 3392
rect 35575 3352 35894 3380
rect 36223 3352 36268 3380
rect 35575 3349 35587 3352
rect 35529 3343 35587 3349
rect 36262 3340 36268 3352
rect 36320 3340 36326 3392
rect 1104 3290 36892 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 36892 3290
rect 1104 3216 36892 3238
rect 11698 3176 11704 3188
rect 11659 3148 11704 3176
rect 11698 3136 11704 3148
rect 11756 3136 11762 3188
rect 12437 3179 12495 3185
rect 12437 3176 12449 3179
rect 12360 3148 12449 3176
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3009 1915 3043
rect 3970 3040 3976 3052
rect 3931 3012 3976 3040
rect 1857 3003 1915 3009
rect 1872 2972 1900 3003
rect 3970 3000 3976 3012
rect 4028 3000 4034 3052
rect 11885 3043 11943 3049
rect 11885 3009 11897 3043
rect 11931 3040 11943 3043
rect 12360 3040 12388 3148
rect 12437 3145 12449 3148
rect 12483 3176 12495 3179
rect 15102 3176 15108 3188
rect 12483 3148 15108 3176
rect 12483 3145 12495 3148
rect 12437 3139 12495 3145
rect 15102 3136 15108 3148
rect 15160 3136 15166 3188
rect 14458 3108 14464 3120
rect 14419 3080 14464 3108
rect 14458 3068 14464 3080
rect 14516 3068 14522 3120
rect 17126 3068 17132 3120
rect 17184 3108 17190 3120
rect 23661 3111 23719 3117
rect 23661 3108 23673 3111
rect 17184 3080 23673 3108
rect 17184 3068 17190 3080
rect 15838 3040 15844 3052
rect 11931 3012 12388 3040
rect 15799 3012 15844 3040
rect 11931 3009 11943 3012
rect 11885 3003 11943 3009
rect 15838 3000 15844 3012
rect 15896 3000 15902 3052
rect 19334 3040 19340 3052
rect 19295 3012 19340 3040
rect 19334 3000 19340 3012
rect 19392 3040 19398 3052
rect 23032 3049 23060 3080
rect 23661 3077 23673 3080
rect 23707 3077 23719 3111
rect 23661 3071 23719 3077
rect 19981 3043 20039 3049
rect 19981 3040 19993 3043
rect 19392 3012 19993 3040
rect 19392 3000 19398 3012
rect 19981 3009 19993 3012
rect 20027 3009 20039 3043
rect 19981 3003 20039 3009
rect 23017 3043 23075 3049
rect 23017 3009 23029 3043
rect 23063 3009 23075 3043
rect 23017 3003 23075 3009
rect 30006 3000 30012 3052
rect 30064 3040 30070 3052
rect 33045 3043 33103 3049
rect 33045 3040 33057 3043
rect 30064 3012 33057 3040
rect 30064 3000 30070 3012
rect 33045 3009 33057 3012
rect 33091 3009 33103 3043
rect 34793 3043 34851 3049
rect 34793 3040 34805 3043
rect 33045 3003 33103 3009
rect 33244 3012 34805 3040
rect 14918 2972 14924 2984
rect 1872 2944 14924 2972
rect 14918 2932 14924 2944
rect 14976 2932 14982 2984
rect 23109 2975 23167 2981
rect 23109 2941 23121 2975
rect 23155 2972 23167 2975
rect 24670 2972 24676 2984
rect 23155 2944 24676 2972
rect 23155 2941 23167 2944
rect 23109 2935 23167 2941
rect 24670 2932 24676 2944
rect 24728 2932 24734 2984
rect 10962 2864 10968 2916
rect 11020 2904 11026 2916
rect 14458 2904 14464 2916
rect 11020 2876 14464 2904
rect 11020 2864 11026 2876
rect 14458 2864 14464 2876
rect 14516 2864 14522 2916
rect 14645 2907 14703 2913
rect 14645 2873 14657 2907
rect 14691 2904 14703 2907
rect 33134 2904 33140 2916
rect 14691 2876 33140 2904
rect 14691 2873 14703 2876
rect 14645 2867 14703 2873
rect 33134 2864 33140 2876
rect 33192 2864 33198 2916
rect 33244 2913 33272 3012
rect 34793 3009 34805 3012
rect 34839 3009 34851 3043
rect 34793 3003 34851 3009
rect 34882 3000 34888 3052
rect 34940 3040 34946 3052
rect 36081 3043 36139 3049
rect 36081 3040 36093 3043
rect 34940 3012 36093 3040
rect 34940 3000 34946 3012
rect 36081 3009 36093 3012
rect 36127 3009 36139 3043
rect 36081 3003 36139 3009
rect 36354 2972 36360 2984
rect 36267 2944 36360 2972
rect 36354 2932 36360 2944
rect 36412 2972 36418 2984
rect 37366 2972 37372 2984
rect 36412 2944 37372 2972
rect 36412 2932 36418 2944
rect 37366 2932 37372 2944
rect 37424 2932 37430 2984
rect 33229 2907 33287 2913
rect 33229 2873 33241 2907
rect 33275 2873 33287 2907
rect 33229 2867 33287 2873
rect 1670 2836 1676 2848
rect 1631 2808 1676 2836
rect 1670 2796 1676 2808
rect 1728 2796 1734 2848
rect 2314 2836 2320 2848
rect 2275 2808 2320 2836
rect 2314 2796 2320 2808
rect 2372 2796 2378 2848
rect 4157 2839 4215 2845
rect 4157 2805 4169 2839
rect 4203 2836 4215 2839
rect 4614 2836 4620 2848
rect 4203 2808 4620 2836
rect 4203 2805 4215 2808
rect 4157 2799 4215 2805
rect 4614 2796 4620 2808
rect 4672 2796 4678 2848
rect 10226 2836 10232 2848
rect 10187 2808 10232 2836
rect 10226 2796 10232 2808
rect 10284 2796 10290 2848
rect 15194 2796 15200 2848
rect 15252 2836 15258 2848
rect 15657 2839 15715 2845
rect 15657 2836 15669 2839
rect 15252 2808 15669 2836
rect 15252 2796 15258 2808
rect 15657 2805 15669 2808
rect 15703 2805 15715 2839
rect 15657 2799 15715 2805
rect 19429 2839 19487 2845
rect 19429 2805 19441 2839
rect 19475 2836 19487 2839
rect 22002 2836 22008 2848
rect 19475 2808 22008 2836
rect 19475 2805 19487 2808
rect 19429 2799 19487 2805
rect 22002 2796 22008 2808
rect 22060 2796 22066 2848
rect 32214 2796 32220 2848
rect 32272 2836 32278 2848
rect 32309 2839 32367 2845
rect 32309 2836 32321 2839
rect 32272 2808 32321 2836
rect 32272 2796 32278 2808
rect 32309 2805 32321 2808
rect 32355 2805 32367 2839
rect 32309 2799 32367 2805
rect 34977 2839 35035 2845
rect 34977 2805 34989 2839
rect 35023 2836 35035 2839
rect 36538 2836 36544 2848
rect 35023 2808 36544 2836
rect 35023 2805 35035 2808
rect 34977 2799 35035 2805
rect 36538 2796 36544 2808
rect 36596 2796 36602 2848
rect 1104 2746 36892 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 36892 2746
rect 1104 2672 36892 2694
rect 2498 2632 2504 2644
rect 2459 2604 2504 2632
rect 2498 2592 2504 2604
rect 2556 2592 2562 2644
rect 3234 2632 3240 2644
rect 3195 2604 3240 2632
rect 3234 2592 3240 2604
rect 3292 2592 3298 2644
rect 11054 2592 11060 2644
rect 11112 2632 11118 2644
rect 11112 2604 15240 2632
rect 11112 2592 11118 2604
rect 10689 2567 10747 2573
rect 10689 2533 10701 2567
rect 10735 2564 10747 2567
rect 11974 2564 11980 2576
rect 10735 2536 11980 2564
rect 10735 2533 10747 2536
rect 10689 2527 10747 2533
rect 11974 2524 11980 2536
rect 12032 2524 12038 2576
rect 13725 2567 13783 2573
rect 13725 2533 13737 2567
rect 13771 2564 13783 2567
rect 14182 2564 14188 2576
rect 13771 2536 14188 2564
rect 13771 2533 13783 2536
rect 13725 2527 13783 2533
rect 14182 2524 14188 2536
rect 14240 2524 14246 2576
rect 15212 2564 15240 2604
rect 15838 2592 15844 2644
rect 15896 2632 15902 2644
rect 19429 2635 19487 2641
rect 19429 2632 19441 2635
rect 15896 2604 19441 2632
rect 15896 2592 15902 2604
rect 19429 2601 19441 2604
rect 19475 2601 19487 2635
rect 20806 2632 20812 2644
rect 20767 2604 20812 2632
rect 19429 2595 19487 2601
rect 20806 2592 20812 2604
rect 20864 2592 20870 2644
rect 22186 2632 22192 2644
rect 22147 2604 22192 2632
rect 22186 2592 22192 2604
rect 22244 2592 22250 2644
rect 25038 2592 25044 2644
rect 25096 2632 25102 2644
rect 32398 2632 32404 2644
rect 25096 2604 31064 2632
rect 32359 2604 32404 2632
rect 25096 2592 25102 2604
rect 16209 2567 16267 2573
rect 16209 2564 16221 2567
rect 15212 2536 16221 2564
rect 16209 2533 16221 2536
rect 16255 2533 16267 2567
rect 16209 2527 16267 2533
rect 9401 2499 9459 2505
rect 9401 2465 9413 2499
rect 9447 2496 9459 2499
rect 10962 2496 10968 2508
rect 9447 2468 10968 2496
rect 9447 2465 9459 2468
rect 9401 2459 9459 2465
rect 10962 2456 10968 2468
rect 11020 2456 11026 2508
rect 1762 2388 1768 2440
rect 1820 2428 1826 2440
rect 1857 2431 1915 2437
rect 1857 2428 1869 2431
rect 1820 2400 1869 2428
rect 1820 2388 1826 2400
rect 1857 2397 1869 2400
rect 1903 2397 1915 2431
rect 2314 2428 2320 2440
rect 2275 2400 2320 2428
rect 1857 2391 1915 2397
rect 2314 2388 2320 2400
rect 2372 2388 2378 2440
rect 4614 2428 4620 2440
rect 4575 2400 4620 2428
rect 4614 2388 4620 2400
rect 4672 2388 4678 2440
rect 6546 2428 6552 2440
rect 6507 2400 6552 2428
rect 6546 2388 6552 2400
rect 6604 2388 6610 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 8496 2400 9137 2428
rect 3234 2320 3240 2372
rect 3292 2360 3298 2372
rect 3329 2363 3387 2369
rect 3329 2360 3341 2363
rect 3292 2332 3341 2360
rect 3292 2320 3298 2332
rect 3329 2329 3341 2332
rect 3375 2360 3387 2363
rect 3973 2363 4031 2369
rect 3973 2360 3985 2363
rect 3375 2332 3985 2360
rect 3375 2329 3387 2332
rect 3329 2323 3387 2329
rect 3973 2329 3985 2332
rect 4019 2329 4031 2363
rect 3973 2323 4031 2329
rect 1302 2252 1308 2304
rect 1360 2292 1366 2304
rect 1673 2295 1731 2301
rect 1673 2292 1685 2295
rect 1360 2264 1685 2292
rect 1360 2252 1366 2264
rect 1673 2261 1685 2264
rect 1719 2261 1731 2295
rect 1673 2255 1731 2261
rect 4522 2252 4528 2304
rect 4580 2292 4586 2304
rect 4801 2295 4859 2301
rect 4801 2292 4813 2295
rect 4580 2264 4813 2292
rect 4580 2252 4586 2264
rect 4801 2261 4813 2264
rect 4847 2261 4859 2295
rect 4801 2255 4859 2261
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 6733 2295 6791 2301
rect 6733 2292 6745 2295
rect 6512 2264 6745 2292
rect 6512 2252 6518 2264
rect 6733 2261 6745 2264
rect 6779 2261 6791 2295
rect 6733 2255 6791 2261
rect 8386 2252 8392 2304
rect 8444 2292 8450 2304
rect 8496 2301 8524 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 11977 2431 12035 2437
rect 11977 2397 11989 2431
rect 12023 2428 12035 2431
rect 13078 2428 13084 2440
rect 12023 2400 13084 2428
rect 12023 2397 12035 2400
rect 11977 2391 12035 2397
rect 13078 2388 13084 2400
rect 13136 2388 13142 2440
rect 15194 2428 15200 2440
rect 15155 2400 15200 2428
rect 15194 2388 15200 2400
rect 15252 2388 15258 2440
rect 16224 2428 16252 2527
rect 22002 2524 22008 2576
rect 22060 2564 22066 2576
rect 22060 2536 25912 2564
rect 22060 2524 22066 2536
rect 24857 2499 24915 2505
rect 24857 2496 24869 2499
rect 16960 2468 24869 2496
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16224 2400 16865 2428
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 9674 2320 9680 2372
rect 9732 2360 9738 2372
rect 10226 2360 10232 2372
rect 9732 2332 10232 2360
rect 9732 2320 9738 2332
rect 10226 2320 10232 2332
rect 10284 2360 10290 2372
rect 10505 2363 10563 2369
rect 10505 2360 10517 2363
rect 10284 2332 10517 2360
rect 10284 2320 10290 2332
rect 10505 2329 10517 2332
rect 10551 2329 10563 2363
rect 13538 2360 13544 2372
rect 13499 2332 13544 2360
rect 10505 2323 10563 2329
rect 13538 2320 13544 2332
rect 13596 2360 13602 2372
rect 14277 2363 14335 2369
rect 14277 2360 14289 2363
rect 13596 2332 14289 2360
rect 13596 2320 13602 2332
rect 14277 2329 14289 2332
rect 14323 2329 14335 2363
rect 14277 2323 14335 2329
rect 15102 2320 15108 2372
rect 15160 2360 15166 2372
rect 16960 2360 16988 2468
rect 24857 2465 24869 2468
rect 24903 2465 24915 2499
rect 24857 2459 24915 2465
rect 19613 2431 19671 2437
rect 19613 2428 19625 2431
rect 15160 2332 16988 2360
rect 18800 2400 19625 2428
rect 15160 2320 15166 2332
rect 8481 2295 8539 2301
rect 8481 2292 8493 2295
rect 8444 2264 8493 2292
rect 8444 2252 8450 2264
rect 8481 2261 8493 2264
rect 8527 2261 8539 2295
rect 8481 2255 8539 2261
rect 11606 2252 11612 2304
rect 11664 2292 11670 2304
rect 11793 2295 11851 2301
rect 11793 2292 11805 2295
rect 11664 2264 11805 2292
rect 11664 2252 11670 2264
rect 11793 2261 11805 2264
rect 11839 2261 11851 2295
rect 11793 2255 11851 2261
rect 14826 2252 14832 2304
rect 14884 2292 14890 2304
rect 15013 2295 15071 2301
rect 15013 2292 15025 2295
rect 14884 2264 15025 2292
rect 14884 2252 14890 2264
rect 15013 2261 15025 2264
rect 15059 2261 15071 2295
rect 15013 2255 15071 2261
rect 16758 2252 16764 2304
rect 16816 2292 16822 2304
rect 17037 2295 17095 2301
rect 17037 2292 17049 2295
rect 16816 2264 17049 2292
rect 16816 2252 16822 2264
rect 17037 2261 17049 2264
rect 17083 2261 17095 2295
rect 17037 2255 17095 2261
rect 18690 2252 18696 2304
rect 18748 2292 18754 2304
rect 18800 2301 18828 2400
rect 19613 2397 19625 2400
rect 19659 2397 19671 2431
rect 19613 2391 19671 2397
rect 20349 2431 20407 2437
rect 20349 2397 20361 2431
rect 20395 2428 20407 2431
rect 20806 2428 20812 2440
rect 20395 2400 20812 2428
rect 20395 2397 20407 2400
rect 20349 2391 20407 2397
rect 20806 2388 20812 2400
rect 20864 2388 20870 2440
rect 25884 2437 25912 2536
rect 30006 2496 30012 2508
rect 29967 2468 30012 2496
rect 30006 2456 30012 2468
rect 30064 2456 30070 2508
rect 31036 2437 31064 2604
rect 32398 2592 32404 2604
rect 32456 2592 32462 2644
rect 34146 2632 34152 2644
rect 34107 2604 34152 2632
rect 34146 2592 34152 2604
rect 34204 2592 34210 2644
rect 35710 2456 35716 2508
rect 35768 2496 35774 2508
rect 35805 2499 35863 2505
rect 35805 2496 35817 2499
rect 35768 2468 35817 2496
rect 35768 2456 35774 2468
rect 35805 2465 35817 2468
rect 35851 2465 35863 2499
rect 35805 2459 35863 2465
rect 24581 2431 24639 2437
rect 24581 2428 24593 2431
rect 23952 2400 24593 2428
rect 21453 2363 21511 2369
rect 21453 2329 21465 2363
rect 21499 2360 21511 2363
rect 21910 2360 21916 2372
rect 21499 2332 21916 2360
rect 21499 2329 21511 2332
rect 21453 2323 21511 2329
rect 21910 2320 21916 2332
rect 21968 2360 21974 2372
rect 22097 2363 22155 2369
rect 22097 2360 22109 2363
rect 21968 2332 22109 2360
rect 21968 2320 21974 2332
rect 22097 2329 22109 2332
rect 22143 2329 22155 2363
rect 22097 2323 22155 2329
rect 18785 2295 18843 2301
rect 18785 2292 18797 2295
rect 18748 2264 18797 2292
rect 18748 2252 18754 2264
rect 18785 2261 18797 2264
rect 18831 2261 18843 2295
rect 18785 2255 18843 2261
rect 19978 2252 19984 2304
rect 20036 2292 20042 2304
rect 20165 2295 20223 2301
rect 20165 2292 20177 2295
rect 20036 2264 20177 2292
rect 20036 2252 20042 2264
rect 20165 2261 20177 2264
rect 20211 2261 20223 2295
rect 20165 2255 20223 2261
rect 23842 2252 23848 2304
rect 23900 2292 23906 2304
rect 23952 2301 23980 2400
rect 24581 2397 24593 2400
rect 24627 2397 24639 2431
rect 24581 2391 24639 2397
rect 25869 2431 25927 2437
rect 25869 2397 25881 2431
rect 25915 2397 25927 2431
rect 27157 2431 27215 2437
rect 27157 2428 27169 2431
rect 25869 2391 25927 2397
rect 26206 2400 27169 2428
rect 24670 2320 24676 2372
rect 24728 2360 24734 2372
rect 26206 2360 26234 2400
rect 27157 2397 27169 2400
rect 27203 2397 27215 2431
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 27157 2391 27215 2397
rect 29104 2400 29745 2428
rect 24728 2332 26234 2360
rect 24728 2320 24734 2332
rect 23937 2295 23995 2301
rect 23937 2292 23949 2295
rect 23900 2264 23949 2292
rect 23900 2252 23906 2264
rect 23937 2261 23949 2264
rect 23983 2261 23995 2295
rect 23937 2255 23995 2261
rect 25130 2252 25136 2304
rect 25188 2292 25194 2304
rect 26053 2295 26111 2301
rect 26053 2292 26065 2295
rect 25188 2264 26065 2292
rect 25188 2252 25194 2264
rect 26053 2261 26065 2264
rect 26099 2261 26111 2295
rect 26053 2255 26111 2261
rect 27062 2252 27068 2304
rect 27120 2292 27126 2304
rect 27341 2295 27399 2301
rect 27341 2292 27353 2295
rect 27120 2264 27353 2292
rect 27120 2252 27126 2264
rect 27341 2261 27353 2264
rect 27387 2261 27399 2295
rect 27341 2255 27399 2261
rect 28994 2252 29000 2304
rect 29052 2292 29058 2304
rect 29104 2301 29132 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 31021 2431 31079 2437
rect 31021 2397 31033 2431
rect 31067 2397 31079 2431
rect 31021 2391 31079 2397
rect 33597 2431 33655 2437
rect 33597 2397 33609 2431
rect 33643 2428 33655 2431
rect 35434 2428 35440 2440
rect 33643 2400 35440 2428
rect 33643 2397 33655 2400
rect 33597 2391 33655 2397
rect 35434 2388 35440 2400
rect 35492 2428 35498 2440
rect 35529 2431 35587 2437
rect 35529 2428 35541 2431
rect 35492 2400 35541 2428
rect 35492 2388 35498 2400
rect 35529 2397 35541 2400
rect 35575 2397 35587 2431
rect 35529 2391 35587 2397
rect 32214 2320 32220 2372
rect 32272 2360 32278 2372
rect 32493 2363 32551 2369
rect 32493 2360 32505 2363
rect 32272 2332 32505 2360
rect 32272 2320 32278 2332
rect 32493 2329 32505 2332
rect 32539 2329 32551 2363
rect 32493 2323 32551 2329
rect 34146 2320 34152 2372
rect 34204 2360 34210 2372
rect 34241 2363 34299 2369
rect 34241 2360 34253 2363
rect 34204 2332 34253 2360
rect 34204 2320 34210 2332
rect 34241 2329 34253 2332
rect 34287 2360 34299 2363
rect 34885 2363 34943 2369
rect 34885 2360 34897 2363
rect 34287 2332 34897 2360
rect 34287 2329 34299 2332
rect 34241 2323 34299 2329
rect 34885 2329 34897 2332
rect 34931 2329 34943 2363
rect 34885 2323 34943 2329
rect 29089 2295 29147 2301
rect 29089 2292 29101 2295
rect 29052 2264 29101 2292
rect 29052 2252 29058 2264
rect 29089 2261 29101 2264
rect 29135 2261 29147 2295
rect 29089 2255 29147 2261
rect 30282 2252 30288 2304
rect 30340 2292 30346 2304
rect 31205 2295 31263 2301
rect 31205 2292 31217 2295
rect 30340 2264 31217 2292
rect 30340 2252 30346 2264
rect 31205 2261 31217 2264
rect 31251 2261 31263 2295
rect 31205 2255 31263 2261
rect 1104 2202 36892 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 36892 2202
rect 1104 2128 36892 2150
rect 14 1300 20 1352
rect 72 1340 78 1352
rect 2314 1340 2320 1352
rect 72 1312 2320 1340
rect 72 1300 78 1312
rect 2314 1300 2320 1312
rect 2372 1300 2378 1352
<< via1 >>
rect 664 37612 716 37664
rect 5172 37612 5224 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 3424 37272 3476 37324
rect 4528 37272 4580 37324
rect 25136 37408 25188 37460
rect 35440 37408 35492 37460
rect 9312 37272 9364 37324
rect 10600 37315 10652 37324
rect 10600 37281 10609 37315
rect 10609 37281 10643 37315
rect 10643 37281 10652 37315
rect 10600 37272 10652 37281
rect 1768 37136 1820 37188
rect 3148 37136 3200 37188
rect 5632 37204 5684 37256
rect 1584 37068 1636 37120
rect 2596 37068 2648 37120
rect 3332 37111 3384 37120
rect 3332 37077 3341 37111
rect 3341 37077 3375 37111
rect 3375 37077 3384 37111
rect 10876 37247 10928 37256
rect 10876 37213 10885 37247
rect 10885 37213 10919 37247
rect 10919 37213 10928 37247
rect 11704 37247 11756 37256
rect 10876 37204 10928 37213
rect 11704 37213 11713 37247
rect 11713 37213 11747 37247
rect 11747 37213 11756 37247
rect 11704 37204 11756 37213
rect 12900 37204 12952 37256
rect 14832 37204 14884 37256
rect 30288 37272 30340 37324
rect 16580 37204 16632 37256
rect 18144 37247 18196 37256
rect 18144 37213 18153 37247
rect 18153 37213 18187 37247
rect 18187 37213 18196 37247
rect 18144 37204 18196 37213
rect 18788 37204 18840 37256
rect 22008 37247 22060 37256
rect 22008 37213 22017 37247
rect 22017 37213 22051 37247
rect 22051 37213 22060 37247
rect 22008 37204 22060 37213
rect 23480 37247 23532 37256
rect 23480 37213 23489 37247
rect 23489 37213 23523 37247
rect 23523 37213 23532 37247
rect 23480 37204 23532 37213
rect 25136 37204 25188 37256
rect 28448 37247 28500 37256
rect 7840 37136 7892 37188
rect 8576 37136 8628 37188
rect 3332 37068 3384 37077
rect 6644 37068 6696 37120
rect 8300 37111 8352 37120
rect 8300 37077 8309 37111
rect 8309 37077 8343 37111
rect 8343 37077 8352 37111
rect 8300 37068 8352 37077
rect 8668 37068 8720 37120
rect 11796 37136 11848 37188
rect 16120 37179 16172 37188
rect 16120 37145 16129 37179
rect 16129 37145 16163 37179
rect 16163 37145 16172 37179
rect 16120 37136 16172 37145
rect 21824 37136 21876 37188
rect 28448 37213 28457 37247
rect 28457 37213 28491 37247
rect 28491 37213 28500 37247
rect 28448 37204 28500 37213
rect 31484 37204 31536 37256
rect 33600 37247 33652 37256
rect 33600 37213 33609 37247
rect 33609 37213 33643 37247
rect 33643 37213 33652 37247
rect 33600 37204 33652 37213
rect 35440 37204 35492 37256
rect 11060 37068 11112 37120
rect 13176 37111 13228 37120
rect 13176 37077 13185 37111
rect 13185 37077 13219 37111
rect 13219 37077 13228 37111
rect 13176 37068 13228 37077
rect 13544 37068 13596 37120
rect 15108 37111 15160 37120
rect 15108 37077 15117 37111
rect 15117 37077 15151 37111
rect 15151 37077 15160 37111
rect 15108 37068 15160 37077
rect 15200 37068 15252 37120
rect 18052 37068 18104 37120
rect 19984 37068 20036 37120
rect 21272 37068 21324 37120
rect 31852 37136 31904 37188
rect 35532 37179 35584 37188
rect 35532 37145 35541 37179
rect 35541 37145 35575 37179
rect 35575 37145 35584 37179
rect 35532 37136 35584 37145
rect 25320 37111 25372 37120
rect 25320 37077 25329 37111
rect 25329 37077 25363 37111
rect 25363 37077 25372 37111
rect 25320 37068 25372 37077
rect 26424 37068 26476 37120
rect 28356 37068 28408 37120
rect 30564 37111 30616 37120
rect 30564 37077 30573 37111
rect 30573 37077 30607 37111
rect 30607 37077 30616 37111
rect 30564 37068 30616 37077
rect 31760 37068 31812 37120
rect 33508 37068 33560 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 4620 36864 4672 36916
rect 5816 36864 5868 36916
rect 7748 36907 7800 36916
rect 7748 36873 7757 36907
rect 7757 36873 7791 36907
rect 7791 36873 7800 36907
rect 7748 36864 7800 36873
rect 11704 36907 11756 36916
rect 2964 36839 3016 36848
rect 2964 36805 2973 36839
rect 2973 36805 3007 36839
rect 3007 36805 3016 36839
rect 2964 36796 3016 36805
rect 6828 36796 6880 36848
rect 2228 36771 2280 36780
rect 2228 36737 2237 36771
rect 2237 36737 2271 36771
rect 2271 36737 2280 36771
rect 2228 36728 2280 36737
rect 2596 36728 2648 36780
rect 6552 36771 6604 36780
rect 4712 36703 4764 36712
rect 4712 36669 4721 36703
rect 4721 36669 4755 36703
rect 4755 36669 4764 36703
rect 4712 36660 4764 36669
rect 4896 36592 4948 36644
rect 6552 36737 6561 36771
rect 6561 36737 6595 36771
rect 6595 36737 6604 36771
rect 6552 36728 6604 36737
rect 10784 36796 10836 36848
rect 6460 36660 6512 36712
rect 8392 36703 8444 36712
rect 8392 36669 8401 36703
rect 8401 36669 8435 36703
rect 8435 36669 8444 36703
rect 8392 36660 8444 36669
rect 10416 36703 10468 36712
rect 10416 36669 10425 36703
rect 10425 36669 10459 36703
rect 10459 36669 10468 36703
rect 10416 36660 10468 36669
rect 10876 36660 10928 36712
rect 11704 36873 11713 36907
rect 11713 36873 11747 36907
rect 11747 36873 11756 36907
rect 11704 36864 11756 36873
rect 11796 36864 11848 36916
rect 13820 36864 13872 36916
rect 18144 36864 18196 36916
rect 35624 36864 35676 36916
rect 35808 36864 35860 36916
rect 11060 36771 11112 36780
rect 11060 36737 11069 36771
rect 11069 36737 11103 36771
rect 11103 36737 11112 36771
rect 11060 36728 11112 36737
rect 13360 36796 13412 36848
rect 15200 36796 15252 36848
rect 13084 36771 13136 36780
rect 13084 36737 13093 36771
rect 13093 36737 13127 36771
rect 13127 36737 13136 36771
rect 13084 36728 13136 36737
rect 14004 36728 14056 36780
rect 15108 36728 15160 36780
rect 35624 36771 35676 36780
rect 35624 36737 35633 36771
rect 35633 36737 35667 36771
rect 35667 36737 35676 36771
rect 35624 36728 35676 36737
rect 36176 36728 36228 36780
rect 11980 36660 12032 36712
rect 13544 36703 13596 36712
rect 13544 36669 13553 36703
rect 13553 36669 13587 36703
rect 13587 36669 13596 36703
rect 13544 36660 13596 36669
rect 16120 36660 16172 36712
rect 3148 36524 3200 36576
rect 5816 36524 5868 36576
rect 6368 36524 6420 36576
rect 7656 36524 7708 36576
rect 9036 36524 9088 36576
rect 9128 36524 9180 36576
rect 10416 36524 10468 36576
rect 14372 36592 14424 36644
rect 35532 36592 35584 36644
rect 22008 36524 22060 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 2228 36320 2280 36372
rect 4988 36252 5040 36304
rect 5172 36320 5224 36372
rect 1584 36227 1636 36236
rect 1584 36193 1593 36227
rect 1593 36193 1627 36227
rect 1627 36193 1636 36227
rect 1584 36184 1636 36193
rect 2412 36184 2464 36236
rect 5080 36184 5132 36236
rect 8300 36252 8352 36304
rect 10876 36320 10928 36372
rect 11980 36363 12032 36372
rect 11980 36329 11989 36363
rect 11989 36329 12023 36363
rect 12023 36329 12032 36363
rect 11980 36320 12032 36329
rect 13820 36320 13872 36372
rect 14832 36363 14884 36372
rect 14832 36329 14841 36363
rect 14841 36329 14875 36363
rect 14875 36329 14884 36363
rect 14832 36320 14884 36329
rect 9128 36227 9180 36236
rect 5172 36116 5224 36168
rect 5448 36159 5500 36168
rect 5448 36125 5457 36159
rect 5457 36125 5491 36159
rect 5491 36125 5500 36159
rect 5448 36116 5500 36125
rect 8300 36116 8352 36168
rect 9128 36193 9137 36227
rect 9137 36193 9171 36227
rect 9171 36193 9180 36227
rect 9128 36184 9180 36193
rect 10968 36184 11020 36236
rect 8668 36116 8720 36168
rect 12532 36252 12584 36304
rect 36728 36320 36780 36372
rect 30564 36252 30616 36304
rect 12532 36116 12584 36168
rect 15108 36116 15160 36168
rect 5908 36091 5960 36100
rect 5908 36057 5917 36091
rect 5917 36057 5951 36091
rect 5951 36057 5960 36091
rect 5908 36048 5960 36057
rect 6276 36048 6328 36100
rect 7656 36091 7708 36100
rect 7656 36057 7665 36091
rect 7665 36057 7699 36091
rect 7699 36057 7708 36091
rect 7656 36048 7708 36057
rect 4068 35980 4120 36032
rect 9680 35980 9732 36032
rect 9864 36048 9916 36100
rect 11060 36048 11112 36100
rect 14372 36048 14424 36100
rect 10416 35980 10468 36032
rect 10876 36023 10928 36032
rect 10876 35989 10885 36023
rect 10885 35989 10919 36023
rect 10919 35989 10928 36023
rect 10876 35980 10928 35989
rect 12440 35980 12492 36032
rect 13544 35980 13596 36032
rect 15936 36023 15988 36032
rect 15936 35989 15945 36023
rect 15945 35989 15979 36023
rect 15979 35989 15988 36023
rect 15936 35980 15988 35989
rect 35348 35980 35400 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 3332 35776 3384 35828
rect 3792 35776 3844 35828
rect 6736 35776 6788 35828
rect 6184 35708 6236 35760
rect 1584 35683 1636 35692
rect 1584 35649 1593 35683
rect 1593 35649 1627 35683
rect 1627 35649 1636 35683
rect 1584 35640 1636 35649
rect 5724 35640 5776 35692
rect 7104 35708 7156 35760
rect 9036 35708 9088 35760
rect 2596 35572 2648 35624
rect 4712 35572 4764 35624
rect 6368 35572 6420 35624
rect 6552 35572 6604 35624
rect 8668 35572 8720 35624
rect 9772 35683 9824 35692
rect 9772 35649 9781 35683
rect 9781 35649 9815 35683
rect 9815 35649 9824 35683
rect 9772 35640 9824 35649
rect 10416 35640 10468 35692
rect 9220 35572 9272 35624
rect 2964 35436 3016 35488
rect 5724 35436 5776 35488
rect 6552 35479 6604 35488
rect 6552 35445 6561 35479
rect 6561 35445 6595 35479
rect 6595 35445 6604 35479
rect 6552 35436 6604 35445
rect 10508 35504 10560 35556
rect 9956 35479 10008 35488
rect 9956 35445 9965 35479
rect 9965 35445 9999 35479
rect 9999 35445 10008 35479
rect 9956 35436 10008 35445
rect 10416 35479 10468 35488
rect 10416 35445 10425 35479
rect 10425 35445 10459 35479
rect 10459 35445 10468 35479
rect 10416 35436 10468 35445
rect 12992 35776 13044 35828
rect 13544 35819 13596 35828
rect 13544 35785 13553 35819
rect 13553 35785 13587 35819
rect 13587 35785 13596 35819
rect 13544 35776 13596 35785
rect 15108 35776 15160 35828
rect 15936 35776 15988 35828
rect 12440 35751 12492 35760
rect 12440 35717 12449 35751
rect 12449 35717 12483 35751
rect 12483 35717 12492 35751
rect 12440 35708 12492 35717
rect 12624 35640 12676 35692
rect 15476 35640 15528 35692
rect 11980 35615 12032 35624
rect 11980 35581 11989 35615
rect 11989 35581 12023 35615
rect 12023 35581 12032 35615
rect 11980 35572 12032 35581
rect 15568 35572 15620 35624
rect 35440 35436 35492 35488
rect 36268 35479 36320 35488
rect 36268 35445 36277 35479
rect 36277 35445 36311 35479
rect 36311 35445 36320 35479
rect 36268 35436 36320 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 1768 35232 1820 35284
rect 2596 35096 2648 35148
rect 3884 35096 3936 35148
rect 4988 35028 5040 35080
rect 5448 35028 5500 35080
rect 1584 34935 1636 34944
rect 1584 34901 1593 34935
rect 1593 34901 1627 34935
rect 1627 34901 1636 34935
rect 1584 34892 1636 34901
rect 4068 34960 4120 35012
rect 4712 34960 4764 35012
rect 7288 35232 7340 35284
rect 7380 35232 7432 35284
rect 9772 35232 9824 35284
rect 9956 35232 10008 35284
rect 13544 35232 13596 35284
rect 14832 35275 14884 35284
rect 14832 35241 14841 35275
rect 14841 35241 14875 35275
rect 14875 35241 14884 35275
rect 14832 35232 14884 35241
rect 28448 35232 28500 35284
rect 6552 35096 6604 35148
rect 8300 35096 8352 35148
rect 8760 35096 8812 35148
rect 9128 35139 9180 35148
rect 9128 35105 9137 35139
rect 9137 35105 9171 35139
rect 9171 35105 9180 35139
rect 9128 35096 9180 35105
rect 14004 35164 14056 35216
rect 10692 35096 10744 35148
rect 11704 35096 11756 35148
rect 11796 35139 11848 35148
rect 11796 35105 11805 35139
rect 11805 35105 11839 35139
rect 11839 35105 11848 35139
rect 11796 35096 11848 35105
rect 12900 35096 12952 35148
rect 13176 35096 13228 35148
rect 15568 35071 15620 35080
rect 15568 35037 15577 35071
rect 15577 35037 15611 35071
rect 15611 35037 15620 35071
rect 15568 35028 15620 35037
rect 27896 35071 27948 35080
rect 27896 35037 27905 35071
rect 27905 35037 27939 35071
rect 27939 35037 27948 35071
rect 27896 35028 27948 35037
rect 35900 35028 35952 35080
rect 5632 34960 5684 35012
rect 7472 34960 7524 35012
rect 6184 34892 6236 34944
rect 7012 34892 7064 34944
rect 8484 34960 8536 35012
rect 9036 34960 9088 35012
rect 9680 34960 9732 35012
rect 8392 34892 8444 34944
rect 10784 34892 10836 34944
rect 11612 35003 11664 35012
rect 11612 34969 11621 35003
rect 11621 34969 11655 35003
rect 11655 34969 11664 35003
rect 11612 34960 11664 34969
rect 12532 34892 12584 34944
rect 15660 34935 15712 34944
rect 15660 34901 15669 34935
rect 15669 34901 15703 34935
rect 15703 34901 15712 34935
rect 15660 34892 15712 34901
rect 16948 34892 17000 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 2412 34688 2464 34740
rect 2688 34688 2740 34740
rect 3240 34620 3292 34672
rect 3700 34663 3752 34672
rect 3700 34629 3709 34663
rect 3709 34629 3743 34663
rect 3743 34629 3752 34663
rect 3700 34620 3752 34629
rect 5724 34688 5776 34740
rect 6828 34688 6880 34740
rect 1768 34595 1820 34604
rect 1768 34561 1777 34595
rect 1777 34561 1811 34595
rect 1811 34561 1820 34595
rect 1768 34552 1820 34561
rect 3976 34595 4028 34604
rect 3976 34561 3985 34595
rect 3985 34561 4019 34595
rect 4019 34561 4028 34595
rect 5172 34620 5224 34672
rect 5356 34620 5408 34672
rect 9864 34688 9916 34740
rect 9956 34688 10008 34740
rect 14832 34688 14884 34740
rect 15108 34731 15160 34740
rect 15108 34697 15117 34731
rect 15117 34697 15151 34731
rect 15151 34697 15160 34731
rect 15108 34688 15160 34697
rect 8484 34620 8536 34672
rect 9496 34620 9548 34672
rect 10140 34620 10192 34672
rect 10600 34620 10652 34672
rect 11796 34663 11848 34672
rect 11796 34629 11805 34663
rect 11805 34629 11839 34663
rect 11839 34629 11848 34663
rect 11796 34620 11848 34629
rect 15660 34620 15712 34672
rect 3976 34552 4028 34561
rect 4988 34552 5040 34604
rect 5540 34595 5592 34604
rect 5540 34561 5549 34595
rect 5549 34561 5583 34595
rect 5583 34561 5592 34595
rect 5540 34552 5592 34561
rect 6828 34552 6880 34604
rect 10968 34595 11020 34604
rect 10968 34561 10977 34595
rect 10977 34561 11011 34595
rect 11011 34561 11020 34595
rect 10968 34552 11020 34561
rect 13268 34552 13320 34604
rect 5356 34527 5408 34536
rect 5356 34493 5365 34527
rect 5365 34493 5399 34527
rect 5399 34493 5408 34527
rect 5356 34484 5408 34493
rect 9404 34484 9456 34536
rect 9772 34527 9824 34536
rect 9772 34493 9781 34527
rect 9781 34493 9815 34527
rect 9815 34493 9824 34527
rect 9772 34484 9824 34493
rect 5540 34416 5592 34468
rect 5908 34416 5960 34468
rect 6644 34416 6696 34468
rect 9588 34348 9640 34400
rect 11980 34484 12032 34536
rect 13176 34484 13228 34536
rect 16948 34527 17000 34536
rect 11796 34416 11848 34468
rect 12348 34416 12400 34468
rect 16948 34493 16957 34527
rect 16957 34493 16991 34527
rect 16991 34493 17000 34527
rect 16948 34484 17000 34493
rect 11520 34348 11572 34400
rect 34796 34348 34848 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 3976 34187 4028 34196
rect 3976 34153 3985 34187
rect 3985 34153 4019 34187
rect 4019 34153 4028 34187
rect 3976 34144 4028 34153
rect 5816 34144 5868 34196
rect 7840 34144 7892 34196
rect 12992 34187 13044 34196
rect 6644 34076 6696 34128
rect 8760 34076 8812 34128
rect 9588 34076 9640 34128
rect 12992 34153 13001 34187
rect 13001 34153 13035 34187
rect 13035 34153 13044 34187
rect 12992 34144 13044 34153
rect 14372 34187 14424 34196
rect 14372 34153 14381 34187
rect 14381 34153 14415 34187
rect 14415 34153 14424 34187
rect 14372 34144 14424 34153
rect 15108 34144 15160 34196
rect 5908 34008 5960 34060
rect 6184 34008 6236 34060
rect 6552 34051 6604 34060
rect 6552 34017 6561 34051
rect 6561 34017 6595 34051
rect 6595 34017 6604 34051
rect 6552 34008 6604 34017
rect 6736 34008 6788 34060
rect 7196 33983 7248 33992
rect 2228 33804 2280 33856
rect 7196 33949 7205 33983
rect 7205 33949 7239 33983
rect 7239 33949 7248 33983
rect 7196 33940 7248 33949
rect 7380 33940 7432 33992
rect 14464 34076 14516 34128
rect 9772 34008 9824 34060
rect 4804 33872 4856 33924
rect 5908 33804 5960 33856
rect 6368 33872 6420 33924
rect 7932 33872 7984 33924
rect 7196 33804 7248 33856
rect 10784 33940 10836 33992
rect 14372 33940 14424 33992
rect 34796 33940 34848 33992
rect 8208 33872 8260 33924
rect 11428 33915 11480 33924
rect 11428 33881 11437 33915
rect 11437 33881 11471 33915
rect 11471 33881 11480 33915
rect 11428 33872 11480 33881
rect 11520 33915 11572 33924
rect 11520 33881 11529 33915
rect 11529 33881 11563 33915
rect 11563 33881 11572 33915
rect 11520 33872 11572 33881
rect 12348 33872 12400 33924
rect 8668 33804 8720 33856
rect 10968 33804 11020 33856
rect 13268 33804 13320 33856
rect 13636 33847 13688 33856
rect 13636 33813 13645 33847
rect 13645 33813 13679 33847
rect 13679 33813 13688 33847
rect 13636 33804 13688 33813
rect 34980 33847 35032 33856
rect 34980 33813 34989 33847
rect 34989 33813 35023 33847
rect 35023 33813 35032 33847
rect 34980 33804 35032 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 2228 33600 2280 33652
rect 4988 33600 5040 33652
rect 7104 33600 7156 33652
rect 7288 33643 7340 33652
rect 7288 33609 7297 33643
rect 7297 33609 7331 33643
rect 7331 33609 7340 33643
rect 7288 33600 7340 33609
rect 9312 33600 9364 33652
rect 1676 33464 1728 33516
rect 2504 33532 2556 33584
rect 3608 33532 3660 33584
rect 5448 33532 5500 33584
rect 8208 33532 8260 33584
rect 8392 33532 8444 33584
rect 10416 33532 10468 33584
rect 6552 33507 6604 33516
rect 6552 33473 6561 33507
rect 6561 33473 6595 33507
rect 6595 33473 6604 33507
rect 6552 33464 6604 33473
rect 6828 33464 6880 33516
rect 7196 33464 7248 33516
rect 11612 33600 11664 33652
rect 15108 33600 15160 33652
rect 31484 33643 31536 33652
rect 31484 33609 31493 33643
rect 31493 33609 31527 33643
rect 31527 33609 31536 33643
rect 31484 33600 31536 33609
rect 10784 33532 10836 33584
rect 12256 33532 12308 33584
rect 13268 33507 13320 33516
rect 13268 33473 13277 33507
rect 13277 33473 13311 33507
rect 13311 33473 13320 33507
rect 13268 33464 13320 33473
rect 14004 33464 14056 33516
rect 2228 33439 2280 33448
rect 2228 33405 2237 33439
rect 2237 33405 2271 33439
rect 2271 33405 2280 33439
rect 2228 33396 2280 33405
rect 3700 33439 3752 33448
rect 3700 33405 3709 33439
rect 3709 33405 3743 33439
rect 3743 33405 3752 33439
rect 3700 33396 3752 33405
rect 6092 33396 6144 33448
rect 7288 33396 7340 33448
rect 8852 33396 8904 33448
rect 9588 33396 9640 33448
rect 34980 33464 35032 33516
rect 36452 33396 36504 33448
rect 7840 33328 7892 33380
rect 36268 33371 36320 33380
rect 36268 33337 36277 33371
rect 36277 33337 36311 33371
rect 36311 33337 36320 33371
rect 36268 33328 36320 33337
rect 4160 33260 4212 33312
rect 10968 33260 11020 33312
rect 13544 33260 13596 33312
rect 14372 33260 14424 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 1584 33056 1636 33108
rect 5448 33099 5500 33108
rect 1676 32963 1728 32972
rect 1676 32929 1685 32963
rect 1685 32929 1719 32963
rect 1719 32929 1728 32963
rect 1676 32920 1728 32929
rect 4804 32988 4856 33040
rect 5448 33065 5457 33099
rect 5457 33065 5491 33099
rect 5491 33065 5500 33099
rect 5448 33056 5500 33065
rect 6276 33056 6328 33108
rect 3332 32852 3384 32904
rect 4896 32920 4948 32972
rect 5264 32920 5316 32972
rect 5448 32852 5500 32904
rect 5540 32895 5592 32904
rect 5540 32861 5549 32895
rect 5549 32861 5583 32895
rect 5583 32861 5592 32895
rect 5540 32852 5592 32861
rect 5908 32852 5960 32904
rect 4620 32784 4672 32836
rect 4896 32784 4948 32836
rect 8760 32920 8812 32972
rect 9128 32920 9180 32972
rect 10232 32920 10284 32972
rect 10968 32895 11020 32904
rect 10968 32861 10977 32895
rect 10977 32861 11011 32895
rect 11011 32861 11020 32895
rect 12716 33056 12768 33108
rect 14740 33056 14792 33108
rect 13728 32988 13780 33040
rect 10968 32852 11020 32861
rect 6644 32784 6696 32836
rect 3700 32716 3752 32768
rect 4528 32716 4580 32768
rect 5264 32716 5316 32768
rect 6552 32716 6604 32768
rect 6828 32759 6880 32768
rect 6828 32725 6837 32759
rect 6837 32725 6871 32759
rect 6871 32725 6880 32759
rect 6828 32716 6880 32725
rect 8944 32784 8996 32836
rect 10692 32827 10744 32836
rect 10692 32793 10701 32827
rect 10701 32793 10735 32827
rect 10735 32793 10744 32827
rect 13544 32827 13596 32836
rect 10692 32784 10744 32793
rect 12164 32716 12216 32768
rect 12440 32759 12492 32768
rect 12440 32725 12449 32759
rect 12449 32725 12483 32759
rect 12483 32725 12492 32759
rect 12440 32716 12492 32725
rect 13544 32793 13553 32827
rect 13553 32793 13587 32827
rect 13587 32793 13596 32827
rect 13544 32784 13596 32793
rect 13636 32827 13688 32836
rect 13636 32793 13645 32827
rect 13645 32793 13679 32827
rect 13679 32793 13688 32827
rect 13636 32784 13688 32793
rect 14832 32784 14884 32836
rect 36360 32759 36412 32768
rect 36360 32725 36369 32759
rect 36369 32725 36403 32759
rect 36403 32725 36412 32759
rect 36360 32716 36412 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 1676 32512 1728 32564
rect 1952 32512 2004 32564
rect 6644 32555 6696 32564
rect 1676 32376 1728 32428
rect 2412 32376 2464 32428
rect 3700 32351 3752 32360
rect 3700 32317 3709 32351
rect 3709 32317 3743 32351
rect 3743 32317 3752 32351
rect 3700 32308 3752 32317
rect 4160 32376 4212 32428
rect 4896 32376 4948 32428
rect 4068 32308 4120 32360
rect 2596 32240 2648 32292
rect 6644 32521 6653 32555
rect 6653 32521 6687 32555
rect 6687 32521 6696 32555
rect 6644 32512 6696 32521
rect 7012 32512 7064 32564
rect 7472 32444 7524 32496
rect 5540 32376 5592 32428
rect 7196 32376 7248 32428
rect 7288 32376 7340 32428
rect 8944 32512 8996 32564
rect 9128 32512 9180 32564
rect 7748 32444 7800 32496
rect 10232 32444 10284 32496
rect 12716 32512 12768 32564
rect 12808 32512 12860 32564
rect 13176 32512 13228 32564
rect 12440 32444 12492 32496
rect 10324 32376 10376 32428
rect 10784 32376 10836 32428
rect 8668 32308 8720 32360
rect 9496 32308 9548 32360
rect 13728 32308 13780 32360
rect 36084 32351 36136 32360
rect 36084 32317 36093 32351
rect 36093 32317 36127 32351
rect 36127 32317 36136 32351
rect 36084 32308 36136 32317
rect 36360 32351 36412 32360
rect 36360 32317 36369 32351
rect 36369 32317 36403 32351
rect 36403 32317 36412 32351
rect 36360 32308 36412 32317
rect 10324 32240 10376 32292
rect 10968 32240 11020 32292
rect 14004 32240 14056 32292
rect 3976 32172 4028 32224
rect 8484 32172 8536 32224
rect 14188 32172 14240 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 3240 31968 3292 32020
rect 4620 31968 4672 32020
rect 8392 31968 8444 32020
rect 9128 32011 9180 32020
rect 9128 31977 9137 32011
rect 9137 31977 9171 32011
rect 9171 31977 9180 32011
rect 9128 31968 9180 31977
rect 10416 31968 10468 32020
rect 4804 31900 4856 31952
rect 2228 31832 2280 31884
rect 3700 31832 3752 31884
rect 4896 31832 4948 31884
rect 2136 31807 2188 31816
rect 2136 31773 2145 31807
rect 2145 31773 2179 31807
rect 2179 31773 2188 31807
rect 2136 31764 2188 31773
rect 2964 31764 3016 31816
rect 3884 31764 3936 31816
rect 4620 31764 4672 31816
rect 5080 31764 5132 31816
rect 5264 31900 5316 31952
rect 6460 31900 6512 31952
rect 6552 31900 6604 31952
rect 5816 31832 5868 31884
rect 6092 31832 6144 31884
rect 10692 31900 10744 31952
rect 35624 31968 35676 32020
rect 5448 31764 5500 31816
rect 6552 31764 6604 31816
rect 9772 31764 9824 31816
rect 9956 31807 10008 31816
rect 9956 31773 9965 31807
rect 9965 31773 9999 31807
rect 9999 31773 10008 31807
rect 10600 31832 10652 31884
rect 9956 31764 10008 31773
rect 11336 31764 11388 31816
rect 12716 31832 12768 31884
rect 13544 31875 13596 31884
rect 13544 31841 13553 31875
rect 13553 31841 13587 31875
rect 13587 31841 13596 31875
rect 13544 31832 13596 31841
rect 6000 31696 6052 31748
rect 7012 31739 7064 31748
rect 7012 31705 7021 31739
rect 7021 31705 7055 31739
rect 7055 31705 7064 31739
rect 7012 31696 7064 31705
rect 7288 31696 7340 31748
rect 11060 31696 11112 31748
rect 13360 31764 13412 31816
rect 14096 31764 14148 31816
rect 15384 31764 15436 31816
rect 19432 31764 19484 31816
rect 27896 31764 27948 31816
rect 35992 31764 36044 31816
rect 13452 31696 13504 31748
rect 13820 31696 13872 31748
rect 4436 31628 4488 31680
rect 9588 31628 9640 31680
rect 11888 31628 11940 31680
rect 13728 31628 13780 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 4712 31424 4764 31476
rect 5080 31424 5132 31476
rect 5172 31424 5224 31476
rect 5356 31424 5408 31476
rect 5724 31424 5776 31476
rect 7288 31467 7340 31476
rect 7288 31433 7297 31467
rect 7297 31433 7331 31467
rect 7331 31433 7340 31467
rect 7288 31424 7340 31433
rect 7932 31467 7984 31476
rect 7932 31433 7941 31467
rect 7941 31433 7975 31467
rect 7975 31433 7984 31467
rect 7932 31424 7984 31433
rect 9128 31424 9180 31476
rect 9588 31424 9640 31476
rect 36084 31424 36136 31476
rect 3976 31356 4028 31408
rect 4436 31399 4488 31408
rect 4436 31365 4445 31399
rect 4445 31365 4479 31399
rect 4479 31365 4488 31399
rect 4436 31356 4488 31365
rect 1952 31331 2004 31340
rect 1952 31297 1961 31331
rect 1961 31297 1995 31331
rect 1995 31297 2004 31331
rect 1952 31288 2004 31297
rect 5724 31288 5776 31340
rect 6000 31288 6052 31340
rect 2596 31220 2648 31272
rect 4160 31263 4212 31272
rect 4160 31229 4169 31263
rect 4169 31229 4203 31263
rect 4203 31229 4212 31263
rect 4160 31220 4212 31229
rect 3884 31152 3936 31204
rect 5448 31220 5500 31272
rect 7380 31288 7432 31340
rect 8852 31356 8904 31408
rect 9220 31356 9272 31408
rect 11336 31356 11388 31408
rect 12808 31399 12860 31408
rect 12808 31365 12817 31399
rect 12817 31365 12851 31399
rect 12851 31365 12860 31399
rect 12808 31356 12860 31365
rect 14188 31399 14240 31408
rect 14188 31365 14197 31399
rect 14197 31365 14231 31399
rect 14231 31365 14240 31399
rect 14188 31356 14240 31365
rect 15384 31399 15436 31408
rect 15384 31365 15393 31399
rect 15393 31365 15427 31399
rect 15427 31365 15436 31399
rect 15384 31356 15436 31365
rect 19432 31356 19484 31408
rect 9128 31220 9180 31272
rect 12624 31220 12676 31272
rect 12808 31220 12860 31272
rect 15200 31220 15252 31272
rect 3700 31127 3752 31136
rect 3700 31093 3709 31127
rect 3709 31093 3743 31127
rect 3743 31093 3752 31127
rect 3700 31084 3752 31093
rect 4436 31084 4488 31136
rect 5448 31084 5500 31136
rect 10048 31084 10100 31136
rect 10416 31084 10468 31136
rect 10968 31084 11020 31136
rect 11428 31084 11480 31136
rect 12348 31084 12400 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 6460 30880 6512 30932
rect 10784 30880 10836 30932
rect 2412 30676 2464 30728
rect 1492 30608 1544 30660
rect 8300 30744 8352 30796
rect 8852 30744 8904 30796
rect 11152 30744 11204 30796
rect 14372 30787 14424 30796
rect 14372 30753 14381 30787
rect 14381 30753 14415 30787
rect 14415 30753 14424 30787
rect 14372 30744 14424 30753
rect 2964 30719 3016 30728
rect 2964 30685 2973 30719
rect 2973 30685 3007 30719
rect 3007 30685 3016 30719
rect 2964 30676 3016 30685
rect 5816 30719 5868 30728
rect 5816 30685 5825 30719
rect 5825 30685 5859 30719
rect 5859 30685 5868 30719
rect 5816 30676 5868 30685
rect 7196 30676 7248 30728
rect 13084 30676 13136 30728
rect 15476 30676 15528 30728
rect 15844 30676 15896 30728
rect 3056 30540 3108 30592
rect 4804 30608 4856 30660
rect 5540 30651 5592 30660
rect 5540 30617 5549 30651
rect 5549 30617 5583 30651
rect 5583 30617 5592 30651
rect 5540 30608 5592 30617
rect 6644 30540 6696 30592
rect 9312 30608 9364 30660
rect 10600 30651 10652 30660
rect 10600 30617 10609 30651
rect 10609 30617 10643 30651
rect 10643 30617 10652 30651
rect 10600 30608 10652 30617
rect 11336 30608 11388 30660
rect 11888 30651 11940 30660
rect 11888 30617 11897 30651
rect 11897 30617 11931 30651
rect 11931 30617 11940 30651
rect 12808 30651 12860 30660
rect 11888 30608 11940 30617
rect 12808 30617 12817 30651
rect 12817 30617 12851 30651
rect 12851 30617 12860 30651
rect 12808 30608 12860 30617
rect 14188 30608 14240 30660
rect 13084 30540 13136 30592
rect 13728 30540 13780 30592
rect 15200 30608 15252 30660
rect 16212 30608 16264 30660
rect 15568 30583 15620 30592
rect 15568 30549 15577 30583
rect 15577 30549 15611 30583
rect 15611 30549 15620 30583
rect 15568 30540 15620 30549
rect 15844 30540 15896 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 7932 30336 7984 30388
rect 8300 30336 8352 30388
rect 12808 30336 12860 30388
rect 19340 30336 19392 30388
rect 1952 30268 2004 30320
rect 2320 30268 2372 30320
rect 5540 30268 5592 30320
rect 4160 30200 4212 30252
rect 6552 30243 6604 30252
rect 6552 30209 6561 30243
rect 6561 30209 6595 30243
rect 6595 30209 6604 30243
rect 6552 30200 6604 30209
rect 3148 30132 3200 30184
rect 5908 30132 5960 30184
rect 8024 30268 8076 30320
rect 10140 30200 10192 30252
rect 12164 30243 12216 30252
rect 12164 30209 12173 30243
rect 12173 30209 12207 30243
rect 12207 30209 12216 30243
rect 12164 30200 12216 30209
rect 13912 30200 13964 30252
rect 14096 30200 14148 30252
rect 14280 30200 14332 30252
rect 15108 30200 15160 30252
rect 35900 30200 35952 30252
rect 6828 30132 6880 30184
rect 3700 30064 3752 30116
rect 3240 29996 3292 30048
rect 7380 30064 7432 30116
rect 7932 30175 7984 30184
rect 7932 30141 7941 30175
rect 7941 30141 7975 30175
rect 7975 30141 7984 30175
rect 7932 30132 7984 30141
rect 8024 30132 8076 30184
rect 11060 30132 11112 30184
rect 12992 30132 13044 30184
rect 14372 30132 14424 30184
rect 16028 30175 16080 30184
rect 16028 30141 16037 30175
rect 16037 30141 16071 30175
rect 16071 30141 16080 30175
rect 16028 30132 16080 30141
rect 36360 30175 36412 30184
rect 36360 30141 36369 30175
rect 36369 30141 36403 30175
rect 36403 30141 36412 30175
rect 36360 30132 36412 30141
rect 13176 30064 13228 30116
rect 8576 29996 8628 30048
rect 9772 29996 9824 30048
rect 10508 29996 10560 30048
rect 11980 29996 12032 30048
rect 12440 29996 12492 30048
rect 12900 29996 12952 30048
rect 13728 29996 13780 30048
rect 14096 30039 14148 30048
rect 14096 30005 14105 30039
rect 14105 30005 14139 30039
rect 14139 30005 14148 30039
rect 14096 29996 14148 30005
rect 15016 29996 15068 30048
rect 15108 29996 15160 30048
rect 25872 29996 25924 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 1676 29835 1728 29844
rect 1676 29801 1685 29835
rect 1685 29801 1719 29835
rect 1719 29801 1728 29835
rect 1676 29792 1728 29801
rect 2320 29835 2372 29844
rect 2320 29801 2329 29835
rect 2329 29801 2363 29835
rect 2363 29801 2372 29835
rect 2320 29792 2372 29801
rect 3976 29792 4028 29844
rect 4160 29792 4212 29844
rect 5816 29792 5868 29844
rect 5908 29792 5960 29844
rect 8852 29792 8904 29844
rect 9496 29792 9548 29844
rect 3608 29724 3660 29776
rect 2964 29656 3016 29708
rect 2412 29588 2464 29640
rect 4620 29656 4672 29708
rect 4160 29631 4212 29640
rect 4160 29597 4169 29631
rect 4169 29597 4203 29631
rect 4203 29597 4212 29631
rect 4160 29588 4212 29597
rect 4712 29588 4764 29640
rect 5264 29588 5316 29640
rect 6552 29656 6604 29708
rect 6828 29699 6880 29708
rect 6828 29665 6837 29699
rect 6837 29665 6871 29699
rect 6871 29665 6880 29699
rect 6828 29656 6880 29665
rect 8116 29724 8168 29776
rect 10600 29792 10652 29844
rect 11704 29792 11756 29844
rect 12348 29792 12400 29844
rect 36360 29835 36412 29844
rect 12164 29724 12216 29776
rect 12808 29724 12860 29776
rect 36360 29801 36369 29835
rect 36369 29801 36403 29835
rect 36403 29801 36412 29835
rect 36360 29792 36412 29801
rect 14280 29724 14332 29776
rect 13636 29656 13688 29708
rect 16212 29699 16264 29708
rect 16212 29665 16221 29699
rect 16221 29665 16255 29699
rect 16255 29665 16264 29699
rect 16212 29656 16264 29665
rect 6276 29520 6328 29572
rect 6736 29520 6788 29572
rect 7380 29520 7432 29572
rect 7564 29520 7616 29572
rect 11152 29588 11204 29640
rect 12532 29588 12584 29640
rect 12808 29588 12860 29640
rect 11060 29520 11112 29572
rect 4160 29452 4212 29504
rect 8484 29452 8536 29504
rect 11520 29563 11572 29572
rect 11520 29529 11529 29563
rect 11529 29529 11563 29563
rect 11563 29529 11572 29563
rect 12992 29563 13044 29572
rect 11520 29520 11572 29529
rect 12992 29529 13001 29563
rect 13001 29529 13035 29563
rect 13035 29529 13044 29563
rect 12992 29520 13044 29529
rect 13176 29520 13228 29572
rect 16396 29563 16448 29572
rect 12900 29452 12952 29504
rect 16396 29529 16405 29563
rect 16405 29529 16439 29563
rect 16439 29529 16448 29563
rect 16396 29520 16448 29529
rect 16856 29520 16908 29572
rect 15568 29452 15620 29504
rect 17500 29452 17552 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 1584 29087 1636 29096
rect 1584 29053 1593 29087
rect 1593 29053 1627 29087
rect 1627 29053 1636 29087
rect 1584 29044 1636 29053
rect 3148 29248 3200 29300
rect 3056 29180 3108 29232
rect 5816 29248 5868 29300
rect 6276 29248 6328 29300
rect 6460 29180 6512 29232
rect 7288 29180 7340 29232
rect 6552 29155 6604 29164
rect 6552 29121 6561 29155
rect 6561 29121 6595 29155
rect 6595 29121 6604 29155
rect 6552 29112 6604 29121
rect 11520 29248 11572 29300
rect 12164 29248 12216 29300
rect 13912 29248 13964 29300
rect 14556 29248 14608 29300
rect 9680 29180 9732 29232
rect 9956 29180 10008 29232
rect 11704 29180 11756 29232
rect 12440 29223 12492 29232
rect 12440 29189 12449 29223
rect 12449 29189 12483 29223
rect 12483 29189 12492 29223
rect 12440 29180 12492 29189
rect 12716 29180 12768 29232
rect 14004 29180 14056 29232
rect 17132 29248 17184 29300
rect 16212 29180 16264 29232
rect 18144 29248 18196 29300
rect 17500 29223 17552 29232
rect 17500 29189 17509 29223
rect 17509 29189 17543 29223
rect 17543 29189 17552 29223
rect 17500 29180 17552 29189
rect 8852 29112 8904 29164
rect 18052 29155 18104 29164
rect 18052 29121 18061 29155
rect 18061 29121 18095 29155
rect 18095 29121 18104 29155
rect 18052 29112 18104 29121
rect 5172 28976 5224 29028
rect 4804 28908 4856 28960
rect 5356 28908 5408 28960
rect 7380 28908 7432 28960
rect 8484 29044 8536 29096
rect 10784 29044 10836 29096
rect 8300 29019 8352 29028
rect 8300 28985 8309 29019
rect 8309 28985 8343 29019
rect 8343 28985 8352 29019
rect 8300 28976 8352 28985
rect 9128 28976 9180 29028
rect 10232 28976 10284 29028
rect 10324 28976 10376 29028
rect 13360 28976 13412 29028
rect 13636 29044 13688 29096
rect 14556 29087 14608 29096
rect 14556 29053 14565 29087
rect 14565 29053 14599 29087
rect 14599 29053 14608 29087
rect 14556 29044 14608 29053
rect 16396 29044 16448 29096
rect 16304 28976 16356 29028
rect 12532 28908 12584 28960
rect 13636 28908 13688 28960
rect 18052 28908 18104 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 4068 28747 4120 28756
rect 4068 28713 4077 28747
rect 4077 28713 4111 28747
rect 4111 28713 4120 28747
rect 4068 28704 4120 28713
rect 5816 28747 5868 28756
rect 5816 28713 5825 28747
rect 5825 28713 5859 28747
rect 5859 28713 5868 28747
rect 5816 28704 5868 28713
rect 7288 28704 7340 28756
rect 7380 28704 7432 28756
rect 2504 28568 2556 28620
rect 4988 28568 5040 28620
rect 6552 28568 6604 28620
rect 2872 28543 2924 28552
rect 2872 28509 2881 28543
rect 2881 28509 2915 28543
rect 2915 28509 2924 28543
rect 2872 28500 2924 28509
rect 13360 28704 13412 28756
rect 13820 28704 13872 28756
rect 14832 28704 14884 28756
rect 18144 28747 18196 28756
rect 10784 28568 10836 28620
rect 11612 28568 11664 28620
rect 12348 28568 12400 28620
rect 15016 28636 15068 28688
rect 15292 28611 15344 28620
rect 15292 28577 15301 28611
rect 15301 28577 15335 28611
rect 15335 28577 15344 28611
rect 15292 28568 15344 28577
rect 16028 28568 16080 28620
rect 16488 28568 16540 28620
rect 1676 28407 1728 28416
rect 1676 28373 1685 28407
rect 1685 28373 1719 28407
rect 1719 28373 1728 28407
rect 1676 28364 1728 28373
rect 8300 28432 8352 28484
rect 8392 28432 8444 28484
rect 14648 28500 14700 28552
rect 18144 28713 18153 28747
rect 18153 28713 18187 28747
rect 18187 28713 18196 28747
rect 18144 28704 18196 28713
rect 18052 28500 18104 28552
rect 35992 28500 36044 28552
rect 11060 28432 11112 28484
rect 11336 28475 11388 28484
rect 11336 28441 11345 28475
rect 11345 28441 11379 28475
rect 11379 28441 11388 28475
rect 11336 28432 11388 28441
rect 2872 28364 2924 28416
rect 3884 28364 3936 28416
rect 5264 28407 5316 28416
rect 5264 28373 5273 28407
rect 5273 28373 5307 28407
rect 5307 28373 5316 28407
rect 5264 28364 5316 28373
rect 7012 28364 7064 28416
rect 7932 28364 7984 28416
rect 11428 28364 11480 28416
rect 11980 28475 12032 28484
rect 11980 28441 11989 28475
rect 11989 28441 12023 28475
rect 12023 28441 12032 28475
rect 12532 28475 12584 28484
rect 11980 28432 12032 28441
rect 12532 28441 12541 28475
rect 12541 28441 12575 28475
rect 12575 28441 12584 28475
rect 12532 28432 12584 28441
rect 15476 28475 15528 28484
rect 15476 28441 15485 28475
rect 15485 28441 15519 28475
rect 15519 28441 15528 28475
rect 15476 28432 15528 28441
rect 15568 28475 15620 28484
rect 15568 28441 15577 28475
rect 15577 28441 15611 28475
rect 15611 28441 15620 28475
rect 15568 28432 15620 28441
rect 14096 28364 14148 28416
rect 14372 28407 14424 28416
rect 14372 28373 14381 28407
rect 14381 28373 14415 28407
rect 14415 28373 14424 28407
rect 14372 28364 14424 28373
rect 16856 28475 16908 28484
rect 16856 28441 16865 28475
rect 16865 28441 16899 28475
rect 16899 28441 16908 28475
rect 16856 28432 16908 28441
rect 18696 28407 18748 28416
rect 18696 28373 18705 28407
rect 18705 28373 18739 28407
rect 18739 28373 18748 28407
rect 18696 28364 18748 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 3240 28160 3292 28212
rect 4068 28203 4120 28212
rect 4068 28169 4077 28203
rect 4077 28169 4111 28203
rect 4111 28169 4120 28203
rect 4068 28160 4120 28169
rect 1676 28092 1728 28144
rect 9312 28160 9364 28212
rect 11060 28203 11112 28212
rect 11060 28169 11069 28203
rect 11069 28169 11103 28203
rect 11103 28169 11112 28203
rect 11060 28160 11112 28169
rect 12256 28160 12308 28212
rect 15476 28160 15528 28212
rect 4988 28092 5040 28144
rect 9496 28135 9548 28144
rect 2412 28024 2464 28076
rect 2872 28067 2924 28076
rect 2872 28033 2881 28067
rect 2881 28033 2915 28067
rect 2915 28033 2924 28067
rect 2872 28024 2924 28033
rect 5080 28024 5132 28076
rect 9496 28101 9505 28135
rect 9505 28101 9539 28135
rect 9539 28101 9548 28135
rect 9496 28092 9548 28101
rect 12440 28092 12492 28144
rect 13544 28135 13596 28144
rect 13544 28101 13553 28135
rect 13553 28101 13587 28135
rect 13587 28101 13596 28135
rect 13544 28092 13596 28101
rect 15752 28135 15804 28144
rect 15752 28101 15761 28135
rect 15761 28101 15795 28135
rect 15795 28101 15804 28135
rect 15752 28092 15804 28101
rect 16304 28135 16356 28144
rect 16304 28101 16313 28135
rect 16313 28101 16347 28135
rect 16347 28101 16356 28135
rect 16304 28092 16356 28101
rect 7840 28067 7892 28076
rect 7840 28033 7849 28067
rect 7849 28033 7883 28067
rect 7883 28033 7892 28067
rect 7840 28024 7892 28033
rect 7932 28024 7984 28076
rect 10416 28024 10468 28076
rect 11244 28024 11296 28076
rect 11888 28024 11940 28076
rect 18052 28067 18104 28076
rect 18052 28033 18061 28067
rect 18061 28033 18095 28067
rect 18095 28033 18104 28067
rect 18052 28024 18104 28033
rect 18696 28067 18748 28076
rect 18696 28033 18705 28067
rect 18705 28033 18739 28067
rect 18739 28033 18748 28067
rect 18696 28024 18748 28033
rect 36452 28024 36504 28076
rect 5540 27956 5592 28008
rect 5816 27956 5868 28008
rect 12624 27956 12676 28008
rect 14280 27956 14332 28008
rect 15016 27999 15068 28008
rect 15016 27965 15025 27999
rect 15025 27965 15059 27999
rect 15059 27965 15068 27999
rect 15016 27956 15068 27965
rect 4620 27888 4672 27940
rect 1584 27863 1636 27872
rect 1584 27829 1593 27863
rect 1593 27829 1627 27863
rect 1627 27829 1636 27863
rect 1584 27820 1636 27829
rect 2136 27820 2188 27872
rect 8392 27888 8444 27940
rect 9312 27888 9364 27940
rect 12992 27931 13044 27940
rect 12992 27897 13001 27931
rect 13001 27897 13035 27931
rect 13035 27897 13044 27931
rect 12992 27888 13044 27897
rect 15568 27888 15620 27940
rect 17316 27956 17368 28008
rect 36360 27999 36412 28008
rect 36360 27965 36369 27999
rect 36369 27965 36403 27999
rect 36403 27965 36412 27999
rect 36360 27956 36412 27965
rect 18604 27888 18656 27940
rect 5172 27820 5224 27872
rect 5448 27863 5500 27872
rect 5448 27829 5457 27863
rect 5457 27829 5491 27863
rect 5491 27829 5500 27863
rect 5448 27820 5500 27829
rect 6644 27863 6696 27872
rect 6644 27829 6653 27863
rect 6653 27829 6687 27863
rect 6687 27829 6696 27863
rect 6644 27820 6696 27829
rect 7288 27863 7340 27872
rect 7288 27829 7297 27863
rect 7297 27829 7331 27863
rect 7331 27829 7340 27863
rect 7288 27820 7340 27829
rect 8208 27820 8260 27872
rect 12256 27820 12308 27872
rect 16028 27820 16080 27872
rect 19248 27863 19300 27872
rect 19248 27829 19257 27863
rect 19257 27829 19291 27863
rect 19291 27829 19300 27863
rect 19248 27820 19300 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 4068 27659 4120 27668
rect 4068 27625 4077 27659
rect 4077 27625 4111 27659
rect 4111 27625 4120 27659
rect 4068 27616 4120 27625
rect 5172 27616 5224 27668
rect 8576 27616 8628 27668
rect 8760 27616 8812 27668
rect 1676 27591 1728 27600
rect 1676 27557 1685 27591
rect 1685 27557 1719 27591
rect 1719 27557 1728 27591
rect 1676 27548 1728 27557
rect 7196 27548 7248 27600
rect 12440 27548 12492 27600
rect 2412 27455 2464 27464
rect 2412 27421 2421 27455
rect 2421 27421 2455 27455
rect 2455 27421 2464 27455
rect 2412 27412 2464 27421
rect 2872 27412 2924 27464
rect 4896 27480 4948 27532
rect 5724 27412 5776 27464
rect 6828 27480 6880 27532
rect 3700 27344 3752 27396
rect 7656 27344 7708 27396
rect 5632 27276 5684 27328
rect 9312 27344 9364 27396
rect 9772 27387 9824 27396
rect 9772 27353 9781 27387
rect 9781 27353 9815 27387
rect 9815 27353 9824 27387
rect 10508 27480 10560 27532
rect 11244 27412 11296 27464
rect 12164 27412 12216 27464
rect 13728 27616 13780 27668
rect 18604 27659 18656 27668
rect 12624 27480 12676 27532
rect 13728 27480 13780 27532
rect 15752 27548 15804 27600
rect 15108 27480 15160 27532
rect 15292 27480 15344 27532
rect 15660 27480 15712 27532
rect 18052 27548 18104 27600
rect 16304 27480 16356 27532
rect 18604 27625 18613 27659
rect 18613 27625 18647 27659
rect 18647 27625 18656 27659
rect 18604 27616 18656 27625
rect 36360 27659 36412 27668
rect 36360 27625 36369 27659
rect 36369 27625 36403 27659
rect 36403 27625 36412 27659
rect 36360 27616 36412 27625
rect 14832 27455 14884 27464
rect 14832 27421 14841 27455
rect 14841 27421 14875 27455
rect 14875 27421 14884 27455
rect 14832 27412 14884 27421
rect 18604 27412 18656 27464
rect 19156 27480 19208 27532
rect 9772 27344 9824 27353
rect 10508 27344 10560 27396
rect 12624 27344 12676 27396
rect 12716 27344 12768 27396
rect 13084 27387 13136 27396
rect 13084 27353 13093 27387
rect 13093 27353 13127 27387
rect 13127 27353 13136 27387
rect 13084 27344 13136 27353
rect 12440 27276 12492 27328
rect 15660 27344 15712 27396
rect 16028 27387 16080 27396
rect 16028 27353 16037 27387
rect 16037 27353 16071 27387
rect 16071 27353 16080 27387
rect 16028 27344 16080 27353
rect 17224 27387 17276 27396
rect 14556 27276 14608 27328
rect 15200 27276 15252 27328
rect 17224 27353 17233 27387
rect 17233 27353 17267 27387
rect 17267 27353 17276 27387
rect 17224 27344 17276 27353
rect 36452 27412 36504 27464
rect 19156 27276 19208 27328
rect 24860 27276 24912 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 3332 27072 3384 27124
rect 4068 27072 4120 27124
rect 9496 27072 9548 27124
rect 9772 27072 9824 27124
rect 10508 27072 10560 27124
rect 14280 27072 14332 27124
rect 14556 27072 14608 27124
rect 15844 27072 15896 27124
rect 16304 27072 16356 27124
rect 18788 27115 18840 27124
rect 18788 27081 18797 27115
rect 18797 27081 18831 27115
rect 18831 27081 18840 27115
rect 18788 27072 18840 27081
rect 35992 27072 36044 27124
rect 6276 27004 6328 27056
rect 12716 27047 12768 27056
rect 1584 26979 1636 26988
rect 1584 26945 1593 26979
rect 1593 26945 1627 26979
rect 1627 26945 1636 26979
rect 1584 26936 1636 26945
rect 2136 26936 2188 26988
rect 9036 26979 9088 26988
rect 9036 26945 9045 26979
rect 9045 26945 9079 26979
rect 9079 26945 9088 26979
rect 9036 26936 9088 26945
rect 10508 26979 10560 26988
rect 10508 26945 10517 26979
rect 10517 26945 10551 26979
rect 10551 26945 10560 26979
rect 10508 26936 10560 26945
rect 6828 26868 6880 26920
rect 8576 26911 8628 26920
rect 8576 26877 8585 26911
rect 8585 26877 8619 26911
rect 8619 26877 8628 26911
rect 12440 26936 12492 26988
rect 12716 27013 12725 27047
rect 12725 27013 12759 27047
rect 12759 27013 12768 27047
rect 12716 27004 12768 27013
rect 13084 27004 13136 27056
rect 13728 27004 13780 27056
rect 14372 27047 14424 27056
rect 14372 27013 14381 27047
rect 14381 27013 14415 27047
rect 14415 27013 14424 27047
rect 14372 27004 14424 27013
rect 16120 27047 16172 27056
rect 16120 27013 16129 27047
rect 16129 27013 16163 27047
rect 16163 27013 16172 27047
rect 16120 27004 16172 27013
rect 17132 27004 17184 27056
rect 18420 27004 18472 27056
rect 14740 26936 14792 26988
rect 15016 26979 15068 26988
rect 15016 26945 15025 26979
rect 15025 26945 15059 26979
rect 15059 26945 15068 26979
rect 15016 26936 15068 26945
rect 16488 26936 16540 26988
rect 18604 26979 18656 26988
rect 8576 26868 8628 26877
rect 6736 26800 6788 26852
rect 9588 26800 9640 26852
rect 1768 26775 1820 26784
rect 1768 26741 1777 26775
rect 1777 26741 1811 26775
rect 1811 26741 1820 26775
rect 1768 26732 1820 26741
rect 5632 26732 5684 26784
rect 10876 26800 10928 26852
rect 12164 26800 12216 26852
rect 13268 26843 13320 26852
rect 13268 26809 13277 26843
rect 13277 26809 13311 26843
rect 13311 26809 13320 26843
rect 13268 26800 13320 26809
rect 15200 26800 15252 26852
rect 16212 26868 16264 26920
rect 18604 26945 18613 26979
rect 18613 26945 18647 26979
rect 18647 26945 18656 26979
rect 18604 26936 18656 26945
rect 19248 26936 19300 26988
rect 17500 26868 17552 26920
rect 16120 26800 16172 26852
rect 17868 26800 17920 26852
rect 26148 27004 26200 27056
rect 36360 26979 36412 26988
rect 36360 26945 36369 26979
rect 36369 26945 36403 26979
rect 36403 26945 36412 26979
rect 36360 26936 36412 26945
rect 10600 26732 10652 26784
rect 13544 26732 13596 26784
rect 13820 26732 13872 26784
rect 15476 26732 15528 26784
rect 15568 26732 15620 26784
rect 19248 26775 19300 26784
rect 19248 26741 19257 26775
rect 19257 26741 19291 26775
rect 19291 26741 19300 26775
rect 19248 26732 19300 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 1492 26528 1544 26580
rect 2228 26571 2280 26580
rect 2228 26537 2237 26571
rect 2237 26537 2271 26571
rect 2271 26537 2280 26571
rect 2228 26528 2280 26537
rect 6276 26571 6328 26580
rect 6276 26537 6285 26571
rect 6285 26537 6319 26571
rect 6319 26537 6328 26571
rect 6276 26528 6328 26537
rect 6368 26528 6420 26580
rect 8300 26528 8352 26580
rect 9312 26528 9364 26580
rect 1768 26460 1820 26512
rect 2596 26324 2648 26376
rect 6092 26256 6144 26308
rect 6828 26256 6880 26308
rect 7656 26299 7708 26308
rect 7656 26265 7665 26299
rect 7665 26265 7699 26299
rect 7699 26265 7708 26299
rect 7656 26256 7708 26265
rect 12532 26528 12584 26580
rect 9588 26460 9640 26512
rect 13268 26460 13320 26512
rect 15476 26460 15528 26512
rect 11428 26435 11480 26444
rect 11428 26401 11437 26435
rect 11437 26401 11471 26435
rect 11471 26401 11480 26435
rect 11428 26392 11480 26401
rect 12164 26392 12216 26444
rect 15292 26392 15344 26444
rect 15568 26435 15620 26444
rect 15568 26401 15577 26435
rect 15577 26401 15611 26435
rect 15611 26401 15620 26435
rect 15568 26392 15620 26401
rect 10416 26324 10468 26376
rect 10692 26367 10744 26376
rect 10692 26333 10701 26367
rect 10701 26333 10735 26367
rect 10735 26333 10744 26367
rect 10692 26324 10744 26333
rect 12716 26324 12768 26376
rect 12900 26324 12952 26376
rect 14832 26324 14884 26376
rect 16856 26460 16908 26512
rect 18236 26460 18288 26512
rect 9496 26256 9548 26308
rect 12992 26299 13044 26308
rect 12992 26265 13001 26299
rect 13001 26265 13035 26299
rect 13035 26265 13044 26299
rect 12992 26256 13044 26265
rect 13544 26299 13596 26308
rect 13544 26265 13553 26299
rect 13553 26265 13587 26299
rect 13587 26265 13596 26299
rect 13544 26256 13596 26265
rect 14004 26256 14056 26308
rect 16856 26256 16908 26308
rect 12532 26188 12584 26240
rect 15384 26188 15436 26240
rect 17316 26392 17368 26444
rect 17500 26435 17552 26444
rect 17500 26401 17509 26435
rect 17509 26401 17543 26435
rect 17543 26401 17552 26435
rect 17500 26392 17552 26401
rect 17960 26256 18012 26308
rect 18420 26299 18472 26308
rect 18420 26265 18429 26299
rect 18429 26265 18463 26299
rect 18463 26265 18472 26299
rect 18420 26256 18472 26265
rect 19248 26324 19300 26376
rect 32404 26324 32456 26376
rect 35532 26256 35584 26308
rect 19984 26231 20036 26240
rect 19984 26197 19993 26231
rect 19993 26197 20027 26231
rect 20027 26197 20036 26231
rect 19984 26188 20036 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 8300 25984 8352 26036
rect 10508 25984 10560 26036
rect 10968 25984 11020 26036
rect 17224 26027 17276 26036
rect 12164 25959 12216 25968
rect 12164 25925 12173 25959
rect 12173 25925 12207 25959
rect 12207 25925 12216 25959
rect 12164 25916 12216 25925
rect 15292 25959 15344 25968
rect 15292 25925 15301 25959
rect 15301 25925 15335 25959
rect 15335 25925 15344 25959
rect 15292 25916 15344 25925
rect 17224 25993 17233 26027
rect 17233 25993 17267 26027
rect 17267 25993 17276 26027
rect 17224 25984 17276 25993
rect 17868 26027 17920 26036
rect 17868 25993 17877 26027
rect 17877 25993 17911 26027
rect 17911 25993 17920 26027
rect 17868 25984 17920 25993
rect 10232 25891 10284 25900
rect 10232 25857 10241 25891
rect 10241 25857 10275 25891
rect 10275 25857 10284 25891
rect 10232 25848 10284 25857
rect 17960 25891 18012 25900
rect 10508 25780 10560 25832
rect 13176 25823 13228 25832
rect 12072 25712 12124 25764
rect 9772 25687 9824 25696
rect 9772 25653 9781 25687
rect 9781 25653 9815 25687
rect 9815 25653 9824 25687
rect 9772 25644 9824 25653
rect 11060 25687 11112 25696
rect 11060 25653 11069 25687
rect 11069 25653 11103 25687
rect 11103 25653 11112 25687
rect 11060 25644 11112 25653
rect 13176 25789 13185 25823
rect 13185 25789 13219 25823
rect 13219 25789 13228 25823
rect 13176 25780 13228 25789
rect 14004 25823 14056 25832
rect 14004 25789 14013 25823
rect 14013 25789 14047 25823
rect 14047 25789 14056 25823
rect 14004 25780 14056 25789
rect 14924 25780 14976 25832
rect 13636 25712 13688 25764
rect 17960 25857 17969 25891
rect 17969 25857 18003 25891
rect 18003 25857 18012 25891
rect 17960 25848 18012 25857
rect 19984 25848 20036 25900
rect 16948 25644 17000 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 13084 25440 13136 25492
rect 14648 25440 14700 25492
rect 18236 25483 18288 25492
rect 11796 25372 11848 25424
rect 15200 25415 15252 25424
rect 15200 25381 15209 25415
rect 15209 25381 15243 25415
rect 15243 25381 15252 25415
rect 15200 25372 15252 25381
rect 13452 25304 13504 25356
rect 17868 25304 17920 25356
rect 18236 25449 18245 25483
rect 18245 25449 18279 25483
rect 18279 25449 18288 25483
rect 18236 25440 18288 25449
rect 1584 25279 1636 25288
rect 1584 25245 1593 25279
rect 1593 25245 1627 25279
rect 1627 25245 1636 25279
rect 1584 25236 1636 25245
rect 10140 25236 10192 25288
rect 10876 25236 10928 25288
rect 7932 25168 7984 25220
rect 9312 25211 9364 25220
rect 9312 25177 9321 25211
rect 9321 25177 9355 25211
rect 9355 25177 9364 25211
rect 9312 25168 9364 25177
rect 11244 25168 11296 25220
rect 11612 25211 11664 25220
rect 11612 25177 11621 25211
rect 11621 25177 11655 25211
rect 11655 25177 11664 25211
rect 11612 25168 11664 25177
rect 12164 25211 12216 25220
rect 12164 25177 12173 25211
rect 12173 25177 12207 25211
rect 12207 25177 12216 25211
rect 12164 25168 12216 25177
rect 12624 25168 12676 25220
rect 13728 25168 13780 25220
rect 15016 25236 15068 25288
rect 18328 25279 18380 25288
rect 18328 25245 18337 25279
rect 18337 25245 18371 25279
rect 18371 25245 18380 25279
rect 18328 25236 18380 25245
rect 16856 25211 16908 25220
rect 1768 25143 1820 25152
rect 1768 25109 1777 25143
rect 1777 25109 1811 25143
rect 1811 25109 1820 25143
rect 1768 25100 1820 25109
rect 2504 25100 2556 25152
rect 9772 25100 9824 25152
rect 14372 25100 14424 25152
rect 16856 25177 16865 25211
rect 16865 25177 16899 25211
rect 16899 25177 16908 25211
rect 16856 25168 16908 25177
rect 17500 25168 17552 25220
rect 16580 25100 16632 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 9312 24896 9364 24948
rect 12532 24896 12584 24948
rect 15108 24896 15160 24948
rect 8392 24760 8444 24812
rect 8668 24760 8720 24812
rect 10140 24828 10192 24880
rect 10600 24871 10652 24880
rect 10600 24837 10609 24871
rect 10609 24837 10643 24871
rect 10643 24837 10652 24871
rect 10600 24828 10652 24837
rect 16580 24828 16632 24880
rect 10508 24735 10560 24744
rect 10508 24701 10517 24735
rect 10517 24701 10551 24735
rect 10551 24701 10560 24735
rect 10508 24692 10560 24701
rect 9680 24624 9732 24676
rect 11704 24692 11756 24744
rect 13176 24735 13228 24744
rect 13176 24701 13185 24735
rect 13185 24701 13219 24735
rect 13219 24701 13228 24735
rect 13176 24692 13228 24701
rect 14372 24760 14424 24812
rect 17868 24760 17920 24812
rect 25872 24803 25924 24812
rect 15844 24692 15896 24744
rect 16488 24692 16540 24744
rect 17500 24735 17552 24744
rect 17500 24701 17509 24735
rect 17509 24701 17543 24735
rect 17543 24701 17552 24735
rect 17500 24692 17552 24701
rect 12164 24556 12216 24608
rect 15752 24624 15804 24676
rect 25872 24769 25881 24803
rect 25881 24769 25915 24803
rect 25915 24769 25924 24803
rect 25872 24760 25924 24769
rect 33416 24803 33468 24812
rect 33416 24769 33425 24803
rect 33425 24769 33459 24803
rect 33459 24769 33468 24803
rect 33416 24760 33468 24769
rect 35532 24803 35584 24812
rect 35532 24769 35541 24803
rect 35541 24769 35575 24803
rect 35575 24769 35584 24803
rect 35532 24760 35584 24769
rect 22192 24624 22244 24676
rect 33600 24667 33652 24676
rect 13360 24556 13412 24608
rect 14832 24556 14884 24608
rect 16028 24556 16080 24608
rect 17868 24556 17920 24608
rect 24492 24556 24544 24608
rect 33600 24633 33609 24667
rect 33609 24633 33643 24667
rect 33643 24633 33652 24667
rect 33600 24624 33652 24633
rect 36084 24624 36136 24676
rect 35992 24556 36044 24608
rect 36268 24599 36320 24608
rect 36268 24565 36277 24599
rect 36277 24565 36311 24599
rect 36311 24565 36320 24599
rect 36268 24556 36320 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 11796 24352 11848 24404
rect 12348 24352 12400 24404
rect 15752 24352 15804 24404
rect 16856 24352 16908 24404
rect 17868 24352 17920 24404
rect 26148 24352 26200 24404
rect 12992 24284 13044 24336
rect 11152 24216 11204 24268
rect 11796 24216 11848 24268
rect 12072 24216 12124 24268
rect 12532 24216 12584 24268
rect 13452 24216 13504 24268
rect 12348 24191 12400 24200
rect 12348 24157 12357 24191
rect 12357 24157 12391 24191
rect 12391 24157 12400 24191
rect 12348 24148 12400 24157
rect 14924 24259 14976 24268
rect 14924 24225 14933 24259
rect 14933 24225 14967 24259
rect 14967 24225 14976 24259
rect 14924 24216 14976 24225
rect 15384 24216 15436 24268
rect 15844 24216 15896 24268
rect 7840 24123 7892 24132
rect 7840 24089 7849 24123
rect 7849 24089 7883 24123
rect 7883 24089 7892 24123
rect 7840 24080 7892 24089
rect 6644 24012 6696 24064
rect 8484 24123 8536 24132
rect 8484 24089 8493 24123
rect 8493 24089 8527 24123
rect 8527 24089 8536 24123
rect 8484 24080 8536 24089
rect 8944 24080 8996 24132
rect 9496 24123 9548 24132
rect 9496 24089 9505 24123
rect 9505 24089 9539 24123
rect 9539 24089 9548 24123
rect 9496 24080 9548 24089
rect 11244 24080 11296 24132
rect 11796 24080 11848 24132
rect 12808 24055 12860 24064
rect 12808 24021 12817 24055
rect 12817 24021 12851 24055
rect 12851 24021 12860 24055
rect 12808 24012 12860 24021
rect 14188 24080 14240 24132
rect 16028 24123 16080 24132
rect 16028 24089 16037 24123
rect 16037 24089 16071 24123
rect 16071 24089 16080 24123
rect 16028 24080 16080 24089
rect 16120 24123 16172 24132
rect 16120 24089 16129 24123
rect 16129 24089 16163 24123
rect 16163 24089 16172 24123
rect 25320 24216 25372 24268
rect 16948 24148 17000 24200
rect 17500 24191 17552 24200
rect 17500 24157 17509 24191
rect 17509 24157 17543 24191
rect 17543 24157 17552 24191
rect 17500 24148 17552 24157
rect 33416 24148 33468 24200
rect 16120 24080 16172 24089
rect 15384 24012 15436 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 7932 23808 7984 23860
rect 10876 23808 10928 23860
rect 11796 23808 11848 23860
rect 12348 23808 12400 23860
rect 16120 23808 16172 23860
rect 17500 23851 17552 23860
rect 17500 23817 17509 23851
rect 17509 23817 17543 23851
rect 17543 23817 17552 23851
rect 17500 23808 17552 23817
rect 36176 23808 36228 23860
rect 12256 23783 12308 23792
rect 12256 23749 12265 23783
rect 12265 23749 12299 23783
rect 12299 23749 12308 23783
rect 12256 23740 12308 23749
rect 13176 23783 13228 23792
rect 13176 23749 13185 23783
rect 13185 23749 13219 23783
rect 13219 23749 13228 23783
rect 13176 23740 13228 23749
rect 13820 23783 13872 23792
rect 13820 23749 13829 23783
rect 13829 23749 13863 23783
rect 13863 23749 13872 23783
rect 13820 23740 13872 23749
rect 15384 23783 15436 23792
rect 15384 23749 15393 23783
rect 15393 23749 15427 23783
rect 15427 23749 15436 23783
rect 15384 23740 15436 23749
rect 1860 23715 1912 23724
rect 1860 23681 1869 23715
rect 1869 23681 1903 23715
rect 1903 23681 1912 23715
rect 1860 23672 1912 23681
rect 2504 23715 2556 23724
rect 2504 23681 2513 23715
rect 2513 23681 2547 23715
rect 2547 23681 2556 23715
rect 2504 23672 2556 23681
rect 6552 23715 6604 23724
rect 6552 23681 6561 23715
rect 6561 23681 6595 23715
rect 6595 23681 6604 23715
rect 6552 23672 6604 23681
rect 10324 23715 10376 23724
rect 10324 23681 10333 23715
rect 10333 23681 10367 23715
rect 10367 23681 10376 23715
rect 10324 23672 10376 23681
rect 10692 23672 10744 23724
rect 10876 23672 10928 23724
rect 11980 23672 12032 23724
rect 22192 23672 22244 23724
rect 35900 23715 35952 23724
rect 35900 23681 35909 23715
rect 35909 23681 35943 23715
rect 35943 23681 35952 23715
rect 35900 23672 35952 23681
rect 12808 23604 12860 23656
rect 13728 23647 13780 23656
rect 13728 23613 13737 23647
rect 13737 23613 13771 23647
rect 13771 23613 13780 23647
rect 13728 23604 13780 23613
rect 11704 23536 11756 23588
rect 14188 23604 14240 23656
rect 15384 23604 15436 23656
rect 15476 23604 15528 23656
rect 1676 23511 1728 23520
rect 1676 23477 1685 23511
rect 1685 23477 1719 23511
rect 1719 23477 1728 23511
rect 1676 23468 1728 23477
rect 2320 23511 2372 23520
rect 2320 23477 2329 23511
rect 2329 23477 2363 23511
rect 2363 23477 2372 23511
rect 2320 23468 2372 23477
rect 35440 23468 35492 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 13820 23264 13872 23316
rect 11704 23239 11756 23248
rect 11704 23205 11713 23239
rect 11713 23205 11747 23239
rect 11747 23205 11756 23239
rect 11704 23196 11756 23205
rect 15200 23239 15252 23248
rect 15200 23205 15209 23239
rect 15209 23205 15243 23239
rect 15243 23205 15252 23239
rect 15200 23196 15252 23205
rect 6092 23103 6144 23112
rect 6092 23069 6101 23103
rect 6101 23069 6135 23103
rect 6135 23069 6144 23103
rect 6092 23060 6144 23069
rect 12348 23060 12400 23112
rect 12624 23060 12676 23112
rect 14188 23060 14240 23112
rect 16488 23128 16540 23180
rect 22192 23103 22244 23112
rect 22192 23069 22201 23103
rect 22201 23069 22235 23103
rect 22235 23069 22244 23103
rect 22192 23060 22244 23069
rect 35900 23060 35952 23112
rect 36452 23060 36504 23112
rect 11152 23035 11204 23044
rect 11152 23001 11161 23035
rect 11161 23001 11195 23035
rect 11195 23001 11204 23035
rect 11152 22992 11204 23001
rect 11520 22992 11572 23044
rect 15660 23035 15712 23044
rect 15660 23001 15669 23035
rect 15669 23001 15703 23035
rect 15703 23001 15712 23035
rect 15660 22992 15712 23001
rect 16488 22992 16540 23044
rect 6000 22967 6052 22976
rect 6000 22933 6009 22967
rect 6009 22933 6043 22967
rect 6043 22933 6052 22967
rect 6000 22924 6052 22933
rect 12808 22924 12860 22976
rect 13544 22924 13596 22976
rect 14740 22924 14792 22976
rect 35348 22924 35400 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 1860 22720 1912 22772
rect 8484 22720 8536 22772
rect 12348 22763 12400 22772
rect 8208 22695 8260 22704
rect 8208 22661 8217 22695
rect 8217 22661 8251 22695
rect 8251 22661 8260 22695
rect 8208 22652 8260 22661
rect 9036 22695 9088 22704
rect 9036 22661 9045 22695
rect 9045 22661 9079 22695
rect 9079 22661 9088 22695
rect 9036 22652 9088 22661
rect 10600 22695 10652 22704
rect 10600 22661 10609 22695
rect 10609 22661 10643 22695
rect 10643 22661 10652 22695
rect 10600 22652 10652 22661
rect 12348 22729 12357 22763
rect 12357 22729 12391 22763
rect 12391 22729 12400 22763
rect 12348 22720 12400 22729
rect 15660 22720 15712 22772
rect 11612 22652 11664 22704
rect 13544 22695 13596 22704
rect 13544 22661 13553 22695
rect 13553 22661 13587 22695
rect 13587 22661 13596 22695
rect 13544 22652 13596 22661
rect 14740 22695 14792 22704
rect 14740 22661 14749 22695
rect 14749 22661 14783 22695
rect 14783 22661 14792 22695
rect 14740 22652 14792 22661
rect 14832 22695 14884 22704
rect 14832 22661 14841 22695
rect 14841 22661 14875 22695
rect 14875 22661 14884 22695
rect 14832 22652 14884 22661
rect 15476 22652 15528 22704
rect 11980 22584 12032 22636
rect 12256 22627 12308 22636
rect 12256 22593 12265 22627
rect 12265 22593 12299 22627
rect 12299 22593 12308 22627
rect 12256 22584 12308 22593
rect 7472 22516 7524 22568
rect 7840 22559 7892 22568
rect 7840 22525 7849 22559
rect 7849 22525 7883 22559
rect 7883 22525 7892 22559
rect 7840 22516 7892 22525
rect 8300 22559 8352 22568
rect 8300 22525 8309 22559
rect 8309 22525 8343 22559
rect 8343 22525 8352 22559
rect 8300 22516 8352 22525
rect 8944 22559 8996 22568
rect 8944 22525 8953 22559
rect 8953 22525 8987 22559
rect 8987 22525 8996 22559
rect 8944 22516 8996 22525
rect 10508 22559 10560 22568
rect 10508 22525 10517 22559
rect 10517 22525 10551 22559
rect 10551 22525 10560 22559
rect 10508 22516 10560 22525
rect 10876 22516 10928 22568
rect 8392 22448 8444 22500
rect 15016 22448 15068 22500
rect 3240 22380 3292 22432
rect 6552 22380 6604 22432
rect 12624 22380 12676 22432
rect 18328 22584 18380 22636
rect 36084 22627 36136 22636
rect 36084 22593 36093 22627
rect 36093 22593 36127 22627
rect 36127 22593 36136 22627
rect 36084 22584 36136 22593
rect 36268 22491 36320 22500
rect 36268 22457 36277 22491
rect 36277 22457 36311 22491
rect 36311 22457 36320 22491
rect 36268 22448 36320 22457
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 9036 22176 9088 22228
rect 10600 22176 10652 22228
rect 11520 22219 11572 22228
rect 11520 22185 11529 22219
rect 11529 22185 11563 22219
rect 11563 22185 11572 22219
rect 11520 22176 11572 22185
rect 8300 22108 8352 22160
rect 8944 22040 8996 22092
rect 10324 22040 10376 22092
rect 9404 21972 9456 22024
rect 12716 22040 12768 22092
rect 14004 22040 14056 22092
rect 15200 22108 15252 22160
rect 15292 22040 15344 22092
rect 5908 21879 5960 21888
rect 5908 21845 5917 21879
rect 5917 21845 5951 21879
rect 5951 21845 5960 21879
rect 5908 21836 5960 21845
rect 6276 21836 6328 21888
rect 11980 21972 12032 22024
rect 14096 21972 14148 22024
rect 16212 22015 16264 22024
rect 16212 21981 16221 22015
rect 16221 21981 16255 22015
rect 16255 21981 16264 22015
rect 16212 21972 16264 21981
rect 13912 21904 13964 21956
rect 15292 21904 15344 21956
rect 14096 21836 14148 21888
rect 30564 21904 30616 21956
rect 31760 21879 31812 21888
rect 31760 21845 31769 21879
rect 31769 21845 31803 21879
rect 31803 21845 31812 21879
rect 31760 21836 31812 21845
rect 35900 21836 35952 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 12624 21675 12676 21684
rect 12624 21641 12633 21675
rect 12633 21641 12667 21675
rect 12667 21641 12676 21675
rect 12624 21632 12676 21641
rect 13728 21632 13780 21684
rect 7288 21564 7340 21616
rect 11980 21564 12032 21616
rect 27160 21632 27212 21684
rect 2320 21496 2372 21548
rect 12992 21496 13044 21548
rect 13820 21539 13872 21548
rect 13820 21505 13829 21539
rect 13829 21505 13863 21539
rect 13863 21505 13872 21539
rect 13820 21496 13872 21505
rect 35992 21496 36044 21548
rect 7288 21428 7340 21480
rect 8208 21428 8260 21480
rect 14740 21428 14792 21480
rect 15752 21471 15804 21480
rect 15752 21437 15761 21471
rect 15761 21437 15795 21471
rect 15795 21437 15804 21471
rect 15752 21428 15804 21437
rect 15200 21403 15252 21412
rect 15200 21369 15209 21403
rect 15209 21369 15243 21403
rect 15243 21369 15252 21403
rect 15200 21360 15252 21369
rect 1676 21335 1728 21344
rect 1676 21301 1685 21335
rect 1685 21301 1719 21335
rect 1719 21301 1728 21335
rect 1676 21292 1728 21301
rect 11980 21292 12032 21344
rect 36268 21335 36320 21344
rect 36268 21301 36277 21335
rect 36277 21301 36311 21335
rect 36311 21301 36320 21335
rect 36268 21292 36320 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 12256 21088 12308 21140
rect 12992 21088 13044 21140
rect 25412 21088 25464 21140
rect 30564 21131 30616 21140
rect 30564 21097 30573 21131
rect 30573 21097 30607 21131
rect 30607 21097 30616 21131
rect 30564 21088 30616 21097
rect 36084 21131 36136 21140
rect 36084 21097 36093 21131
rect 36093 21097 36127 21131
rect 36127 21097 36136 21131
rect 36084 21088 36136 21097
rect 13820 21020 13872 21072
rect 14740 20995 14792 21004
rect 14740 20961 14749 20995
rect 14749 20961 14783 20995
rect 14783 20961 14792 20995
rect 14740 20952 14792 20961
rect 35716 20884 35768 20936
rect 14832 20859 14884 20868
rect 14832 20825 14841 20859
rect 14841 20825 14875 20859
rect 14875 20825 14884 20859
rect 14832 20816 14884 20825
rect 16396 20816 16448 20868
rect 12992 20791 13044 20800
rect 12992 20757 13001 20791
rect 13001 20757 13035 20791
rect 13035 20757 13044 20791
rect 12992 20748 13044 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 14832 20544 14884 20596
rect 16212 20587 16264 20596
rect 16212 20553 16221 20587
rect 16221 20553 16255 20587
rect 16255 20553 16264 20587
rect 16212 20544 16264 20553
rect 13820 20408 13872 20460
rect 16948 20272 17000 20324
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 5264 20000 5316 20052
rect 8392 20000 8444 20052
rect 11152 20000 11204 20052
rect 21824 20043 21876 20052
rect 21824 20009 21833 20043
rect 21833 20009 21867 20043
rect 21867 20009 21876 20043
rect 21824 20000 21876 20009
rect 6000 19728 6052 19780
rect 6184 19728 6236 19780
rect 21824 19796 21876 19848
rect 1676 19703 1728 19712
rect 1676 19669 1685 19703
rect 1685 19669 1719 19703
rect 1719 19669 1728 19703
rect 1676 19660 1728 19669
rect 1952 19660 2004 19712
rect 7564 19703 7616 19712
rect 7564 19669 7573 19703
rect 7573 19669 7607 19703
rect 7607 19669 7616 19703
rect 7564 19660 7616 19669
rect 20812 19660 20864 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 2504 18819 2556 18828
rect 2504 18785 2513 18819
rect 2513 18785 2547 18819
rect 2547 18785 2556 18819
rect 2504 18776 2556 18785
rect 8208 18776 8260 18828
rect 16396 18819 16448 18828
rect 16396 18785 16405 18819
rect 16405 18785 16439 18819
rect 16439 18785 16448 18819
rect 16396 18776 16448 18785
rect 7564 18683 7616 18692
rect 7564 18649 7573 18683
rect 7573 18649 7607 18683
rect 7607 18649 7616 18683
rect 16948 18683 17000 18692
rect 7564 18640 7616 18649
rect 16948 18649 16957 18683
rect 16957 18649 16991 18683
rect 16991 18649 17000 18683
rect 16948 18640 17000 18649
rect 1768 18615 1820 18624
rect 1768 18581 1777 18615
rect 1777 18581 1811 18615
rect 1811 18581 1820 18615
rect 1768 18572 1820 18581
rect 7380 18572 7432 18624
rect 17684 18615 17736 18624
rect 17684 18581 17693 18615
rect 17693 18581 17727 18615
rect 17727 18581 17736 18615
rect 17684 18572 17736 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 1584 18232 1636 18284
rect 12992 18028 13044 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 1584 17799 1636 17808
rect 1584 17765 1593 17799
rect 1593 17765 1627 17799
rect 1627 17765 1636 17799
rect 1584 17756 1636 17765
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 27160 17187 27212 17196
rect 27160 17153 27169 17187
rect 27169 17153 27203 17187
rect 27203 17153 27212 17187
rect 27160 17144 27212 17153
rect 36268 17051 36320 17060
rect 36268 17017 36277 17051
rect 36277 17017 36311 17051
rect 36311 17017 36320 17051
rect 36268 17008 36320 17017
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 14096 16056 14148 16108
rect 25412 16099 25464 16108
rect 25412 16065 25421 16099
rect 25421 16065 25455 16099
rect 25455 16065 25464 16099
rect 25412 16056 25464 16065
rect 36176 16056 36228 16108
rect 36360 16031 36412 16040
rect 36360 15997 36369 16031
rect 36369 15997 36403 16031
rect 36403 15997 36412 16031
rect 36360 15988 36412 15997
rect 34152 15920 34204 15972
rect 1676 15895 1728 15904
rect 1676 15861 1685 15895
rect 1685 15861 1719 15895
rect 1719 15861 1728 15895
rect 1676 15852 1728 15861
rect 25596 15895 25648 15904
rect 25596 15861 25605 15895
rect 25605 15861 25639 15895
rect 25639 15861 25648 15895
rect 25596 15852 25648 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 25596 15648 25648 15700
rect 34520 15648 34572 15700
rect 36360 15691 36412 15700
rect 36360 15657 36369 15691
rect 36369 15657 36403 15691
rect 36403 15657 36412 15691
rect 36360 15648 36412 15657
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 24860 14399 24912 14408
rect 24860 14365 24869 14399
rect 24869 14365 24903 14399
rect 24903 14365 24912 14399
rect 24860 14356 24912 14365
rect 36176 14356 36228 14408
rect 1676 14331 1728 14340
rect 1676 14297 1685 14331
rect 1685 14297 1719 14331
rect 1719 14297 1728 14331
rect 1676 14288 1728 14297
rect 6184 14288 6236 14340
rect 17684 14288 17736 14340
rect 25044 14263 25096 14272
rect 25044 14229 25053 14263
rect 25053 14229 25087 14263
rect 25087 14229 25096 14263
rect 25044 14220 25096 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 1676 14059 1728 14068
rect 1676 14025 1685 14059
rect 1685 14025 1719 14059
rect 1719 14025 1728 14059
rect 1676 14016 1728 14025
rect 13084 14016 13136 14068
rect 13452 13880 13504 13932
rect 34520 13880 34572 13932
rect 36268 13719 36320 13728
rect 36268 13685 36277 13719
rect 36277 13685 36311 13719
rect 36311 13685 36320 13719
rect 36268 13676 36320 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 7288 13268 7340 13320
rect 1860 13175 1912 13184
rect 1860 13141 1869 13175
rect 1869 13141 1903 13175
rect 1903 13141 1912 13175
rect 1860 13132 1912 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 1860 12835 1912 12844
rect 1860 12801 1869 12835
rect 1869 12801 1903 12835
rect 1903 12801 1912 12835
rect 1860 12792 1912 12801
rect 1676 12631 1728 12640
rect 1676 12597 1685 12631
rect 1685 12597 1719 12631
rect 1719 12597 1728 12631
rect 1676 12588 1728 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 36360 11747 36412 11756
rect 36360 11713 36369 11747
rect 36369 11713 36403 11747
rect 36403 11713 36412 11747
rect 36360 11704 36412 11713
rect 36176 11543 36228 11552
rect 36176 11509 36185 11543
rect 36185 11509 36219 11543
rect 36219 11509 36228 11543
rect 36176 11500 36228 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 1952 10616 2004 10668
rect 36452 10616 36504 10668
rect 36360 10591 36412 10600
rect 36360 10557 36369 10591
rect 36369 10557 36403 10591
rect 36403 10557 36412 10591
rect 36360 10548 36412 10557
rect 1676 10455 1728 10464
rect 1676 10421 1685 10455
rect 1685 10421 1719 10455
rect 1719 10421 1728 10455
rect 1676 10412 1728 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 36360 10251 36412 10260
rect 36360 10217 36369 10251
rect 36369 10217 36403 10251
rect 36403 10217 36412 10251
rect 36360 10208 36412 10217
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 7380 9596 7432 9648
rect 2780 9528 2832 9580
rect 13176 9324 13228 9376
rect 36084 9367 36136 9376
rect 36084 9333 36093 9367
rect 36093 9333 36127 9367
rect 36127 9333 36136 9367
rect 36084 9324 36136 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 6276 8984 6328 9036
rect 1584 8959 1636 8968
rect 1584 8925 1593 8959
rect 1593 8925 1627 8959
rect 1627 8925 1636 8959
rect 1584 8916 1636 8925
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 10876 8619 10928 8628
rect 10876 8585 10885 8619
rect 10885 8585 10919 8619
rect 10919 8585 10928 8619
rect 10876 8576 10928 8585
rect 15384 8576 15436 8628
rect 24492 8619 24544 8628
rect 24492 8585 24501 8619
rect 24501 8585 24535 8619
rect 24535 8585 24544 8619
rect 24492 8576 24544 8585
rect 10968 8483 11020 8492
rect 10968 8449 10977 8483
rect 10977 8449 11011 8483
rect 11011 8449 11020 8483
rect 10968 8440 11020 8449
rect 15108 8483 15160 8492
rect 15108 8449 15117 8483
rect 15117 8449 15151 8483
rect 15151 8449 15160 8483
rect 15108 8440 15160 8449
rect 30012 8440 30064 8492
rect 36176 8508 36228 8560
rect 36084 8483 36136 8492
rect 36084 8449 36093 8483
rect 36093 8449 36127 8483
rect 36127 8449 36136 8483
rect 36084 8440 36136 8449
rect 36084 8304 36136 8356
rect 36268 8347 36320 8356
rect 36268 8313 36277 8347
rect 36277 8313 36311 8347
rect 36311 8313 36320 8347
rect 36268 8304 36320 8313
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 15752 8075 15804 8084
rect 15752 8041 15761 8075
rect 15761 8041 15795 8075
rect 15795 8041 15804 8075
rect 15752 8032 15804 8041
rect 15844 7871 15896 7880
rect 15844 7837 15853 7871
rect 15853 7837 15887 7871
rect 15887 7837 15896 7871
rect 15844 7828 15896 7837
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 1860 7395 1912 7404
rect 1860 7361 1869 7395
rect 1869 7361 1903 7395
rect 1903 7361 1912 7395
rect 1860 7352 1912 7361
rect 1676 7191 1728 7200
rect 1676 7157 1685 7191
rect 1685 7157 1719 7191
rect 1719 7157 1728 7191
rect 1676 7148 1728 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 6368 6783 6420 6792
rect 6368 6749 6377 6783
rect 6377 6749 6411 6783
rect 6411 6749 6420 6783
rect 6368 6740 6420 6749
rect 6552 6647 6604 6656
rect 6552 6613 6561 6647
rect 6561 6613 6595 6647
rect 6595 6613 6604 6647
rect 6552 6604 6604 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 15016 6443 15068 6452
rect 15016 6409 15025 6443
rect 15025 6409 15059 6443
rect 15059 6409 15068 6443
rect 15016 6400 15068 6409
rect 35900 6400 35952 6452
rect 15568 6307 15620 6316
rect 15568 6273 15577 6307
rect 15577 6273 15611 6307
rect 15611 6273 15620 6307
rect 15568 6264 15620 6273
rect 36360 6307 36412 6316
rect 36360 6273 36369 6307
rect 36369 6273 36403 6307
rect 36403 6273 36412 6307
rect 36360 6264 36412 6273
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 1584 5219 1636 5228
rect 1584 5185 1593 5219
rect 1593 5185 1627 5219
rect 1627 5185 1636 5219
rect 1584 5176 1636 5185
rect 36084 5219 36136 5228
rect 36084 5185 36093 5219
rect 36093 5185 36127 5219
rect 36127 5185 36136 5219
rect 36084 5176 36136 5185
rect 2780 4972 2832 5024
rect 3976 4972 4028 5024
rect 36268 5015 36320 5024
rect 36268 4981 36277 5015
rect 36277 4981 36311 5015
rect 36311 4981 36320 5015
rect 36268 4972 36320 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 36360 3927 36412 3936
rect 36360 3893 36369 3927
rect 36369 3893 36403 3927
rect 36403 3893 36412 3927
rect 36360 3884 36412 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 1860 3680 1912 3732
rect 15568 3723 15620 3732
rect 15568 3689 15577 3723
rect 15577 3689 15611 3723
rect 15611 3689 15620 3723
rect 15568 3680 15620 3689
rect 2504 3519 2556 3528
rect 2504 3485 2513 3519
rect 2513 3485 2547 3519
rect 2547 3485 2556 3519
rect 2504 3476 2556 3485
rect 15568 3476 15620 3528
rect 11704 3408 11756 3460
rect 34888 3408 34940 3460
rect 1676 3383 1728 3392
rect 1676 3349 1685 3383
rect 1685 3349 1719 3383
rect 1719 3349 1728 3383
rect 1676 3340 1728 3349
rect 14924 3383 14976 3392
rect 14924 3349 14933 3383
rect 14933 3349 14967 3383
rect 14967 3349 14976 3383
rect 14924 3340 14976 3349
rect 33140 3340 33192 3392
rect 36268 3383 36320 3392
rect 36268 3349 36277 3383
rect 36277 3349 36311 3383
rect 36311 3349 36320 3383
rect 36268 3340 36320 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 11704 3179 11756 3188
rect 11704 3145 11713 3179
rect 11713 3145 11747 3179
rect 11747 3145 11756 3179
rect 11704 3136 11756 3145
rect 3976 3043 4028 3052
rect 3976 3009 3985 3043
rect 3985 3009 4019 3043
rect 4019 3009 4028 3043
rect 3976 3000 4028 3009
rect 15108 3136 15160 3188
rect 14464 3111 14516 3120
rect 14464 3077 14473 3111
rect 14473 3077 14507 3111
rect 14507 3077 14516 3111
rect 14464 3068 14516 3077
rect 17132 3068 17184 3120
rect 15844 3043 15896 3052
rect 15844 3009 15853 3043
rect 15853 3009 15887 3043
rect 15887 3009 15896 3043
rect 15844 3000 15896 3009
rect 19340 3043 19392 3052
rect 19340 3009 19349 3043
rect 19349 3009 19383 3043
rect 19383 3009 19392 3043
rect 19340 3000 19392 3009
rect 30012 3000 30064 3052
rect 14924 2932 14976 2984
rect 24676 2932 24728 2984
rect 10968 2864 11020 2916
rect 14464 2864 14516 2916
rect 33140 2864 33192 2916
rect 34888 3000 34940 3052
rect 36360 2975 36412 2984
rect 36360 2941 36369 2975
rect 36369 2941 36403 2975
rect 36403 2941 36412 2975
rect 36360 2932 36412 2941
rect 37372 2932 37424 2984
rect 1676 2839 1728 2848
rect 1676 2805 1685 2839
rect 1685 2805 1719 2839
rect 1719 2805 1728 2839
rect 1676 2796 1728 2805
rect 2320 2839 2372 2848
rect 2320 2805 2329 2839
rect 2329 2805 2363 2839
rect 2363 2805 2372 2839
rect 2320 2796 2372 2805
rect 4620 2796 4672 2848
rect 10232 2839 10284 2848
rect 10232 2805 10241 2839
rect 10241 2805 10275 2839
rect 10275 2805 10284 2839
rect 10232 2796 10284 2805
rect 15200 2796 15252 2848
rect 22008 2796 22060 2848
rect 32220 2796 32272 2848
rect 36544 2796 36596 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 2504 2635 2556 2644
rect 2504 2601 2513 2635
rect 2513 2601 2547 2635
rect 2547 2601 2556 2635
rect 2504 2592 2556 2601
rect 3240 2635 3292 2644
rect 3240 2601 3249 2635
rect 3249 2601 3283 2635
rect 3283 2601 3292 2635
rect 3240 2592 3292 2601
rect 11060 2592 11112 2644
rect 11980 2524 12032 2576
rect 14188 2524 14240 2576
rect 15844 2592 15896 2644
rect 20812 2635 20864 2644
rect 20812 2601 20821 2635
rect 20821 2601 20855 2635
rect 20855 2601 20864 2635
rect 20812 2592 20864 2601
rect 22192 2635 22244 2644
rect 22192 2601 22201 2635
rect 22201 2601 22235 2635
rect 22235 2601 22244 2635
rect 22192 2592 22244 2601
rect 25044 2592 25096 2644
rect 32404 2635 32456 2644
rect 10968 2456 11020 2508
rect 1768 2388 1820 2440
rect 2320 2431 2372 2440
rect 2320 2397 2329 2431
rect 2329 2397 2363 2431
rect 2363 2397 2372 2431
rect 2320 2388 2372 2397
rect 4620 2431 4672 2440
rect 4620 2397 4629 2431
rect 4629 2397 4663 2431
rect 4663 2397 4672 2431
rect 4620 2388 4672 2397
rect 6552 2431 6604 2440
rect 6552 2397 6561 2431
rect 6561 2397 6595 2431
rect 6595 2397 6604 2431
rect 6552 2388 6604 2397
rect 3240 2320 3292 2372
rect 1308 2252 1360 2304
rect 4528 2252 4580 2304
rect 6460 2252 6512 2304
rect 8392 2252 8444 2304
rect 13084 2388 13136 2440
rect 15200 2431 15252 2440
rect 15200 2397 15209 2431
rect 15209 2397 15243 2431
rect 15243 2397 15252 2431
rect 15200 2388 15252 2397
rect 22008 2524 22060 2576
rect 9680 2320 9732 2372
rect 10232 2320 10284 2372
rect 13544 2363 13596 2372
rect 13544 2329 13553 2363
rect 13553 2329 13587 2363
rect 13587 2329 13596 2363
rect 13544 2320 13596 2329
rect 15108 2320 15160 2372
rect 11612 2252 11664 2304
rect 14832 2252 14884 2304
rect 16764 2252 16816 2304
rect 18696 2252 18748 2304
rect 20812 2388 20864 2440
rect 30012 2499 30064 2508
rect 30012 2465 30021 2499
rect 30021 2465 30055 2499
rect 30055 2465 30064 2499
rect 30012 2456 30064 2465
rect 32404 2601 32413 2635
rect 32413 2601 32447 2635
rect 32447 2601 32456 2635
rect 32404 2592 32456 2601
rect 34152 2635 34204 2644
rect 34152 2601 34161 2635
rect 34161 2601 34195 2635
rect 34195 2601 34204 2635
rect 34152 2592 34204 2601
rect 35716 2456 35768 2508
rect 21916 2320 21968 2372
rect 19984 2252 20036 2304
rect 23848 2252 23900 2304
rect 24676 2320 24728 2372
rect 25136 2252 25188 2304
rect 27068 2252 27120 2304
rect 29000 2252 29052 2304
rect 35440 2388 35492 2440
rect 32220 2320 32272 2372
rect 34152 2320 34204 2372
rect 30288 2252 30340 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 20 1300 72 1352
rect 2320 1300 2372 1352
<< metal2 >>
rect 662 39200 718 39800
rect 2594 39200 2650 39800
rect 3422 39536 3478 39545
rect 3422 39471 3478 39480
rect 676 37670 704 39200
rect 664 37664 716 37670
rect 664 37606 716 37612
rect 1768 37188 1820 37194
rect 1688 37148 1768 37176
rect 1584 37120 1636 37126
rect 1584 37062 1636 37068
rect 1596 36242 1624 37062
rect 1584 36236 1636 36242
rect 1584 36178 1636 36184
rect 1596 35698 1624 36178
rect 1584 35692 1636 35698
rect 1584 35634 1636 35640
rect 1584 34944 1636 34950
rect 1688 34932 1716 37148
rect 1768 37130 1820 37136
rect 2608 37126 2636 39200
rect 3436 37330 3464 39471
rect 4526 39200 4582 39800
rect 5814 39200 5870 39800
rect 7746 39200 7802 39800
rect 9678 39200 9734 39800
rect 10966 39200 11022 39800
rect 12898 39200 12954 39800
rect 14830 39200 14886 39800
rect 16118 39200 16174 39800
rect 16224 39222 16620 39250
rect 4540 37754 4568 39200
rect 4540 37726 4660 37754
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 3424 37324 3476 37330
rect 3424 37266 3476 37272
rect 4528 37324 4580 37330
rect 4528 37266 4580 37272
rect 3148 37188 3200 37194
rect 3148 37130 3200 37136
rect 2596 37120 2648 37126
rect 2596 37062 2648 37068
rect 2608 36786 2636 37062
rect 2964 36848 3016 36854
rect 2964 36790 3016 36796
rect 2228 36780 2280 36786
rect 2228 36722 2280 36728
rect 2596 36780 2648 36786
rect 2596 36722 2648 36728
rect 2240 36378 2268 36722
rect 2228 36372 2280 36378
rect 2228 36314 2280 36320
rect 2412 36236 2464 36242
rect 2412 36178 2464 36184
rect 1768 35284 1820 35290
rect 1768 35226 1820 35232
rect 1636 34904 1716 34932
rect 1584 34886 1636 34892
rect 1596 33114 1624 34886
rect 1780 34610 1808 35226
rect 2424 34746 2452 36178
rect 2608 35630 2636 36722
rect 2596 35624 2648 35630
rect 2596 35566 2648 35572
rect 2608 35154 2636 35566
rect 2976 35494 3004 36790
rect 3160 36582 3188 37130
rect 3332 37120 3384 37126
rect 3332 37062 3384 37068
rect 3148 36576 3200 36582
rect 3148 36518 3200 36524
rect 3344 35834 3372 37062
rect 4540 36666 4568 37266
rect 4632 36922 4660 37726
rect 5172 37664 5224 37670
rect 5172 37606 5224 37612
rect 4620 36916 4672 36922
rect 4620 36858 4672 36864
rect 4712 36712 4764 36718
rect 4540 36638 4660 36666
rect 4712 36654 4764 36660
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4066 36136 4122 36145
rect 4066 36071 4122 36080
rect 4080 36038 4108 36071
rect 4068 36032 4120 36038
rect 4068 35974 4120 35980
rect 3332 35828 3384 35834
rect 3332 35770 3384 35776
rect 3792 35828 3844 35834
rect 3792 35770 3844 35776
rect 2964 35488 3016 35494
rect 2964 35430 3016 35436
rect 2596 35148 2648 35154
rect 2596 35090 2648 35096
rect 2608 34762 2636 35090
rect 2516 34746 2728 34762
rect 2412 34740 2464 34746
rect 2412 34682 2464 34688
rect 2516 34740 2740 34746
rect 2516 34734 2688 34740
rect 1768 34604 1820 34610
rect 1768 34546 1820 34552
rect 2228 33856 2280 33862
rect 2228 33798 2280 33804
rect 2240 33658 2268 33798
rect 2228 33652 2280 33658
rect 2228 33594 2280 33600
rect 1676 33516 1728 33522
rect 1676 33458 1728 33464
rect 1584 33108 1636 33114
rect 1584 33050 1636 33056
rect 1688 32978 1716 33458
rect 2240 33454 2268 33594
rect 2228 33448 2280 33454
rect 2228 33390 2280 33396
rect 2424 33402 2452 34682
rect 2516 33590 2544 34734
rect 2688 34682 2740 34688
rect 3240 34672 3292 34678
rect 3240 34614 3292 34620
rect 3700 34672 3752 34678
rect 3700 34614 3752 34620
rect 2504 33584 2556 33590
rect 2504 33526 2556 33532
rect 2424 33374 2544 33402
rect 1676 32972 1728 32978
rect 1676 32914 1728 32920
rect 1688 32570 1716 32914
rect 1676 32564 1728 32570
rect 1676 32506 1728 32512
rect 1952 32564 2004 32570
rect 1952 32506 2004 32512
rect 1676 32428 1728 32434
rect 1676 32370 1728 32376
rect 1490 30696 1546 30705
rect 1490 30631 1492 30640
rect 1544 30631 1546 30640
rect 1492 30602 1544 30608
rect 1504 26586 1532 30602
rect 1688 29850 1716 32370
rect 1964 31346 1992 32506
rect 2412 32428 2464 32434
rect 2412 32370 2464 32376
rect 2226 32056 2282 32065
rect 2226 31991 2282 32000
rect 2240 31890 2268 31991
rect 2228 31884 2280 31890
rect 2228 31826 2280 31832
rect 2136 31816 2188 31822
rect 2136 31758 2188 31764
rect 1952 31340 2004 31346
rect 1952 31282 2004 31288
rect 1964 30326 1992 31282
rect 1952 30320 2004 30326
rect 1952 30262 2004 30268
rect 1676 29844 1728 29850
rect 1676 29786 1728 29792
rect 1584 29096 1636 29102
rect 1584 29038 1636 29044
rect 1596 28665 1624 29038
rect 1582 28656 1638 28665
rect 1582 28591 1638 28600
rect 1596 27962 1624 28591
rect 1676 28416 1728 28422
rect 1676 28358 1728 28364
rect 1688 28150 1716 28358
rect 1676 28144 1728 28150
rect 1676 28086 1728 28092
rect 1596 27934 1716 27962
rect 1584 27872 1636 27878
rect 1584 27814 1636 27820
rect 1596 26994 1624 27814
rect 1688 27606 1716 27934
rect 2148 27878 2176 31758
rect 2136 27872 2188 27878
rect 2136 27814 2188 27820
rect 1676 27600 1728 27606
rect 1676 27542 1728 27548
rect 2148 26994 2176 27814
rect 1584 26988 1636 26994
rect 1584 26930 1636 26936
rect 2136 26988 2188 26994
rect 2136 26930 2188 26936
rect 1768 26784 1820 26790
rect 1768 26726 1820 26732
rect 1780 26625 1808 26726
rect 1766 26616 1822 26625
rect 1492 26580 1544 26586
rect 2240 26586 2268 31826
rect 2424 30734 2452 32370
rect 2412 30728 2464 30734
rect 2412 30670 2464 30676
rect 2320 30320 2372 30326
rect 2320 30262 2372 30268
rect 2332 29850 2360 30262
rect 2320 29844 2372 29850
rect 2320 29786 2372 29792
rect 2424 29646 2452 30670
rect 2412 29640 2464 29646
rect 2412 29582 2464 29588
rect 2424 28082 2452 29582
rect 2516 28626 2544 33374
rect 2596 32292 2648 32298
rect 2596 32234 2648 32240
rect 2608 31278 2636 32234
rect 3252 32026 3280 34614
rect 3608 33584 3660 33590
rect 3608 33526 3660 33532
rect 3332 32904 3384 32910
rect 3332 32846 3384 32852
rect 3240 32020 3292 32026
rect 3240 31962 3292 31968
rect 2964 31816 3016 31822
rect 2964 31758 3016 31764
rect 2596 31272 2648 31278
rect 2596 31214 2648 31220
rect 2504 28620 2556 28626
rect 2504 28562 2556 28568
rect 2412 28076 2464 28082
rect 2412 28018 2464 28024
rect 2424 27470 2452 28018
rect 2412 27464 2464 27470
rect 2412 27406 2464 27412
rect 1766 26551 1822 26560
rect 2228 26580 2280 26586
rect 1492 26522 1544 26528
rect 2228 26522 2280 26528
rect 1768 26512 1820 26518
rect 1768 26454 1820 26460
rect 1584 25288 1636 25294
rect 1582 25256 1584 25265
rect 1636 25256 1638 25265
rect 1582 25191 1638 25200
rect 1780 25158 1808 26454
rect 2608 26382 2636 31214
rect 2976 30734 3004 31758
rect 2964 30728 3016 30734
rect 2964 30670 3016 30676
rect 2976 29714 3004 30670
rect 3056 30592 3108 30598
rect 3056 30534 3108 30540
rect 2964 29708 3016 29714
rect 2964 29650 3016 29656
rect 2976 28948 3004 29650
rect 3068 29238 3096 30534
rect 3148 30184 3200 30190
rect 3148 30126 3200 30132
rect 3160 29306 3188 30126
rect 3240 30048 3292 30054
rect 3240 29990 3292 29996
rect 3148 29300 3200 29306
rect 3148 29242 3200 29248
rect 3056 29232 3108 29238
rect 3056 29174 3108 29180
rect 2884 28920 3004 28948
rect 2884 28558 2912 28920
rect 2872 28552 2924 28558
rect 2872 28494 2924 28500
rect 2872 28416 2924 28422
rect 2872 28358 2924 28364
rect 2884 28082 2912 28358
rect 3252 28218 3280 29990
rect 3240 28212 3292 28218
rect 3240 28154 3292 28160
rect 2872 28076 2924 28082
rect 2872 28018 2924 28024
rect 2884 27470 2912 28018
rect 2872 27464 2924 27470
rect 2872 27406 2924 27412
rect 3344 27130 3372 32846
rect 3620 29782 3648 33526
rect 3712 33454 3740 34614
rect 3700 33448 3752 33454
rect 3700 33390 3752 33396
rect 3700 32768 3752 32774
rect 3700 32710 3752 32716
rect 3712 32366 3740 32710
rect 3700 32360 3752 32366
rect 3700 32302 3752 32308
rect 3712 31890 3740 32302
rect 3804 31929 3832 35770
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 3884 35148 3936 35154
rect 3884 35090 3936 35096
rect 3896 32586 3924 35090
rect 4068 35012 4120 35018
rect 4068 34954 4120 34960
rect 3976 34604 4028 34610
rect 3976 34546 4028 34552
rect 3988 34202 4016 34546
rect 3976 34196 4028 34202
rect 3976 34138 4028 34144
rect 4080 34082 4108 34954
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4080 34054 4200 34082
rect 4172 33318 4200 34054
rect 4160 33312 4212 33318
rect 4160 33254 4212 33260
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4632 32994 4660 36638
rect 4724 35630 4752 36654
rect 4896 36644 4948 36650
rect 4896 36586 4948 36592
rect 4712 35624 4764 35630
rect 4712 35566 4764 35572
rect 4712 35012 4764 35018
rect 4712 34954 4764 34960
rect 4540 32966 4660 32994
rect 4540 32774 4568 32966
rect 4620 32836 4672 32842
rect 4620 32778 4672 32784
rect 4528 32768 4580 32774
rect 4528 32710 4580 32716
rect 3896 32558 4200 32586
rect 3790 31920 3846 31929
rect 3700 31884 3752 31890
rect 3790 31855 3846 31864
rect 3700 31826 3752 31832
rect 3896 31822 3924 32558
rect 4172 32434 4200 32558
rect 4160 32428 4212 32434
rect 4160 32370 4212 32376
rect 4068 32360 4120 32366
rect 4068 32302 4120 32308
rect 3976 32224 4028 32230
rect 3976 32166 4028 32172
rect 3884 31816 3936 31822
rect 3884 31758 3936 31764
rect 3988 31521 4016 32166
rect 3974 31512 4030 31521
rect 3974 31447 4030 31456
rect 3976 31408 4028 31414
rect 3976 31350 4028 31356
rect 3884 31204 3936 31210
rect 3884 31146 3936 31152
rect 3700 31136 3752 31142
rect 3700 31078 3752 31084
rect 3712 30122 3740 31078
rect 3700 30116 3752 30122
rect 3700 30058 3752 30064
rect 3608 29776 3660 29782
rect 3608 29718 3660 29724
rect 3712 27402 3740 30058
rect 3896 28422 3924 31146
rect 3988 29850 4016 31350
rect 4080 31260 4108 32302
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4632 32026 4660 32778
rect 4620 32020 4672 32026
rect 4620 31962 4672 31968
rect 4620 31816 4672 31822
rect 4724 31804 4752 34954
rect 4804 33924 4856 33930
rect 4804 33866 4856 33872
rect 4816 33046 4844 33866
rect 4804 33040 4856 33046
rect 4804 32982 4856 32988
rect 4816 32858 4844 32982
rect 4908 32978 4936 36586
rect 5184 36378 5212 37606
rect 5538 37360 5594 37369
rect 5538 37295 5594 37304
rect 5172 36372 5224 36378
rect 5172 36314 5224 36320
rect 4988 36304 5040 36310
rect 4986 36272 4988 36281
rect 5040 36272 5042 36281
rect 4986 36207 5042 36216
rect 5080 36236 5132 36242
rect 5080 36178 5132 36184
rect 4988 35080 5040 35086
rect 4988 35022 5040 35028
rect 5000 34610 5028 35022
rect 4988 34604 5040 34610
rect 4988 34546 5040 34552
rect 4988 33652 5040 33658
rect 4988 33594 5040 33600
rect 4896 32972 4948 32978
rect 4896 32914 4948 32920
rect 4816 32842 4936 32858
rect 4816 32836 4948 32842
rect 4816 32830 4896 32836
rect 4896 32778 4948 32784
rect 4894 32464 4950 32473
rect 4894 32399 4896 32408
rect 4948 32399 4950 32408
rect 4896 32370 4948 32376
rect 4804 31952 4856 31958
rect 4804 31894 4856 31900
rect 4672 31776 4752 31804
rect 4620 31758 4672 31764
rect 4436 31680 4488 31686
rect 4436 31622 4488 31628
rect 4448 31414 4476 31622
rect 4436 31408 4488 31414
rect 4436 31350 4488 31356
rect 4160 31272 4212 31278
rect 4080 31232 4160 31260
rect 4080 30274 4108 31232
rect 4160 31214 4212 31220
rect 4448 31142 4476 31350
rect 4436 31136 4488 31142
rect 4436 31078 4488 31084
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4080 30258 4200 30274
rect 4080 30252 4212 30258
rect 4080 30246 4160 30252
rect 3976 29844 4028 29850
rect 3976 29786 4028 29792
rect 4080 29832 4108 30246
rect 4160 30194 4212 30200
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4160 29844 4212 29850
rect 4080 29804 4160 29832
rect 4080 28762 4108 29804
rect 4160 29786 4212 29792
rect 4632 29714 4660 31758
rect 4712 31476 4764 31482
rect 4712 31418 4764 31424
rect 4620 29708 4672 29714
rect 4620 29650 4672 29656
rect 4724 29646 4752 31418
rect 4816 30666 4844 31894
rect 4896 31884 4948 31890
rect 4896 31826 4948 31832
rect 4804 30660 4856 30666
rect 4804 30602 4856 30608
rect 4160 29640 4212 29646
rect 4160 29582 4212 29588
rect 4712 29640 4764 29646
rect 4712 29582 4764 29588
rect 4172 29510 4200 29582
rect 4160 29504 4212 29510
rect 4160 29446 4212 29452
rect 4804 28960 4856 28966
rect 4632 28920 4804 28948
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4068 28756 4120 28762
rect 4068 28698 4120 28704
rect 3884 28416 3936 28422
rect 3884 28358 3936 28364
rect 4080 28218 4108 28698
rect 4068 28212 4120 28218
rect 4068 28154 4120 28160
rect 4080 27674 4108 28154
rect 4632 27946 4660 28920
rect 4804 28902 4856 28908
rect 4620 27940 4672 27946
rect 4620 27882 4672 27888
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4068 27668 4120 27674
rect 4068 27610 4120 27616
rect 3700 27396 3752 27402
rect 3700 27338 3752 27344
rect 4080 27130 4108 27610
rect 4908 27538 4936 31826
rect 5000 29866 5028 33594
rect 5092 32314 5120 36178
rect 5184 36174 5212 36314
rect 5172 36168 5224 36174
rect 5172 36110 5224 36116
rect 5448 36168 5500 36174
rect 5448 36110 5500 36116
rect 5460 35086 5488 36110
rect 5448 35080 5500 35086
rect 5448 35022 5500 35028
rect 5172 34672 5224 34678
rect 5356 34672 5408 34678
rect 5224 34632 5356 34660
rect 5172 34614 5224 34620
rect 5552 34649 5580 37295
rect 5632 37256 5684 37262
rect 5632 37198 5684 37204
rect 5644 35136 5672 37198
rect 5828 36922 5856 39200
rect 6644 37120 6696 37126
rect 6644 37062 6696 37068
rect 5816 36916 5868 36922
rect 5816 36858 5868 36864
rect 6552 36780 6604 36786
rect 6552 36722 6604 36728
rect 6460 36712 6512 36718
rect 6460 36654 6512 36660
rect 5816 36576 5868 36582
rect 5816 36518 5868 36524
rect 6368 36576 6420 36582
rect 6368 36518 6420 36524
rect 5724 35692 5776 35698
rect 5724 35634 5776 35640
rect 5736 35494 5764 35634
rect 5724 35488 5776 35494
rect 5724 35430 5776 35436
rect 5644 35108 5764 35136
rect 5632 35012 5684 35018
rect 5632 34954 5684 34960
rect 5356 34614 5408 34620
rect 5538 34640 5594 34649
rect 5538 34575 5540 34584
rect 5592 34575 5594 34584
rect 5540 34546 5592 34552
rect 5356 34536 5408 34542
rect 5356 34478 5408 34484
rect 5264 32972 5316 32978
rect 5264 32914 5316 32920
rect 5276 32774 5304 32914
rect 5264 32768 5316 32774
rect 5264 32710 5316 32716
rect 5092 32286 5212 32314
rect 5080 31816 5132 31822
rect 5080 31758 5132 31764
rect 5092 31482 5120 31758
rect 5184 31482 5212 32286
rect 5276 31958 5304 32710
rect 5264 31952 5316 31958
rect 5264 31894 5316 31900
rect 5368 31754 5396 34478
rect 5540 34468 5592 34474
rect 5540 34410 5592 34416
rect 5448 33584 5500 33590
rect 5448 33526 5500 33532
rect 5460 33114 5488 33526
rect 5448 33108 5500 33114
rect 5448 33050 5500 33056
rect 5552 32910 5580 34410
rect 5448 32904 5500 32910
rect 5446 32872 5448 32881
rect 5540 32904 5592 32910
rect 5500 32872 5502 32881
rect 5540 32846 5592 32852
rect 5446 32807 5502 32816
rect 5446 32464 5502 32473
rect 5552 32434 5580 32846
rect 5446 32399 5502 32408
rect 5540 32428 5592 32434
rect 5460 31822 5488 32399
rect 5540 32370 5592 32376
rect 5448 31816 5500 31822
rect 5448 31758 5500 31764
rect 5276 31726 5396 31754
rect 5080 31476 5132 31482
rect 5080 31418 5132 31424
rect 5172 31476 5224 31482
rect 5172 31418 5224 31424
rect 5000 29838 5120 29866
rect 4988 28620 5040 28626
rect 4988 28562 5040 28568
rect 5000 28150 5028 28562
rect 4988 28144 5040 28150
rect 4988 28086 5040 28092
rect 5092 28082 5120 29838
rect 5276 29646 5304 31726
rect 5356 31476 5408 31482
rect 5356 31418 5408 31424
rect 5264 29640 5316 29646
rect 5264 29582 5316 29588
rect 5172 29028 5224 29034
rect 5172 28970 5224 28976
rect 5080 28076 5132 28082
rect 5080 28018 5132 28024
rect 5184 27878 5212 28970
rect 5276 28422 5304 29582
rect 5368 28966 5396 31418
rect 5448 31272 5500 31278
rect 5552 31260 5580 32370
rect 5500 31232 5580 31260
rect 5448 31214 5500 31220
rect 5448 31136 5500 31142
rect 5448 31078 5500 31084
rect 5356 28960 5408 28966
rect 5356 28902 5408 28908
rect 5264 28416 5316 28422
rect 5264 28358 5316 28364
rect 5172 27872 5224 27878
rect 5172 27814 5224 27820
rect 5184 27674 5212 27814
rect 5172 27668 5224 27674
rect 5172 27610 5224 27616
rect 4896 27532 4948 27538
rect 4896 27474 4948 27480
rect 3332 27124 3384 27130
rect 3332 27066 3384 27072
rect 4068 27124 4120 27130
rect 4068 27066 4120 27072
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 2596 26376 2648 26382
rect 2596 26318 2648 26324
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 1768 25152 1820 25158
rect 1768 25094 1820 25100
rect 2504 25152 2556 25158
rect 2504 25094 2556 25100
rect 2516 23730 2544 25094
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 1860 23724 1912 23730
rect 1860 23666 1912 23672
rect 2504 23724 2556 23730
rect 2504 23666 2556 23672
rect 1676 23520 1728 23526
rect 1676 23462 1728 23468
rect 1688 23225 1716 23462
rect 1674 23216 1730 23225
rect 1674 23151 1730 23160
rect 1872 22778 1900 23666
rect 2320 23520 2372 23526
rect 2320 23462 2372 23468
rect 1860 22772 1912 22778
rect 1860 22714 1912 22720
rect 2332 21554 2360 23462
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 3240 22432 3292 22438
rect 3240 22374 3292 22380
rect 2320 21548 2372 21554
rect 2320 21490 2372 21496
rect 1676 21344 1728 21350
rect 1676 21286 1728 21292
rect 1688 21185 1716 21286
rect 1674 21176 1730 21185
rect 1674 21111 1730 21120
rect 1674 19816 1730 19825
rect 1674 19751 1730 19760
rect 1688 19718 1716 19751
rect 1676 19712 1728 19718
rect 1676 19654 1728 19660
rect 1952 19712 2004 19718
rect 1952 19654 2004 19660
rect 1768 18624 1820 18630
rect 1768 18566 1820 18572
rect 1584 18284 1636 18290
rect 1584 18226 1636 18232
rect 1596 17814 1624 18226
rect 1584 17808 1636 17814
rect 1582 17776 1584 17785
rect 1636 17776 1638 17785
rect 1582 17711 1638 17720
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 1688 15745 1716 15846
rect 1674 15736 1730 15745
rect 1674 15671 1730 15680
rect 1674 14376 1730 14385
rect 1674 14311 1676 14320
rect 1728 14311 1730 14320
rect 1676 14282 1728 14288
rect 1688 14074 1716 14282
rect 1676 14068 1728 14074
rect 1676 14010 1728 14016
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 1688 12345 1716 12582
rect 1674 12336 1730 12345
rect 1674 12271 1730 12280
rect 1676 10464 1728 10470
rect 1676 10406 1728 10412
rect 1688 10305 1716 10406
rect 1674 10296 1730 10305
rect 1674 10231 1730 10240
rect 1584 8968 1636 8974
rect 1582 8936 1584 8945
rect 1636 8936 1638 8945
rect 1582 8871 1638 8880
rect 1596 8634 1624 8871
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 1676 7200 1728 7206
rect 1676 7142 1728 7148
rect 1688 6905 1716 7142
rect 1674 6896 1730 6905
rect 1674 6831 1730 6840
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1596 4865 1624 5170
rect 1582 4856 1638 4865
rect 1582 4791 1638 4800
rect 1674 3496 1730 3505
rect 1674 3431 1730 3440
rect 1688 3398 1716 3431
rect 1676 3392 1728 3398
rect 1676 3334 1728 3340
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 1308 2304 1360 2310
rect 1308 2246 1360 2252
rect 20 1352 72 1358
rect 20 1294 72 1300
rect 32 800 60 1294
rect 1320 800 1348 2246
rect 1688 1465 1716 2790
rect 1780 2446 1808 18566
rect 1860 13184 1912 13190
rect 1860 13126 1912 13132
rect 1872 12850 1900 13126
rect 1860 12844 1912 12850
rect 1860 12786 1912 12792
rect 1964 10674 1992 19654
rect 2502 18864 2558 18873
rect 2502 18799 2504 18808
rect 2556 18799 2558 18808
rect 2504 18770 2556 18776
rect 1952 10668 2004 10674
rect 1952 10610 2004 10616
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 1860 7404 1912 7410
rect 1860 7346 1912 7352
rect 1872 3738 1900 7346
rect 2792 5030 2820 9522
rect 2780 5024 2832 5030
rect 2780 4966 2832 4972
rect 1860 3732 1912 3738
rect 1860 3674 1912 3680
rect 2504 3528 2556 3534
rect 2504 3470 2556 3476
rect 2320 2848 2372 2854
rect 2320 2790 2372 2796
rect 2332 2446 2360 2790
rect 2516 2650 2544 3470
rect 3252 2650 3280 22374
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 5276 20058 5304 28358
rect 5460 27878 5488 31078
rect 5540 30660 5592 30666
rect 5644 30648 5672 34954
rect 5736 34746 5764 35108
rect 5724 34740 5776 34746
rect 5724 34682 5776 34688
rect 5828 34202 5856 36518
rect 5908 36100 5960 36106
rect 5908 36042 5960 36048
rect 6276 36100 6328 36106
rect 6276 36042 6328 36048
rect 5920 34474 5948 36042
rect 6184 35760 6236 35766
rect 6184 35702 6236 35708
rect 6196 34950 6224 35702
rect 6184 34944 6236 34950
rect 6184 34886 6236 34892
rect 5908 34468 5960 34474
rect 5908 34410 5960 34416
rect 5816 34196 5868 34202
rect 5816 34138 5868 34144
rect 5920 34066 5948 34410
rect 5908 34060 5960 34066
rect 5908 34002 5960 34008
rect 6184 34060 6236 34066
rect 6184 34002 6236 34008
rect 6196 33946 6224 34002
rect 6104 33918 6224 33946
rect 5908 33856 5960 33862
rect 5736 33804 5908 33810
rect 5736 33798 5960 33804
rect 5736 33782 5948 33798
rect 5736 31482 5764 33782
rect 6104 33454 6132 33918
rect 6092 33448 6144 33454
rect 6092 33390 6144 33396
rect 5908 32904 5960 32910
rect 5908 32846 5960 32852
rect 5816 31884 5868 31890
rect 5816 31826 5868 31832
rect 5724 31476 5776 31482
rect 5724 31418 5776 31424
rect 5724 31340 5776 31346
rect 5724 31282 5776 31288
rect 5592 30620 5672 30648
rect 5540 30602 5592 30608
rect 5540 30320 5592 30326
rect 5540 30262 5592 30268
rect 5552 28014 5580 30262
rect 5540 28008 5592 28014
rect 5540 27950 5592 27956
rect 5448 27872 5500 27878
rect 5448 27814 5500 27820
rect 5644 27334 5672 30620
rect 5736 27470 5764 31282
rect 5828 30734 5856 31826
rect 5920 31736 5948 32846
rect 6104 31890 6132 33390
rect 6288 33114 6316 36042
rect 6380 35630 6408 36518
rect 6368 35624 6420 35630
rect 6368 35566 6420 35572
rect 6380 33930 6408 35566
rect 6368 33924 6420 33930
rect 6368 33866 6420 33872
rect 6276 33108 6328 33114
rect 6276 33050 6328 33056
rect 6092 31884 6144 31890
rect 6092 31826 6144 31832
rect 6000 31748 6052 31754
rect 5920 31708 6000 31736
rect 6000 31690 6052 31696
rect 6012 31346 6040 31690
rect 6000 31340 6052 31346
rect 6000 31282 6052 31288
rect 5816 30728 5868 30734
rect 5816 30670 5868 30676
rect 5828 29850 5856 30670
rect 5908 30184 5960 30190
rect 5908 30126 5960 30132
rect 5920 29850 5948 30126
rect 5816 29844 5868 29850
rect 5816 29786 5868 29792
rect 5908 29844 5960 29850
rect 5908 29786 5960 29792
rect 5828 29306 5856 29786
rect 6276 29572 6328 29578
rect 6276 29514 6328 29520
rect 6288 29306 6316 29514
rect 5816 29300 5868 29306
rect 5816 29242 5868 29248
rect 6276 29300 6328 29306
rect 6276 29242 6328 29248
rect 5828 28762 5856 29242
rect 5816 28756 5868 28762
rect 5816 28698 5868 28704
rect 5828 28014 5856 28698
rect 5816 28008 5868 28014
rect 5816 27950 5868 27956
rect 5724 27464 5776 27470
rect 5724 27406 5776 27412
rect 5632 27328 5684 27334
rect 5632 27270 5684 27276
rect 5644 26790 5672 27270
rect 6276 27056 6328 27062
rect 6276 26998 6328 27004
rect 5632 26784 5684 26790
rect 5632 26726 5684 26732
rect 6288 26586 6316 26998
rect 6380 26586 6408 33866
rect 6472 31958 6500 36654
rect 6564 36009 6592 36722
rect 6550 36000 6606 36009
rect 6550 35935 6606 35944
rect 6552 35624 6604 35630
rect 6552 35566 6604 35572
rect 6564 35494 6592 35566
rect 6552 35488 6604 35494
rect 6552 35430 6604 35436
rect 6564 35154 6592 35430
rect 6656 35329 6684 37062
rect 7760 36922 7788 39200
rect 9312 37324 9364 37330
rect 9312 37266 9364 37272
rect 7840 37188 7892 37194
rect 7840 37130 7892 37136
rect 8576 37188 8628 37194
rect 8576 37130 8628 37136
rect 7748 36916 7800 36922
rect 7748 36858 7800 36864
rect 6828 36848 6880 36854
rect 6828 36790 6880 36796
rect 6736 35828 6788 35834
rect 6736 35770 6788 35776
rect 6642 35320 6698 35329
rect 6642 35255 6698 35264
rect 6552 35148 6604 35154
rect 6552 35090 6604 35096
rect 6564 34066 6592 35090
rect 6644 34468 6696 34474
rect 6644 34410 6696 34416
rect 6656 34134 6684 34410
rect 6644 34128 6696 34134
rect 6644 34070 6696 34076
rect 6748 34066 6776 35770
rect 6840 34746 6868 36790
rect 7656 36576 7708 36582
rect 7656 36518 7708 36524
rect 7668 36106 7696 36518
rect 7656 36100 7708 36106
rect 7656 36042 7708 36048
rect 7104 35760 7156 35766
rect 7104 35702 7156 35708
rect 7012 34944 7064 34950
rect 7012 34886 7064 34892
rect 6828 34740 6880 34746
rect 6828 34682 6880 34688
rect 6828 34604 6880 34610
rect 6828 34546 6880 34552
rect 6552 34060 6604 34066
rect 6552 34002 6604 34008
rect 6736 34060 6788 34066
rect 6736 34002 6788 34008
rect 6840 33522 6868 34546
rect 6552 33516 6604 33522
rect 6552 33458 6604 33464
rect 6828 33516 6880 33522
rect 6828 33458 6880 33464
rect 6564 32774 6592 33458
rect 6644 32836 6696 32842
rect 6644 32778 6696 32784
rect 6552 32768 6604 32774
rect 6552 32710 6604 32716
rect 6656 32570 6684 32778
rect 6828 32768 6880 32774
rect 6828 32710 6880 32716
rect 6644 32564 6696 32570
rect 6644 32506 6696 32512
rect 6460 31952 6512 31958
rect 6552 31952 6604 31958
rect 6460 31894 6512 31900
rect 6550 31920 6552 31929
rect 6604 31920 6606 31929
rect 6550 31855 6606 31864
rect 6552 31816 6604 31822
rect 6552 31758 6604 31764
rect 6460 30932 6512 30938
rect 6460 30874 6512 30880
rect 6472 29238 6500 30874
rect 6564 30258 6592 31758
rect 6840 31754 6868 32710
rect 7024 32570 7052 34886
rect 7116 33658 7144 35702
rect 7378 35320 7434 35329
rect 7288 35284 7340 35290
rect 7378 35255 7380 35264
rect 7288 35226 7340 35232
rect 7432 35255 7434 35264
rect 7380 35226 7432 35232
rect 7196 33992 7248 33998
rect 7196 33934 7248 33940
rect 7208 33862 7236 33934
rect 7196 33856 7248 33862
rect 7196 33798 7248 33804
rect 7104 33652 7156 33658
rect 7104 33594 7156 33600
rect 7208 33522 7236 33798
rect 7300 33658 7328 35226
rect 7472 35012 7524 35018
rect 7472 34954 7524 34960
rect 7380 33992 7432 33998
rect 7380 33934 7432 33940
rect 7288 33652 7340 33658
rect 7288 33594 7340 33600
rect 7196 33516 7248 33522
rect 7196 33458 7248 33464
rect 7012 32564 7064 32570
rect 7012 32506 7064 32512
rect 7208 32434 7236 33458
rect 7288 33448 7340 33454
rect 7392 33436 7420 33934
rect 7340 33408 7420 33436
rect 7288 33390 7340 33396
rect 7300 32434 7328 33390
rect 7484 32502 7512 34954
rect 7852 34202 7880 37130
rect 8300 37120 8352 37126
rect 8300 37062 8352 37068
rect 8312 36310 8340 37062
rect 8392 36712 8444 36718
rect 8392 36654 8444 36660
rect 8300 36304 8352 36310
rect 8300 36246 8352 36252
rect 8300 36168 8352 36174
rect 8300 36110 8352 36116
rect 8312 35154 8340 36110
rect 8300 35148 8352 35154
rect 8300 35090 8352 35096
rect 8404 34950 8432 36654
rect 8482 36272 8538 36281
rect 8482 36207 8538 36216
rect 8496 35018 8524 36207
rect 8484 35012 8536 35018
rect 8484 34954 8536 34960
rect 8392 34944 8444 34950
rect 8392 34886 8444 34892
rect 8484 34672 8536 34678
rect 8484 34614 8536 34620
rect 7840 34196 7892 34202
rect 7840 34138 7892 34144
rect 7932 33924 7984 33930
rect 7932 33866 7984 33872
rect 8208 33924 8260 33930
rect 8208 33866 8260 33872
rect 7840 33380 7892 33386
rect 7840 33322 7892 33328
rect 7746 32872 7802 32881
rect 7746 32807 7802 32816
rect 7760 32502 7788 32807
rect 7472 32496 7524 32502
rect 7472 32438 7524 32444
rect 7748 32496 7800 32502
rect 7748 32438 7800 32444
rect 7196 32428 7248 32434
rect 7196 32370 7248 32376
rect 7288 32428 7340 32434
rect 7340 32388 7420 32416
rect 7288 32370 7340 32376
rect 6748 31726 6868 31754
rect 7012 31748 7064 31754
rect 6644 30592 6696 30598
rect 6644 30534 6696 30540
rect 6552 30252 6604 30258
rect 6552 30194 6604 30200
rect 6552 29708 6604 29714
rect 6552 29650 6604 29656
rect 6460 29232 6512 29238
rect 6460 29174 6512 29180
rect 6564 29170 6592 29650
rect 6552 29164 6604 29170
rect 6552 29106 6604 29112
rect 6564 28626 6592 29106
rect 6552 28620 6604 28626
rect 6552 28562 6604 28568
rect 6656 27962 6684 30534
rect 6748 29578 6776 31726
rect 7012 31690 7064 31696
rect 7288 31748 7340 31754
rect 7288 31690 7340 31696
rect 6828 30184 6880 30190
rect 6828 30126 6880 30132
rect 6840 29714 6868 30126
rect 6828 29708 6880 29714
rect 6828 29650 6880 29656
rect 6736 29572 6788 29578
rect 6736 29514 6788 29520
rect 7024 28422 7052 31690
rect 7300 31482 7328 31690
rect 7288 31476 7340 31482
rect 7288 31418 7340 31424
rect 7392 31346 7420 32388
rect 7380 31340 7432 31346
rect 7380 31282 7432 31288
rect 7196 30728 7248 30734
rect 7196 30670 7248 30676
rect 7012 28416 7064 28422
rect 7012 28358 7064 28364
rect 6656 27934 6776 27962
rect 6644 27872 6696 27878
rect 6644 27814 6696 27820
rect 6276 26580 6328 26586
rect 6276 26522 6328 26528
rect 6368 26580 6420 26586
rect 6368 26522 6420 26528
rect 6092 26308 6144 26314
rect 6092 26250 6144 26256
rect 6104 23118 6132 26250
rect 6656 24070 6684 27814
rect 6748 26858 6776 27934
rect 7208 27606 7236 30670
rect 7380 30116 7432 30122
rect 7380 30058 7432 30064
rect 7392 29730 7420 30058
rect 7392 29702 7604 29730
rect 7576 29578 7604 29702
rect 7380 29572 7432 29578
rect 7380 29514 7432 29520
rect 7564 29572 7616 29578
rect 7564 29514 7616 29520
rect 7288 29232 7340 29238
rect 7392 29209 7420 29514
rect 7288 29174 7340 29180
rect 7378 29200 7434 29209
rect 7300 28762 7328 29174
rect 7378 29135 7434 29144
rect 7380 28960 7432 28966
rect 7380 28902 7432 28908
rect 7392 28762 7420 28902
rect 7288 28756 7340 28762
rect 7288 28698 7340 28704
rect 7380 28756 7432 28762
rect 7380 28698 7432 28704
rect 7852 28082 7880 33322
rect 7944 31482 7972 33866
rect 8220 33590 8248 33866
rect 8208 33584 8260 33590
rect 8208 33526 8260 33532
rect 8392 33584 8444 33590
rect 8392 33526 8444 33532
rect 8404 32026 8432 33526
rect 8496 32230 8524 34614
rect 8484 32224 8536 32230
rect 8484 32166 8536 32172
rect 8392 32020 8444 32026
rect 8392 31962 8444 31968
rect 7932 31476 7984 31482
rect 7932 31418 7984 31424
rect 8300 30796 8352 30802
rect 8300 30738 8352 30744
rect 8312 30394 8340 30738
rect 7932 30388 7984 30394
rect 7932 30330 7984 30336
rect 8300 30388 8352 30394
rect 8300 30330 8352 30336
rect 7944 30190 7972 30330
rect 8024 30320 8076 30326
rect 8024 30262 8076 30268
rect 8036 30190 8064 30262
rect 7932 30184 7984 30190
rect 7932 30126 7984 30132
rect 8024 30184 8076 30190
rect 8024 30126 8076 30132
rect 7944 29764 7972 30126
rect 8588 30054 8616 37130
rect 8668 37120 8720 37126
rect 8668 37062 8720 37068
rect 8680 36174 8708 37062
rect 9036 36576 9088 36582
rect 9036 36518 9088 36524
rect 9128 36576 9180 36582
rect 9128 36518 9180 36524
rect 8668 36168 8720 36174
rect 8668 36110 8720 36116
rect 9048 35766 9076 36518
rect 9140 36242 9168 36518
rect 9128 36236 9180 36242
rect 9128 36178 9180 36184
rect 9036 35760 9088 35766
rect 9036 35702 9088 35708
rect 8668 35624 8720 35630
rect 8668 35566 8720 35572
rect 8680 33862 8708 35566
rect 9140 35154 9168 36178
rect 9220 35624 9272 35630
rect 9220 35566 9272 35572
rect 8760 35148 8812 35154
rect 8760 35090 8812 35096
rect 9128 35148 9180 35154
rect 9128 35090 9180 35096
rect 8772 34134 8800 35090
rect 9036 35012 9088 35018
rect 9036 34954 9088 34960
rect 8760 34128 8812 34134
rect 8760 34070 8812 34076
rect 8668 33856 8720 33862
rect 8668 33798 8720 33804
rect 8680 32366 8708 33798
rect 8772 32978 8800 34070
rect 8852 33448 8904 33454
rect 8852 33390 8904 33396
rect 8760 32972 8812 32978
rect 8760 32914 8812 32920
rect 8668 32360 8720 32366
rect 8668 32302 8720 32308
rect 8576 30048 8628 30054
rect 8576 29990 8628 29996
rect 8116 29776 8168 29782
rect 7944 29736 8116 29764
rect 8116 29718 8168 29724
rect 8484 29504 8536 29510
rect 8484 29446 8536 29452
rect 8496 29102 8524 29446
rect 8484 29096 8536 29102
rect 8484 29038 8536 29044
rect 8300 29028 8352 29034
rect 8300 28970 8352 28976
rect 8312 28490 8340 28970
rect 8300 28484 8352 28490
rect 8300 28426 8352 28432
rect 8392 28484 8444 28490
rect 8392 28426 8444 28432
rect 7932 28416 7984 28422
rect 7932 28358 7984 28364
rect 7944 28082 7972 28358
rect 7840 28076 7892 28082
rect 7840 28018 7892 28024
rect 7932 28076 7984 28082
rect 7932 28018 7984 28024
rect 8404 27946 8432 28426
rect 8392 27940 8444 27946
rect 8392 27882 8444 27888
rect 7288 27872 7340 27878
rect 7288 27814 7340 27820
rect 8208 27872 8260 27878
rect 8208 27814 8260 27820
rect 7196 27600 7248 27606
rect 7196 27542 7248 27548
rect 6828 27532 6880 27538
rect 6828 27474 6880 27480
rect 6840 26926 6868 27474
rect 6828 26920 6880 26926
rect 6828 26862 6880 26868
rect 6736 26852 6788 26858
rect 6736 26794 6788 26800
rect 6840 26314 6868 26862
rect 6828 26308 6880 26314
rect 6828 26250 6880 26256
rect 6644 24064 6696 24070
rect 6644 24006 6696 24012
rect 6552 23724 6604 23730
rect 6552 23666 6604 23672
rect 6092 23112 6144 23118
rect 6092 23054 6144 23060
rect 6000 22976 6052 22982
rect 6000 22918 6052 22924
rect 5906 21992 5962 22001
rect 5906 21927 5962 21936
rect 5920 21894 5948 21927
rect 5908 21888 5960 21894
rect 5908 21830 5960 21836
rect 5264 20052 5316 20058
rect 5264 19994 5316 20000
rect 6012 19786 6040 22918
rect 6564 22438 6592 23666
rect 6552 22432 6604 22438
rect 6552 22374 6604 22380
rect 6276 21888 6328 21894
rect 6276 21830 6328 21836
rect 6000 19780 6052 19786
rect 6000 19722 6052 19728
rect 6184 19780 6236 19786
rect 6184 19722 6236 19728
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 6196 14346 6224 19722
rect 6184 14340 6236 14346
rect 6184 14282 6236 14288
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 6196 6914 6224 14282
rect 6288 9042 6316 21830
rect 7300 21622 7328 27814
rect 7656 27396 7708 27402
rect 7656 27338 7708 27344
rect 7668 26314 7696 27338
rect 7656 26308 7708 26314
rect 7656 26250 7708 26256
rect 7932 25220 7984 25226
rect 7932 25162 7984 25168
rect 7840 24132 7892 24138
rect 7840 24074 7892 24080
rect 7852 22574 7880 24074
rect 7944 23866 7972 25162
rect 7932 23860 7984 23866
rect 7932 23802 7984 23808
rect 8220 22710 8248 27814
rect 8576 27668 8628 27674
rect 8576 27610 8628 27616
rect 8588 26926 8616 27610
rect 8576 26920 8628 26926
rect 8576 26862 8628 26868
rect 8300 26580 8352 26586
rect 8300 26522 8352 26528
rect 8312 26042 8340 26522
rect 8300 26036 8352 26042
rect 8300 25978 8352 25984
rect 8680 24818 8708 32302
rect 8864 31754 8892 33390
rect 8944 32836 8996 32842
rect 8944 32778 8996 32784
rect 8956 32570 8984 32778
rect 8944 32564 8996 32570
rect 8944 32506 8996 32512
rect 8772 31726 8892 31754
rect 8772 27674 8800 31726
rect 8852 31408 8904 31414
rect 8852 31350 8904 31356
rect 8864 30802 8892 31350
rect 8852 30796 8904 30802
rect 8852 30738 8904 30744
rect 8852 29844 8904 29850
rect 8852 29786 8904 29792
rect 8864 29170 8892 29786
rect 8852 29164 8904 29170
rect 8852 29106 8904 29112
rect 8760 27668 8812 27674
rect 8760 27610 8812 27616
rect 9048 26994 9076 34954
rect 9232 33538 9260 35566
rect 9324 33658 9352 37266
rect 9692 36666 9720 39200
rect 10600 37324 10652 37330
rect 10600 37266 10652 37272
rect 10416 36712 10468 36718
rect 9692 36638 9812 36666
rect 10416 36654 10468 36660
rect 9680 36032 9732 36038
rect 9680 35974 9732 35980
rect 9692 35018 9720 35974
rect 9784 35698 9812 36638
rect 10428 36582 10456 36654
rect 10416 36576 10468 36582
rect 10416 36518 10468 36524
rect 9864 36100 9916 36106
rect 9864 36042 9916 36048
rect 9772 35692 9824 35698
rect 9772 35634 9824 35640
rect 9784 35290 9812 35634
rect 9772 35284 9824 35290
rect 9772 35226 9824 35232
rect 9680 35012 9732 35018
rect 9680 34954 9732 34960
rect 9876 34746 9904 36042
rect 10416 36032 10468 36038
rect 10416 35974 10468 35980
rect 10428 35698 10456 35974
rect 10416 35692 10468 35698
rect 10416 35634 10468 35640
rect 10508 35556 10560 35562
rect 10508 35498 10560 35504
rect 9956 35488 10008 35494
rect 9956 35430 10008 35436
rect 10416 35488 10468 35494
rect 10416 35430 10468 35436
rect 9968 35290 9996 35430
rect 9956 35284 10008 35290
rect 9956 35226 10008 35232
rect 9864 34740 9916 34746
rect 9864 34682 9916 34688
rect 9956 34740 10008 34746
rect 9956 34682 10008 34688
rect 9496 34672 9548 34678
rect 9416 34620 9496 34626
rect 9416 34614 9548 34620
rect 9586 34640 9642 34649
rect 9416 34598 9536 34614
rect 9416 34542 9444 34598
rect 9968 34626 9996 34682
rect 9586 34575 9642 34584
rect 9692 34598 9996 34626
rect 10140 34672 10192 34678
rect 10428 34649 10456 35430
rect 10520 35329 10548 35498
rect 10506 35320 10562 35329
rect 10506 35255 10562 35264
rect 10612 34678 10640 37266
rect 10876 37256 10928 37262
rect 10876 37198 10928 37204
rect 10784 36848 10836 36854
rect 10784 36790 10836 36796
rect 10796 36020 10824 36790
rect 10888 36718 10916 37198
rect 10980 37108 11008 39200
rect 12912 37262 12940 39200
rect 14844 37262 14872 39200
rect 16132 39114 16160 39200
rect 16224 39114 16252 39222
rect 16132 39086 16252 39114
rect 16592 37262 16620 39222
rect 18050 39200 18106 39800
rect 19982 39200 20038 39800
rect 21270 39200 21326 39800
rect 23202 39200 23258 39800
rect 23308 39222 23520 39250
rect 11704 37256 11756 37262
rect 11704 37198 11756 37204
rect 12900 37256 12952 37262
rect 12900 37198 12952 37204
rect 14832 37256 14884 37262
rect 14832 37198 14884 37204
rect 16580 37256 16632 37262
rect 16580 37198 16632 37204
rect 11060 37120 11112 37126
rect 10980 37080 11060 37108
rect 11060 37062 11112 37068
rect 11716 36922 11744 37198
rect 11796 37188 11848 37194
rect 11796 37130 11848 37136
rect 16120 37188 16172 37194
rect 16120 37130 16172 37136
rect 11808 36922 11836 37130
rect 13176 37120 13228 37126
rect 13176 37062 13228 37068
rect 13544 37120 13596 37126
rect 13544 37062 13596 37068
rect 15108 37120 15160 37126
rect 15108 37062 15160 37068
rect 15200 37120 15252 37126
rect 15200 37062 15252 37068
rect 11704 36916 11756 36922
rect 11704 36858 11756 36864
rect 11796 36916 11848 36922
rect 11796 36858 11848 36864
rect 11060 36780 11112 36786
rect 11060 36722 11112 36728
rect 13084 36780 13136 36786
rect 13084 36722 13136 36728
rect 10876 36712 10928 36718
rect 10876 36654 10928 36660
rect 10888 36378 10916 36654
rect 10876 36372 10928 36378
rect 10876 36314 10928 36320
rect 10968 36236 11020 36242
rect 10968 36178 11020 36184
rect 10876 36032 10928 36038
rect 10796 35992 10876 36020
rect 10876 35974 10928 35980
rect 10692 35148 10744 35154
rect 10692 35090 10744 35096
rect 10704 35057 10732 35090
rect 10690 35048 10746 35057
rect 10690 34983 10746 34992
rect 10784 34944 10836 34950
rect 10784 34886 10836 34892
rect 10600 34672 10652 34678
rect 10140 34614 10192 34620
rect 10414 34640 10470 34649
rect 9404 34536 9456 34542
rect 9404 34478 9456 34484
rect 9600 34490 9628 34575
rect 9692 34490 9720 34598
rect 9600 34462 9720 34490
rect 9772 34536 9824 34542
rect 9772 34478 9824 34484
rect 9588 34400 9640 34406
rect 9588 34342 9640 34348
rect 9600 34134 9628 34342
rect 9588 34128 9640 34134
rect 9588 34070 9640 34076
rect 9312 33652 9364 33658
rect 9312 33594 9364 33600
rect 9232 33510 9352 33538
rect 9128 32972 9180 32978
rect 9128 32914 9180 32920
rect 9140 32570 9168 32914
rect 9128 32564 9180 32570
rect 9128 32506 9180 32512
rect 9140 32026 9168 32506
rect 9128 32020 9180 32026
rect 9128 31962 9180 31968
rect 9140 31482 9168 31962
rect 9324 31754 9352 33510
rect 9600 33454 9628 34070
rect 9784 34066 9812 34478
rect 9772 34060 9824 34066
rect 9772 34002 9824 34008
rect 9588 33448 9640 33454
rect 9588 33390 9640 33396
rect 9496 32360 9548 32366
rect 9496 32302 9548 32308
rect 9324 31726 9444 31754
rect 9218 31512 9274 31521
rect 9128 31476 9180 31482
rect 9218 31447 9274 31456
rect 9128 31418 9180 31424
rect 9232 31414 9260 31447
rect 9220 31408 9272 31414
rect 9220 31350 9272 31356
rect 9128 31272 9180 31278
rect 9128 31214 9180 31220
rect 9140 29034 9168 31214
rect 9312 30660 9364 30666
rect 9312 30602 9364 30608
rect 9128 29028 9180 29034
rect 9128 28970 9180 28976
rect 9324 28218 9352 30602
rect 9312 28212 9364 28218
rect 9312 28154 9364 28160
rect 9312 27940 9364 27946
rect 9312 27882 9364 27888
rect 9324 27402 9352 27882
rect 9312 27396 9364 27402
rect 9312 27338 9364 27344
rect 9036 26988 9088 26994
rect 9036 26930 9088 26936
rect 9324 26586 9352 27338
rect 9312 26580 9364 26586
rect 9312 26522 9364 26528
rect 9312 25220 9364 25226
rect 9312 25162 9364 25168
rect 9324 24954 9352 25162
rect 9312 24948 9364 24954
rect 9312 24890 9364 24896
rect 8392 24812 8444 24818
rect 8392 24754 8444 24760
rect 8668 24812 8720 24818
rect 8668 24754 8720 24760
rect 8208 22704 8260 22710
rect 8208 22646 8260 22652
rect 7472 22568 7524 22574
rect 7472 22510 7524 22516
rect 7840 22568 7892 22574
rect 7840 22510 7892 22516
rect 8300 22568 8352 22574
rect 8300 22510 8352 22516
rect 7288 21616 7340 21622
rect 7288 21558 7340 21564
rect 7288 21480 7340 21486
rect 7484 21434 7512 22510
rect 8312 22166 8340 22510
rect 8404 22506 8432 24754
rect 8484 24132 8536 24138
rect 8484 24074 8536 24080
rect 8944 24132 8996 24138
rect 8944 24074 8996 24080
rect 8496 22778 8524 24074
rect 8484 22772 8536 22778
rect 8484 22714 8536 22720
rect 8956 22574 8984 24074
rect 9036 22704 9088 22710
rect 9036 22646 9088 22652
rect 8944 22568 8996 22574
rect 8944 22510 8996 22516
rect 8392 22500 8444 22506
rect 8392 22442 8444 22448
rect 8300 22160 8352 22166
rect 8300 22102 8352 22108
rect 7340 21428 7512 21434
rect 7288 21422 7512 21428
rect 8208 21480 8260 21486
rect 8208 21422 8260 21428
rect 7300 21406 7512 21422
rect 7300 13326 7328 21406
rect 7564 19712 7616 19718
rect 7564 19654 7616 19660
rect 7576 18698 7604 19654
rect 8220 18834 8248 21422
rect 8404 20058 8432 22442
rect 8956 22098 8984 22510
rect 9048 22234 9076 22646
rect 9036 22228 9088 22234
rect 9036 22170 9088 22176
rect 8944 22092 8996 22098
rect 8944 22034 8996 22040
rect 9416 22030 9444 31726
rect 9508 29850 9536 32302
rect 9784 31822 9812 34002
rect 9772 31816 9824 31822
rect 9772 31758 9824 31764
rect 9956 31816 10008 31822
rect 9956 31758 10008 31764
rect 9588 31680 9640 31686
rect 9588 31622 9640 31628
rect 9600 31482 9628 31622
rect 9588 31476 9640 31482
rect 9588 31418 9640 31424
rect 9784 30054 9812 31758
rect 9772 30048 9824 30054
rect 9772 29990 9824 29996
rect 9496 29844 9548 29850
rect 9496 29786 9548 29792
rect 9968 29238 9996 31758
rect 10048 31136 10100 31142
rect 10048 31078 10100 31084
rect 9680 29232 9732 29238
rect 9680 29174 9732 29180
rect 9956 29232 10008 29238
rect 9956 29174 10008 29180
rect 9496 28144 9548 28150
rect 9496 28086 9548 28092
rect 9508 27130 9536 28086
rect 9496 27124 9548 27130
rect 9496 27066 9548 27072
rect 9588 26852 9640 26858
rect 9588 26794 9640 26800
rect 9600 26518 9628 26794
rect 9588 26512 9640 26518
rect 9588 26454 9640 26460
rect 9496 26308 9548 26314
rect 9496 26250 9548 26256
rect 9508 24138 9536 26250
rect 9692 24682 9720 29174
rect 10060 29073 10088 31078
rect 10152 30258 10180 34614
rect 10600 34614 10652 34620
rect 10414 34575 10470 34584
rect 10796 33998 10824 34886
rect 10784 33992 10836 33998
rect 10784 33934 10836 33940
rect 10796 33590 10824 33934
rect 10416 33584 10468 33590
rect 10416 33526 10468 33532
rect 10784 33584 10836 33590
rect 10784 33526 10836 33532
rect 10232 32972 10284 32978
rect 10232 32914 10284 32920
rect 10244 32502 10272 32914
rect 10232 32496 10284 32502
rect 10232 32438 10284 32444
rect 10324 32428 10376 32434
rect 10324 32370 10376 32376
rect 10336 32298 10364 32370
rect 10324 32292 10376 32298
rect 10324 32234 10376 32240
rect 10428 32026 10456 33526
rect 10692 32836 10744 32842
rect 10692 32778 10744 32784
rect 10416 32020 10468 32026
rect 10416 31962 10468 31968
rect 10428 31142 10456 31962
rect 10704 31958 10732 32778
rect 10784 32428 10836 32434
rect 10784 32370 10836 32376
rect 10692 31952 10744 31958
rect 10692 31894 10744 31900
rect 10600 31884 10652 31890
rect 10600 31826 10652 31832
rect 10416 31136 10468 31142
rect 10416 31078 10468 31084
rect 10140 30252 10192 30258
rect 10140 30194 10192 30200
rect 10046 29064 10102 29073
rect 10046 28999 10102 29008
rect 9772 27396 9824 27402
rect 9772 27338 9824 27344
rect 9784 27130 9812 27338
rect 9772 27124 9824 27130
rect 9772 27066 9824 27072
rect 9772 25696 9824 25702
rect 9772 25638 9824 25644
rect 9784 25158 9812 25638
rect 10152 25294 10180 30194
rect 10322 29200 10378 29209
rect 10322 29135 10378 29144
rect 10336 29034 10364 29135
rect 10232 29028 10284 29034
rect 10232 28970 10284 28976
rect 10324 29028 10376 29034
rect 10324 28970 10376 28976
rect 10244 25906 10272 28970
rect 10428 28082 10456 31078
rect 10612 30666 10640 31826
rect 10796 30938 10824 32370
rect 10784 30932 10836 30938
rect 10784 30874 10836 30880
rect 10888 30818 10916 35974
rect 10980 34610 11008 36178
rect 11072 36106 11100 36722
rect 11980 36712 12032 36718
rect 11980 36654 12032 36660
rect 11992 36378 12020 36654
rect 11980 36372 12032 36378
rect 11980 36314 12032 36320
rect 12532 36304 12584 36310
rect 12532 36246 12584 36252
rect 12544 36174 12572 36246
rect 12532 36168 12584 36174
rect 12532 36110 12584 36116
rect 11060 36100 11112 36106
rect 11060 36042 11112 36048
rect 12440 36032 12492 36038
rect 12440 35974 12492 35980
rect 12452 35766 12480 35974
rect 12992 35828 13044 35834
rect 12992 35770 13044 35776
rect 12440 35760 12492 35766
rect 12440 35702 12492 35708
rect 12624 35692 12676 35698
rect 12624 35634 12676 35640
rect 11980 35624 12032 35630
rect 11980 35566 12032 35572
rect 11704 35148 11756 35154
rect 11704 35090 11756 35096
rect 11796 35148 11848 35154
rect 11796 35090 11848 35096
rect 11612 35012 11664 35018
rect 11612 34954 11664 34960
rect 10968 34604 11020 34610
rect 10968 34546 11020 34552
rect 11520 34400 11572 34406
rect 11520 34342 11572 34348
rect 11532 33930 11560 34342
rect 11428 33924 11480 33930
rect 11428 33866 11480 33872
rect 11520 33924 11572 33930
rect 11520 33866 11572 33872
rect 10968 33856 11020 33862
rect 10968 33798 11020 33804
rect 10980 33318 11008 33798
rect 10968 33312 11020 33318
rect 10968 33254 11020 33260
rect 10968 32904 11020 32910
rect 10968 32846 11020 32852
rect 10980 32298 11008 32846
rect 10968 32292 11020 32298
rect 10968 32234 11020 32240
rect 11336 31816 11388 31822
rect 11336 31758 11388 31764
rect 11060 31748 11112 31754
rect 11060 31690 11112 31696
rect 10968 31136 11020 31142
rect 10968 31078 11020 31084
rect 10704 30790 10916 30818
rect 10600 30660 10652 30666
rect 10600 30602 10652 30608
rect 10508 30048 10560 30054
rect 10508 29990 10560 29996
rect 10416 28076 10468 28082
rect 10416 28018 10468 28024
rect 10428 26382 10456 28018
rect 10520 27538 10548 29990
rect 10612 29850 10640 30602
rect 10600 29844 10652 29850
rect 10600 29786 10652 29792
rect 10508 27532 10560 27538
rect 10508 27474 10560 27480
rect 10508 27396 10560 27402
rect 10508 27338 10560 27344
rect 10520 27130 10548 27338
rect 10508 27124 10560 27130
rect 10508 27066 10560 27072
rect 10508 26988 10560 26994
rect 10508 26930 10560 26936
rect 10416 26376 10468 26382
rect 10416 26318 10468 26324
rect 10520 26042 10548 26930
rect 10600 26784 10652 26790
rect 10600 26726 10652 26732
rect 10508 26036 10560 26042
rect 10508 25978 10560 25984
rect 10232 25900 10284 25906
rect 10232 25842 10284 25848
rect 10520 25838 10548 25978
rect 10508 25832 10560 25838
rect 10508 25774 10560 25780
rect 10140 25288 10192 25294
rect 10140 25230 10192 25236
rect 9772 25152 9824 25158
rect 9772 25094 9824 25100
rect 10152 24886 10180 25230
rect 10612 24886 10640 26726
rect 10704 26382 10732 30790
rect 10784 29096 10836 29102
rect 10784 29038 10836 29044
rect 10796 28626 10824 29038
rect 10784 28620 10836 28626
rect 10784 28562 10836 28568
rect 10876 26852 10928 26858
rect 10876 26794 10928 26800
rect 10692 26376 10744 26382
rect 10692 26318 10744 26324
rect 10140 24880 10192 24886
rect 10140 24822 10192 24828
rect 10600 24880 10652 24886
rect 10600 24822 10652 24828
rect 10508 24744 10560 24750
rect 10508 24686 10560 24692
rect 9680 24676 9732 24682
rect 9680 24618 9732 24624
rect 9496 24132 9548 24138
rect 9496 24074 9548 24080
rect 10324 23724 10376 23730
rect 10324 23666 10376 23672
rect 10336 22098 10364 23666
rect 10520 22574 10548 24686
rect 10704 23730 10732 26318
rect 10888 25294 10916 26794
rect 10980 26042 11008 31078
rect 11072 30190 11100 31690
rect 11348 31414 11376 31758
rect 11336 31408 11388 31414
rect 11336 31350 11388 31356
rect 11440 31142 11468 33866
rect 11624 33658 11652 34954
rect 11612 33652 11664 33658
rect 11612 33594 11664 33600
rect 11716 31754 11744 35090
rect 11808 34678 11836 35090
rect 11796 34672 11848 34678
rect 11796 34614 11848 34620
rect 11808 34474 11836 34614
rect 11992 34542 12020 35566
rect 12636 35329 12664 35634
rect 12622 35320 12678 35329
rect 12622 35255 12678 35264
rect 12900 35148 12952 35154
rect 12900 35090 12952 35096
rect 12532 34944 12584 34950
rect 12532 34886 12584 34892
rect 11980 34536 12032 34542
rect 11980 34478 12032 34484
rect 11796 34468 11848 34474
rect 11796 34410 11848 34416
rect 11992 31754 12020 34478
rect 12348 34468 12400 34474
rect 12348 34410 12400 34416
rect 12360 33930 12388 34410
rect 12348 33924 12400 33930
rect 12348 33866 12400 33872
rect 12256 33584 12308 33590
rect 12256 33526 12308 33532
rect 12164 32768 12216 32774
rect 12164 32710 12216 32716
rect 11624 31726 11744 31754
rect 11808 31726 12020 31754
rect 11428 31136 11480 31142
rect 11428 31078 11480 31084
rect 11152 30796 11204 30802
rect 11152 30738 11204 30744
rect 11060 30184 11112 30190
rect 11060 30126 11112 30132
rect 11072 29578 11100 30126
rect 11164 29646 11192 30738
rect 11336 30660 11388 30666
rect 11336 30602 11388 30608
rect 11152 29640 11204 29646
rect 11152 29582 11204 29588
rect 11060 29572 11112 29578
rect 11060 29514 11112 29520
rect 11348 28529 11376 30602
rect 11520 29572 11572 29578
rect 11520 29514 11572 29520
rect 11532 29306 11560 29514
rect 11520 29300 11572 29306
rect 11520 29242 11572 29248
rect 11624 28626 11652 31726
rect 11704 29844 11756 29850
rect 11704 29786 11756 29792
rect 11716 29238 11744 29786
rect 11704 29232 11756 29238
rect 11704 29174 11756 29180
rect 11612 28620 11664 28626
rect 11612 28562 11664 28568
rect 11334 28520 11390 28529
rect 11060 28484 11112 28490
rect 11334 28455 11336 28464
rect 11060 28426 11112 28432
rect 11388 28455 11390 28464
rect 11336 28426 11388 28432
rect 11072 28218 11100 28426
rect 11428 28416 11480 28422
rect 11428 28358 11480 28364
rect 11060 28212 11112 28218
rect 11060 28154 11112 28160
rect 11244 28076 11296 28082
rect 11244 28018 11296 28024
rect 11256 27470 11284 28018
rect 11244 27464 11296 27470
rect 11244 27406 11296 27412
rect 11440 26450 11468 28358
rect 11428 26444 11480 26450
rect 11428 26386 11480 26392
rect 10968 26036 11020 26042
rect 10968 25978 11020 25984
rect 11060 25696 11112 25702
rect 11060 25638 11112 25644
rect 10876 25288 10928 25294
rect 10876 25230 10928 25236
rect 10888 23866 10916 25230
rect 10876 23860 10928 23866
rect 10876 23802 10928 23808
rect 10888 23730 10916 23802
rect 10692 23724 10744 23730
rect 10692 23666 10744 23672
rect 10876 23724 10928 23730
rect 10876 23666 10928 23672
rect 10600 22704 10652 22710
rect 10600 22646 10652 22652
rect 10508 22568 10560 22574
rect 10508 22510 10560 22516
rect 10612 22234 10640 22646
rect 10876 22568 10928 22574
rect 10876 22510 10928 22516
rect 10600 22228 10652 22234
rect 10600 22170 10652 22176
rect 10324 22092 10376 22098
rect 10324 22034 10376 22040
rect 9404 22024 9456 22030
rect 9404 21966 9456 21972
rect 8392 20052 8444 20058
rect 8392 19994 8444 20000
rect 8208 18828 8260 18834
rect 8208 18770 8260 18776
rect 7564 18692 7616 18698
rect 7564 18634 7616 18640
rect 7380 18624 7432 18630
rect 7380 18566 7432 18572
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 7392 9654 7420 18566
rect 7380 9648 7432 9654
rect 7380 9590 7432 9596
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 10888 8634 10916 22510
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 6196 6886 6408 6914
rect 6380 6798 6408 6886
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6552 6656 6604 6662
rect 6552 6598 6604 6604
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 3988 3058 4016 4966
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 3976 3052 4028 3058
rect 3976 2994 4028 3000
rect 4620 2848 4672 2854
rect 4620 2790 4672 2796
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 2504 2644 2556 2650
rect 2504 2586 2556 2592
rect 3240 2644 3292 2650
rect 3240 2586 3292 2592
rect 4632 2446 4660 2790
rect 6564 2446 6592 6598
rect 10980 2922 11008 8434
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 10232 2848 10284 2854
rect 10232 2790 10284 2796
rect 1768 2440 1820 2446
rect 1768 2382 1820 2388
rect 2320 2440 2372 2446
rect 2320 2382 2372 2388
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 6552 2440 6604 2446
rect 6552 2382 6604 2388
rect 1674 1456 1730 1465
rect 1674 1391 1730 1400
rect 2332 1358 2360 2382
rect 10244 2378 10272 2790
rect 10980 2514 11008 2858
rect 11072 2650 11100 25638
rect 11808 25430 11836 31726
rect 11888 31680 11940 31686
rect 11888 31622 11940 31628
rect 11900 30666 11928 31622
rect 11888 30660 11940 30666
rect 11888 30602 11940 30608
rect 12176 30258 12204 32710
rect 12164 30252 12216 30258
rect 12164 30194 12216 30200
rect 11980 30048 12032 30054
rect 11980 29990 12032 29996
rect 11886 29064 11942 29073
rect 11886 28999 11942 29008
rect 11900 28082 11928 28999
rect 11992 28490 12020 29990
rect 12164 29776 12216 29782
rect 12164 29718 12216 29724
rect 12176 29306 12204 29718
rect 12164 29300 12216 29306
rect 12164 29242 12216 29248
rect 11980 28484 12032 28490
rect 11980 28426 12032 28432
rect 11888 28076 11940 28082
rect 11888 28018 11940 28024
rect 12176 27470 12204 29242
rect 12268 28665 12296 33526
rect 12440 32768 12492 32774
rect 12440 32710 12492 32716
rect 12452 32502 12480 32710
rect 12440 32496 12492 32502
rect 12440 32438 12492 32444
rect 12348 31136 12400 31142
rect 12348 31078 12400 31084
rect 12360 29850 12388 31078
rect 12440 30048 12492 30054
rect 12440 29990 12492 29996
rect 12348 29844 12400 29850
rect 12348 29786 12400 29792
rect 12452 29238 12480 29990
rect 12544 29646 12572 34886
rect 12716 33108 12768 33114
rect 12716 33050 12768 33056
rect 12728 32570 12756 33050
rect 12716 32564 12768 32570
rect 12716 32506 12768 32512
rect 12808 32564 12860 32570
rect 12808 32506 12860 32512
rect 12716 31884 12768 31890
rect 12716 31826 12768 31832
rect 12624 31272 12676 31278
rect 12624 31214 12676 31220
rect 12532 29640 12584 29646
rect 12532 29582 12584 29588
rect 12440 29232 12492 29238
rect 12440 29174 12492 29180
rect 12532 28960 12584 28966
rect 12532 28902 12584 28908
rect 12254 28656 12310 28665
rect 12254 28591 12310 28600
rect 12348 28620 12400 28626
rect 12268 28218 12296 28591
rect 12348 28562 12400 28568
rect 12256 28212 12308 28218
rect 12256 28154 12308 28160
rect 12256 27872 12308 27878
rect 12256 27814 12308 27820
rect 12164 27464 12216 27470
rect 12164 27406 12216 27412
rect 12164 26852 12216 26858
rect 12164 26794 12216 26800
rect 12176 26450 12204 26794
rect 12164 26444 12216 26450
rect 12164 26386 12216 26392
rect 12176 25974 12204 26386
rect 12164 25968 12216 25974
rect 12164 25910 12216 25916
rect 12072 25764 12124 25770
rect 12072 25706 12124 25712
rect 11796 25424 11848 25430
rect 11796 25366 11848 25372
rect 11244 25220 11296 25226
rect 11244 25162 11296 25168
rect 11612 25220 11664 25226
rect 11612 25162 11664 25168
rect 11152 24268 11204 24274
rect 11152 24210 11204 24216
rect 11164 23050 11192 24210
rect 11256 24138 11284 25162
rect 11244 24132 11296 24138
rect 11244 24074 11296 24080
rect 11152 23044 11204 23050
rect 11152 22986 11204 22992
rect 11520 23044 11572 23050
rect 11520 22986 11572 22992
rect 11164 20058 11192 22986
rect 11532 22234 11560 22986
rect 11624 22710 11652 25162
rect 11704 24744 11756 24750
rect 11704 24686 11756 24692
rect 11716 23594 11744 24686
rect 11796 24404 11848 24410
rect 11796 24346 11848 24352
rect 11808 24274 11836 24346
rect 12084 24274 12112 25706
rect 12164 25220 12216 25226
rect 12164 25162 12216 25168
rect 12176 24614 12204 25162
rect 12164 24608 12216 24614
rect 12164 24550 12216 24556
rect 11796 24268 11848 24274
rect 11796 24210 11848 24216
rect 12072 24268 12124 24274
rect 12072 24210 12124 24216
rect 11796 24132 11848 24138
rect 11796 24074 11848 24080
rect 11808 23866 11836 24074
rect 11796 23860 11848 23866
rect 11796 23802 11848 23808
rect 12268 23798 12296 27814
rect 12360 24410 12388 28562
rect 12544 28490 12572 28902
rect 12532 28484 12584 28490
rect 12532 28426 12584 28432
rect 12440 28144 12492 28150
rect 12440 28086 12492 28092
rect 12452 27606 12480 28086
rect 12636 28014 12664 31214
rect 12728 29238 12756 31826
rect 12820 31414 12848 32506
rect 12808 31408 12860 31414
rect 12808 31350 12860 31356
rect 12808 31272 12860 31278
rect 12808 31214 12860 31220
rect 12820 30666 12848 31214
rect 12808 30660 12860 30666
rect 12808 30602 12860 30608
rect 12820 30394 12848 30602
rect 12808 30388 12860 30394
rect 12808 30330 12860 30336
rect 12820 29782 12848 30330
rect 12912 30054 12940 35090
rect 13004 34202 13032 35770
rect 13096 35034 13124 36722
rect 13188 35154 13216 37062
rect 13360 36848 13412 36854
rect 13360 36790 13412 36796
rect 13176 35148 13228 35154
rect 13176 35090 13228 35096
rect 13266 35048 13322 35057
rect 13096 35006 13216 35034
rect 13188 34542 13216 35006
rect 13266 34983 13322 34992
rect 13280 34610 13308 34983
rect 13268 34604 13320 34610
rect 13268 34546 13320 34552
rect 13176 34536 13228 34542
rect 13176 34478 13228 34484
rect 12992 34196 13044 34202
rect 12992 34138 13044 34144
rect 13188 32570 13216 34478
rect 13268 33856 13320 33862
rect 13268 33798 13320 33804
rect 13280 33522 13308 33798
rect 13268 33516 13320 33522
rect 13268 33458 13320 33464
rect 13176 32564 13228 32570
rect 13176 32506 13228 32512
rect 13280 32042 13308 33458
rect 13096 32014 13308 32042
rect 13096 30734 13124 32014
rect 13372 31822 13400 36790
rect 13556 36718 13584 37062
rect 13820 36916 13872 36922
rect 13820 36858 13872 36864
rect 13544 36712 13596 36718
rect 13544 36654 13596 36660
rect 13556 36038 13584 36654
rect 13832 36378 13860 36858
rect 15120 36786 15148 37062
rect 15212 36854 15240 37062
rect 15200 36848 15252 36854
rect 15200 36790 15252 36796
rect 14004 36780 14056 36786
rect 14004 36722 14056 36728
rect 15108 36780 15160 36786
rect 15108 36722 15160 36728
rect 13820 36372 13872 36378
rect 13820 36314 13872 36320
rect 13544 36032 13596 36038
rect 13544 35974 13596 35980
rect 13556 35834 13584 35974
rect 13544 35828 13596 35834
rect 13544 35770 13596 35776
rect 13556 35290 13584 35770
rect 13544 35284 13596 35290
rect 13544 35226 13596 35232
rect 14016 35222 14044 36722
rect 14372 36644 14424 36650
rect 14372 36586 14424 36592
rect 14384 36106 14412 36586
rect 14832 36372 14884 36378
rect 14832 36314 14884 36320
rect 14372 36100 14424 36106
rect 14372 36042 14424 36048
rect 14004 35216 14056 35222
rect 14004 35158 14056 35164
rect 13636 33856 13688 33862
rect 13636 33798 13688 33804
rect 13544 33312 13596 33318
rect 13544 33254 13596 33260
rect 13556 32842 13584 33254
rect 13648 32842 13676 33798
rect 14016 33522 14044 35158
rect 14384 34202 14412 36042
rect 14844 35290 14872 36314
rect 15120 36174 15148 36722
rect 16132 36718 16160 37130
rect 18064 37126 18092 39200
rect 18144 37256 18196 37262
rect 18144 37198 18196 37204
rect 18788 37256 18840 37262
rect 18788 37198 18840 37204
rect 18052 37120 18104 37126
rect 18052 37062 18104 37068
rect 18156 36922 18184 37198
rect 18144 36916 18196 36922
rect 18144 36858 18196 36864
rect 16120 36712 16172 36718
rect 16120 36654 16172 36660
rect 15108 36168 15160 36174
rect 15108 36110 15160 36116
rect 15936 36032 15988 36038
rect 15936 35974 15988 35980
rect 15948 35834 15976 35974
rect 15108 35828 15160 35834
rect 15108 35770 15160 35776
rect 15936 35828 15988 35834
rect 15936 35770 15988 35776
rect 14832 35284 14884 35290
rect 14832 35226 14884 35232
rect 14844 34746 14872 35226
rect 15120 34746 15148 35770
rect 15476 35692 15528 35698
rect 15476 35634 15528 35640
rect 14832 34740 14884 34746
rect 14832 34682 14884 34688
rect 15108 34740 15160 34746
rect 15108 34682 15160 34688
rect 15120 34202 15148 34682
rect 14372 34196 14424 34202
rect 14372 34138 14424 34144
rect 15108 34196 15160 34202
rect 15108 34138 15160 34144
rect 14384 33998 14412 34138
rect 14464 34128 14516 34134
rect 14464 34070 14516 34076
rect 14372 33992 14424 33998
rect 14372 33934 14424 33940
rect 14004 33516 14056 33522
rect 14004 33458 14056 33464
rect 14372 33312 14424 33318
rect 14372 33254 14424 33260
rect 13728 33040 13780 33046
rect 13728 32982 13780 32988
rect 13544 32836 13596 32842
rect 13544 32778 13596 32784
rect 13636 32836 13688 32842
rect 13636 32778 13688 32784
rect 13544 31884 13596 31890
rect 13544 31826 13596 31832
rect 13360 31816 13412 31822
rect 13360 31758 13412 31764
rect 13452 31748 13504 31754
rect 13452 31690 13504 31696
rect 13084 30728 13136 30734
rect 13084 30670 13136 30676
rect 13084 30592 13136 30598
rect 13084 30534 13136 30540
rect 12992 30184 13044 30190
rect 12992 30126 13044 30132
rect 12900 30048 12952 30054
rect 12900 29990 12952 29996
rect 12808 29776 12860 29782
rect 12808 29718 12860 29724
rect 12808 29640 12860 29646
rect 12808 29582 12860 29588
rect 12716 29232 12768 29238
rect 12716 29174 12768 29180
rect 12624 28008 12676 28014
rect 12624 27950 12676 27956
rect 12440 27600 12492 27606
rect 12440 27542 12492 27548
rect 12636 27538 12664 27950
rect 12624 27532 12676 27538
rect 12624 27474 12676 27480
rect 12624 27396 12676 27402
rect 12624 27338 12676 27344
rect 12716 27396 12768 27402
rect 12716 27338 12768 27344
rect 12440 27328 12492 27334
rect 12440 27270 12492 27276
rect 12452 26994 12480 27270
rect 12440 26988 12492 26994
rect 12440 26930 12492 26936
rect 12532 26580 12584 26586
rect 12532 26522 12584 26528
rect 12544 26246 12572 26522
rect 12532 26240 12584 26246
rect 12532 26182 12584 26188
rect 12636 25226 12664 27338
rect 12728 27062 12756 27338
rect 12716 27056 12768 27062
rect 12716 26998 12768 27004
rect 12728 26382 12756 26998
rect 12716 26376 12768 26382
rect 12716 26318 12768 26324
rect 12624 25220 12676 25226
rect 12624 25162 12676 25168
rect 12532 24948 12584 24954
rect 12532 24890 12584 24896
rect 12348 24404 12400 24410
rect 12348 24346 12400 24352
rect 12544 24274 12572 24890
rect 12820 24664 12848 29582
rect 13004 29578 13032 30126
rect 12992 29572 13044 29578
rect 12992 29514 13044 29520
rect 12900 29504 12952 29510
rect 12900 29446 12952 29452
rect 12912 27928 12940 29446
rect 12992 27940 13044 27946
rect 12912 27900 12992 27928
rect 12992 27882 13044 27888
rect 12900 26376 12952 26382
rect 12900 26318 12952 26324
rect 12636 24636 12848 24664
rect 12532 24268 12584 24274
rect 12532 24210 12584 24216
rect 12348 24200 12400 24206
rect 12348 24142 12400 24148
rect 12360 23866 12388 24142
rect 12348 23860 12400 23866
rect 12348 23802 12400 23808
rect 12256 23792 12308 23798
rect 12256 23734 12308 23740
rect 11980 23724 12032 23730
rect 11980 23666 12032 23672
rect 11704 23588 11756 23594
rect 11704 23530 11756 23536
rect 11716 23254 11744 23530
rect 11704 23248 11756 23254
rect 11704 23190 11756 23196
rect 11612 22704 11664 22710
rect 11612 22646 11664 22652
rect 11992 22642 12020 23666
rect 12636 23118 12664 24636
rect 12808 24064 12860 24070
rect 12808 24006 12860 24012
rect 12820 23662 12848 24006
rect 12808 23656 12860 23662
rect 12808 23598 12860 23604
rect 12348 23112 12400 23118
rect 12348 23054 12400 23060
rect 12624 23112 12676 23118
rect 12624 23054 12676 23060
rect 12360 22778 12388 23054
rect 12348 22772 12400 22778
rect 12348 22714 12400 22720
rect 11980 22636 12032 22642
rect 11980 22578 12032 22584
rect 12256 22636 12308 22642
rect 12256 22578 12308 22584
rect 11520 22228 11572 22234
rect 11520 22170 11572 22176
rect 11980 22024 12032 22030
rect 11980 21966 12032 21972
rect 11992 21622 12020 21966
rect 11980 21616 12032 21622
rect 11980 21558 12032 21564
rect 11992 21350 12020 21558
rect 11980 21344 12032 21350
rect 11980 21286 12032 21292
rect 11152 20052 11204 20058
rect 11152 19994 11204 20000
rect 11704 3460 11756 3466
rect 11704 3402 11756 3408
rect 11716 3194 11744 3402
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 11992 2582 12020 21286
rect 12268 21146 12296 22578
rect 12636 22438 12664 23054
rect 12820 22982 12848 23598
rect 12808 22976 12860 22982
rect 12808 22918 12860 22924
rect 12624 22432 12676 22438
rect 12624 22374 12676 22380
rect 12636 21690 12664 22374
rect 12716 22094 12768 22098
rect 12912 22094 12940 26318
rect 13004 26314 13032 27882
rect 13096 27402 13124 30534
rect 13176 30116 13228 30122
rect 13176 30058 13228 30064
rect 13188 29578 13216 30058
rect 13176 29572 13228 29578
rect 13176 29514 13228 29520
rect 13360 29028 13412 29034
rect 13360 28970 13412 28976
rect 13372 28762 13400 28970
rect 13360 28756 13412 28762
rect 13360 28698 13412 28704
rect 13464 28234 13492 31690
rect 13372 28206 13492 28234
rect 13084 27396 13136 27402
rect 13084 27338 13136 27344
rect 13084 27056 13136 27062
rect 13084 26998 13136 27004
rect 12992 26308 13044 26314
rect 12992 26250 13044 26256
rect 13004 24342 13032 26250
rect 13096 25498 13124 26998
rect 13268 26852 13320 26858
rect 13268 26794 13320 26800
rect 13280 26518 13308 26794
rect 13268 26512 13320 26518
rect 13268 26454 13320 26460
rect 13176 25832 13228 25838
rect 13176 25774 13228 25780
rect 13084 25492 13136 25498
rect 13084 25434 13136 25440
rect 13188 24750 13216 25774
rect 13176 24744 13228 24750
rect 13176 24686 13228 24692
rect 12992 24336 13044 24342
rect 12992 24278 13044 24284
rect 13188 23798 13216 24686
rect 13372 24614 13400 28206
rect 13556 28150 13584 31826
rect 13648 29714 13676 32778
rect 13740 32366 13768 32982
rect 13728 32360 13780 32366
rect 13728 32302 13780 32308
rect 13740 31754 13768 32302
rect 14004 32292 14056 32298
rect 14004 32234 14056 32240
rect 13740 31748 13872 31754
rect 13740 31726 13820 31748
rect 13820 31690 13872 31696
rect 13728 31680 13780 31686
rect 13728 31622 13780 31628
rect 13740 30598 13768 31622
rect 13728 30592 13780 30598
rect 13728 30534 13780 30540
rect 13912 30252 13964 30258
rect 13912 30194 13964 30200
rect 13728 30048 13780 30054
rect 13728 29990 13780 29996
rect 13636 29708 13688 29714
rect 13636 29650 13688 29656
rect 13636 29096 13688 29102
rect 13636 29038 13688 29044
rect 13648 28966 13676 29038
rect 13636 28960 13688 28966
rect 13636 28902 13688 28908
rect 13544 28144 13596 28150
rect 13544 28086 13596 28092
rect 13556 26874 13584 28086
rect 13464 26846 13584 26874
rect 13464 25362 13492 26846
rect 13544 26784 13596 26790
rect 13544 26726 13596 26732
rect 13556 26314 13584 26726
rect 13544 26308 13596 26314
rect 13544 26250 13596 26256
rect 13648 25770 13676 28902
rect 13740 27674 13768 29990
rect 13924 29306 13952 30194
rect 13912 29300 13964 29306
rect 13912 29242 13964 29248
rect 14016 29238 14044 32234
rect 14188 32224 14240 32230
rect 14188 32166 14240 32172
rect 14096 31816 14148 31822
rect 14096 31758 14148 31764
rect 14108 30258 14136 31758
rect 14200 31414 14228 32166
rect 14188 31408 14240 31414
rect 14188 31350 14240 31356
rect 14384 30802 14412 33254
rect 14372 30796 14424 30802
rect 14372 30738 14424 30744
rect 14188 30660 14240 30666
rect 14188 30602 14240 30608
rect 14096 30252 14148 30258
rect 14200 30240 14228 30602
rect 14280 30252 14332 30258
rect 14200 30212 14280 30240
rect 14096 30194 14148 30200
rect 14280 30194 14332 30200
rect 14384 30190 14412 30738
rect 14372 30184 14424 30190
rect 14372 30126 14424 30132
rect 14096 30048 14148 30054
rect 14096 29990 14148 29996
rect 14004 29232 14056 29238
rect 14004 29174 14056 29180
rect 13820 28756 13872 28762
rect 13820 28698 13872 28704
rect 13728 27668 13780 27674
rect 13728 27610 13780 27616
rect 13728 27532 13780 27538
rect 13728 27474 13780 27480
rect 13740 27062 13768 27474
rect 13728 27056 13780 27062
rect 13728 26998 13780 27004
rect 13832 26790 13860 28698
rect 14108 28422 14136 29990
rect 14280 29776 14332 29782
rect 14280 29718 14332 29724
rect 14096 28416 14148 28422
rect 14096 28358 14148 28364
rect 14292 28014 14320 29718
rect 14372 28416 14424 28422
rect 14372 28358 14424 28364
rect 14280 28008 14332 28014
rect 14280 27950 14332 27956
rect 14292 27130 14320 27950
rect 14280 27124 14332 27130
rect 14280 27066 14332 27072
rect 14384 27062 14412 28358
rect 14372 27056 14424 27062
rect 14372 26998 14424 27004
rect 14476 26874 14504 34070
rect 15120 33658 15148 34138
rect 15108 33652 15160 33658
rect 15108 33594 15160 33600
rect 14740 33108 14792 33114
rect 14740 33050 14792 33056
rect 14556 29300 14608 29306
rect 14556 29242 14608 29248
rect 14568 29102 14596 29242
rect 14556 29096 14608 29102
rect 14556 29038 14608 29044
rect 14646 28656 14702 28665
rect 14646 28591 14702 28600
rect 14660 28558 14688 28591
rect 14648 28552 14700 28558
rect 14648 28494 14700 28500
rect 14556 27328 14608 27334
rect 14556 27270 14608 27276
rect 14568 27130 14596 27270
rect 14556 27124 14608 27130
rect 14556 27066 14608 27072
rect 13924 26846 14504 26874
rect 13820 26784 13872 26790
rect 13820 26726 13872 26732
rect 13636 25764 13688 25770
rect 13636 25706 13688 25712
rect 13452 25356 13504 25362
rect 13452 25298 13504 25304
rect 13728 25220 13780 25226
rect 13728 25162 13780 25168
rect 13360 24608 13412 24614
rect 13360 24550 13412 24556
rect 13452 24268 13504 24274
rect 13452 24210 13504 24216
rect 13176 23792 13228 23798
rect 13176 23734 13228 23740
rect 12716 22092 12940 22094
rect 12768 22066 12940 22092
rect 12716 22034 12768 22040
rect 12624 21684 12676 21690
rect 12624 21626 12676 21632
rect 12992 21548 13044 21554
rect 12992 21490 13044 21496
rect 13004 21146 13032 21490
rect 12256 21140 12308 21146
rect 12256 21082 12308 21088
rect 12992 21140 13044 21146
rect 12992 21082 13044 21088
rect 13004 20806 13032 21082
rect 12992 20800 13044 20806
rect 12992 20742 13044 20748
rect 13004 18086 13032 20742
rect 12992 18080 13044 18086
rect 12992 18022 13044 18028
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 11980 2576 12032 2582
rect 11980 2518 12032 2524
rect 10968 2508 11020 2514
rect 10968 2450 11020 2456
rect 13096 2446 13124 14010
rect 13188 9382 13216 23734
rect 13464 13938 13492 24210
rect 13740 23662 13768 25162
rect 13820 23792 13872 23798
rect 13820 23734 13872 23740
rect 13728 23656 13780 23662
rect 13728 23598 13780 23604
rect 13544 22976 13596 22982
rect 13544 22918 13596 22924
rect 13556 22710 13584 22918
rect 13544 22704 13596 22710
rect 13544 22646 13596 22652
rect 13740 21690 13768 23598
rect 13832 23322 13860 23734
rect 13820 23316 13872 23322
rect 13820 23258 13872 23264
rect 13924 21962 13952 26846
rect 14004 26308 14056 26314
rect 14004 26250 14056 26256
rect 14016 25838 14044 26250
rect 14004 25832 14056 25838
rect 14004 25774 14056 25780
rect 14016 22098 14044 25774
rect 14660 25498 14688 28494
rect 14752 28121 14780 33050
rect 14832 32836 14884 32842
rect 14832 32778 14884 32784
rect 14844 28762 14872 32778
rect 15384 31816 15436 31822
rect 15384 31758 15436 31764
rect 15396 31414 15424 31758
rect 15384 31408 15436 31414
rect 15384 31350 15436 31356
rect 15200 31272 15252 31278
rect 15200 31214 15252 31220
rect 15212 30666 15240 31214
rect 15488 30734 15516 35634
rect 15568 35624 15620 35630
rect 15568 35566 15620 35572
rect 15580 35086 15608 35566
rect 15568 35080 15620 35086
rect 15568 35022 15620 35028
rect 15660 34944 15712 34950
rect 15660 34886 15712 34892
rect 16948 34944 17000 34950
rect 16948 34886 17000 34892
rect 15672 34678 15700 34886
rect 15660 34672 15712 34678
rect 15660 34614 15712 34620
rect 16960 34542 16988 34886
rect 16948 34536 17000 34542
rect 16948 34478 17000 34484
rect 15476 30728 15528 30734
rect 15476 30670 15528 30676
rect 15844 30728 15896 30734
rect 15844 30670 15896 30676
rect 15200 30660 15252 30666
rect 15200 30602 15252 30608
rect 15856 30598 15884 30670
rect 16212 30660 16264 30666
rect 16212 30602 16264 30608
rect 15568 30592 15620 30598
rect 15568 30534 15620 30540
rect 15844 30592 15896 30598
rect 15844 30534 15896 30540
rect 15108 30252 15160 30258
rect 15108 30194 15160 30200
rect 15120 30054 15148 30194
rect 15016 30048 15068 30054
rect 15016 29990 15068 29996
rect 15108 30048 15160 30054
rect 15108 29990 15160 29996
rect 14832 28756 14884 28762
rect 14832 28698 14884 28704
rect 14738 28112 14794 28121
rect 14738 28047 14794 28056
rect 14752 26994 14780 28047
rect 14844 27470 14872 28698
rect 15028 28694 15056 29990
rect 15580 29510 15608 30534
rect 15568 29504 15620 29510
rect 15568 29446 15620 29452
rect 15016 28688 15068 28694
rect 15016 28630 15068 28636
rect 15028 28014 15056 28630
rect 15292 28620 15344 28626
rect 15292 28562 15344 28568
rect 15304 28529 15332 28562
rect 15290 28520 15346 28529
rect 15290 28455 15346 28464
rect 15476 28484 15528 28490
rect 15016 28008 15068 28014
rect 15016 27950 15068 27956
rect 15304 27538 15332 28455
rect 15476 28426 15528 28432
rect 15568 28484 15620 28490
rect 15568 28426 15620 28432
rect 15488 28218 15516 28426
rect 15476 28212 15528 28218
rect 15476 28154 15528 28160
rect 15580 27946 15608 28426
rect 15752 28144 15804 28150
rect 15752 28086 15804 28092
rect 15568 27940 15620 27946
rect 15568 27882 15620 27888
rect 15764 27606 15792 28086
rect 15752 27600 15804 27606
rect 15752 27542 15804 27548
rect 15108 27532 15160 27538
rect 15108 27474 15160 27480
rect 15292 27532 15344 27538
rect 15292 27474 15344 27480
rect 15660 27532 15712 27538
rect 15660 27474 15712 27480
rect 14832 27464 14884 27470
rect 14832 27406 14884 27412
rect 14740 26988 14792 26994
rect 14740 26930 14792 26936
rect 14844 26382 14872 27406
rect 15016 26988 15068 26994
rect 15016 26930 15068 26936
rect 14832 26376 14884 26382
rect 14832 26318 14884 26324
rect 14924 25832 14976 25838
rect 14924 25774 14976 25780
rect 14648 25492 14700 25498
rect 14648 25434 14700 25440
rect 14372 25152 14424 25158
rect 14372 25094 14424 25100
rect 14384 24818 14412 25094
rect 14372 24812 14424 24818
rect 14372 24754 14424 24760
rect 14832 24608 14884 24614
rect 14832 24550 14884 24556
rect 14188 24132 14240 24138
rect 14188 24074 14240 24080
rect 14200 23662 14228 24074
rect 14188 23656 14240 23662
rect 14188 23598 14240 23604
rect 14188 23112 14240 23118
rect 14188 23054 14240 23060
rect 14004 22092 14056 22098
rect 14004 22034 14056 22040
rect 14096 22024 14148 22030
rect 14096 21966 14148 21972
rect 13912 21956 13964 21962
rect 13912 21898 13964 21904
rect 13924 21842 13952 21898
rect 14108 21894 14136 21966
rect 13832 21814 13952 21842
rect 14096 21888 14148 21894
rect 14096 21830 14148 21836
rect 13728 21684 13780 21690
rect 13728 21626 13780 21632
rect 13832 21554 13860 21814
rect 13820 21548 13872 21554
rect 13820 21490 13872 21496
rect 13832 21078 13860 21490
rect 13820 21072 13872 21078
rect 13820 21014 13872 21020
rect 13832 20466 13860 21014
rect 13820 20460 13872 20466
rect 13820 20402 13872 20408
rect 14108 16114 14136 21830
rect 14096 16108 14148 16114
rect 14096 16050 14148 16056
rect 13452 13932 13504 13938
rect 13452 13874 13504 13880
rect 13176 9376 13228 9382
rect 13176 9318 13228 9324
rect 14200 2582 14228 23054
rect 14740 22976 14792 22982
rect 14740 22918 14792 22924
rect 14752 22710 14780 22918
rect 14844 22710 14872 24550
rect 14936 24274 14964 25774
rect 15028 25294 15056 26930
rect 15016 25288 15068 25294
rect 15016 25230 15068 25236
rect 15120 24954 15148 27474
rect 15672 27402 15700 27474
rect 15660 27396 15712 27402
rect 15660 27338 15712 27344
rect 15200 27328 15252 27334
rect 15200 27270 15252 27276
rect 15212 26858 15240 27270
rect 15856 27130 15884 30534
rect 16028 30184 16080 30190
rect 16028 30126 16080 30132
rect 16040 28626 16068 30126
rect 16224 29714 16252 30602
rect 16212 29708 16264 29714
rect 16212 29650 16264 29656
rect 16224 29238 16252 29650
rect 16396 29572 16448 29578
rect 16396 29514 16448 29520
rect 16856 29572 16908 29578
rect 16856 29514 16908 29520
rect 16212 29232 16264 29238
rect 16212 29174 16264 29180
rect 16408 29102 16436 29514
rect 16396 29096 16448 29102
rect 16396 29038 16448 29044
rect 16304 29028 16356 29034
rect 16304 28970 16356 28976
rect 16028 28620 16080 28626
rect 16028 28562 16080 28568
rect 16316 28150 16344 28970
rect 16488 28620 16540 28626
rect 16488 28562 16540 28568
rect 16304 28144 16356 28150
rect 16304 28086 16356 28092
rect 16028 27872 16080 27878
rect 16028 27814 16080 27820
rect 16040 27402 16068 27814
rect 16316 27690 16344 28086
rect 16224 27662 16344 27690
rect 16028 27396 16080 27402
rect 16028 27338 16080 27344
rect 15844 27124 15896 27130
rect 15844 27066 15896 27072
rect 15200 26852 15252 26858
rect 15200 26794 15252 26800
rect 15212 25430 15240 26794
rect 15476 26784 15528 26790
rect 15476 26726 15528 26732
rect 15568 26784 15620 26790
rect 15568 26726 15620 26732
rect 15488 26518 15516 26726
rect 15476 26512 15528 26518
rect 15476 26454 15528 26460
rect 15580 26450 15608 26726
rect 15292 26444 15344 26450
rect 15292 26386 15344 26392
rect 15568 26444 15620 26450
rect 15568 26386 15620 26392
rect 15304 25974 15332 26386
rect 15384 26240 15436 26246
rect 15384 26182 15436 26188
rect 15292 25968 15344 25974
rect 15292 25910 15344 25916
rect 15200 25424 15252 25430
rect 15200 25366 15252 25372
rect 15108 24948 15160 24954
rect 15108 24890 15160 24896
rect 15396 24274 15424 26182
rect 15856 24750 15884 27066
rect 16120 27056 16172 27062
rect 16120 26998 16172 27004
rect 16132 26858 16160 26998
rect 16224 26926 16252 27662
rect 16304 27532 16356 27538
rect 16304 27474 16356 27480
rect 16316 27130 16344 27474
rect 16304 27124 16356 27130
rect 16304 27066 16356 27072
rect 16500 26994 16528 28562
rect 16868 28490 16896 29514
rect 17500 29504 17552 29510
rect 17500 29446 17552 29452
rect 17132 29300 17184 29306
rect 17132 29242 17184 29248
rect 16856 28484 16908 28490
rect 16856 28426 16908 28432
rect 17144 27062 17172 29242
rect 17512 29238 17540 29446
rect 18144 29300 18196 29306
rect 18144 29242 18196 29248
rect 17500 29232 17552 29238
rect 17500 29174 17552 29180
rect 18052 29164 18104 29170
rect 18052 29106 18104 29112
rect 18064 29073 18092 29106
rect 18050 29064 18106 29073
rect 18050 28999 18106 29008
rect 18052 28960 18104 28966
rect 18052 28902 18104 28908
rect 18064 28558 18092 28902
rect 18156 28762 18184 29242
rect 18144 28756 18196 28762
rect 18144 28698 18196 28704
rect 18052 28552 18104 28558
rect 18052 28494 18104 28500
rect 18064 28082 18092 28494
rect 18696 28416 18748 28422
rect 18696 28358 18748 28364
rect 18708 28121 18736 28358
rect 18694 28112 18750 28121
rect 18052 28076 18104 28082
rect 18694 28047 18696 28056
rect 18052 28018 18104 28024
rect 18748 28047 18750 28056
rect 18696 28018 18748 28024
rect 17316 28008 17368 28014
rect 17316 27950 17368 27956
rect 17224 27396 17276 27402
rect 17224 27338 17276 27344
rect 17132 27056 17184 27062
rect 17132 26998 17184 27004
rect 16488 26988 16540 26994
rect 16488 26930 16540 26936
rect 16212 26920 16264 26926
rect 16212 26862 16264 26868
rect 16120 26852 16172 26858
rect 16120 26794 16172 26800
rect 16856 26512 16908 26518
rect 16856 26454 16908 26460
rect 16868 26314 16896 26454
rect 16856 26308 16908 26314
rect 16856 26250 16908 26256
rect 16948 25696 17000 25702
rect 16948 25638 17000 25644
rect 16856 25220 16908 25226
rect 16856 25162 16908 25168
rect 16580 25152 16632 25158
rect 16580 25094 16632 25100
rect 16592 24886 16620 25094
rect 16580 24880 16632 24886
rect 16580 24822 16632 24828
rect 15844 24744 15896 24750
rect 15844 24686 15896 24692
rect 16488 24744 16540 24750
rect 16488 24686 16540 24692
rect 15752 24676 15804 24682
rect 15752 24618 15804 24624
rect 15764 24410 15792 24618
rect 15752 24404 15804 24410
rect 15752 24346 15804 24352
rect 15856 24274 15884 24686
rect 16028 24608 16080 24614
rect 16028 24550 16080 24556
rect 14924 24268 14976 24274
rect 14924 24210 14976 24216
rect 15384 24268 15436 24274
rect 15844 24268 15896 24274
rect 15436 24228 15516 24256
rect 15384 24210 15436 24216
rect 15384 24064 15436 24070
rect 15384 24006 15436 24012
rect 15396 23798 15424 24006
rect 15384 23792 15436 23798
rect 15384 23734 15436 23740
rect 15488 23662 15516 24228
rect 15844 24210 15896 24216
rect 16040 24138 16068 24550
rect 16028 24132 16080 24138
rect 16028 24074 16080 24080
rect 16120 24132 16172 24138
rect 16120 24074 16172 24080
rect 16132 23866 16160 24074
rect 16120 23860 16172 23866
rect 16120 23802 16172 23808
rect 15384 23656 15436 23662
rect 15384 23598 15436 23604
rect 15476 23656 15528 23662
rect 15476 23598 15528 23604
rect 15200 23248 15252 23254
rect 15200 23190 15252 23196
rect 14740 22704 14792 22710
rect 14740 22646 14792 22652
rect 14832 22704 14884 22710
rect 14832 22646 14884 22652
rect 15016 22500 15068 22506
rect 15016 22442 15068 22448
rect 14740 21480 14792 21486
rect 14740 21422 14792 21428
rect 14752 21010 14780 21422
rect 14740 21004 14792 21010
rect 14740 20946 14792 20952
rect 14832 20868 14884 20874
rect 14832 20810 14884 20816
rect 14844 20602 14872 20810
rect 14832 20596 14884 20602
rect 14832 20538 14884 20544
rect 15028 6458 15056 22442
rect 15212 22166 15240 23190
rect 15200 22160 15252 22166
rect 15200 22102 15252 22108
rect 15212 21418 15240 22102
rect 15292 22092 15344 22098
rect 15292 22034 15344 22040
rect 15304 21962 15332 22034
rect 15292 21956 15344 21962
rect 15292 21898 15344 21904
rect 15200 21412 15252 21418
rect 15200 21354 15252 21360
rect 15396 8634 15424 23598
rect 15488 22710 15516 23598
rect 16500 23186 16528 24686
rect 16868 24410 16896 25162
rect 16856 24404 16908 24410
rect 16856 24346 16908 24352
rect 16960 24206 16988 25638
rect 16948 24200 17000 24206
rect 16948 24142 17000 24148
rect 16488 23180 16540 23186
rect 16488 23122 16540 23128
rect 16500 23050 16528 23122
rect 15660 23044 15712 23050
rect 15660 22986 15712 22992
rect 16488 23044 16540 23050
rect 16488 22986 16540 22992
rect 15672 22778 15700 22986
rect 15660 22772 15712 22778
rect 15660 22714 15712 22720
rect 15476 22704 15528 22710
rect 15476 22646 15528 22652
rect 16212 22024 16264 22030
rect 16212 21966 16264 21972
rect 15752 21480 15804 21486
rect 15752 21422 15804 21428
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 15016 6452 15068 6458
rect 15016 6394 15068 6400
rect 14924 3392 14976 3398
rect 14924 3334 14976 3340
rect 14464 3120 14516 3126
rect 14464 3062 14516 3068
rect 14476 2922 14504 3062
rect 14936 2990 14964 3334
rect 15120 3194 15148 8434
rect 15764 8090 15792 21422
rect 16224 20602 16252 21966
rect 16396 20868 16448 20874
rect 16396 20810 16448 20816
rect 16212 20596 16264 20602
rect 16212 20538 16264 20544
rect 16408 18834 16436 20810
rect 16948 20324 17000 20330
rect 16948 20266 17000 20272
rect 16396 18828 16448 18834
rect 16396 18770 16448 18776
rect 16960 18698 16988 20266
rect 16948 18692 17000 18698
rect 16948 18634 17000 18640
rect 15752 8084 15804 8090
rect 15752 8026 15804 8032
rect 15844 7880 15896 7886
rect 15844 7822 15896 7828
rect 15568 6316 15620 6322
rect 15568 6258 15620 6264
rect 15580 3738 15608 6258
rect 15568 3732 15620 3738
rect 15568 3674 15620 3680
rect 15580 3534 15608 3674
rect 15568 3528 15620 3534
rect 15568 3470 15620 3476
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 14924 2984 14976 2990
rect 14924 2926 14976 2932
rect 14464 2916 14516 2922
rect 14464 2858 14516 2864
rect 14188 2576 14240 2582
rect 14188 2518 14240 2524
rect 13084 2440 13136 2446
rect 13084 2382 13136 2388
rect 15120 2378 15148 3130
rect 15856 3058 15884 7822
rect 17144 3126 17172 26998
rect 17236 26042 17264 27338
rect 17328 26450 17356 27950
rect 18064 27606 18092 28018
rect 18604 27940 18656 27946
rect 18604 27882 18656 27888
rect 18616 27674 18644 27882
rect 18604 27668 18656 27674
rect 18604 27610 18656 27616
rect 18052 27600 18104 27606
rect 18052 27542 18104 27548
rect 18604 27464 18656 27470
rect 18604 27406 18656 27412
rect 18420 27056 18472 27062
rect 18420 26998 18472 27004
rect 17500 26920 17552 26926
rect 17500 26862 17552 26868
rect 17512 26450 17540 26862
rect 17868 26852 17920 26858
rect 17868 26794 17920 26800
rect 17316 26444 17368 26450
rect 17316 26386 17368 26392
rect 17500 26444 17552 26450
rect 17500 26386 17552 26392
rect 17880 26042 17908 26794
rect 18236 26512 18288 26518
rect 18236 26454 18288 26460
rect 17960 26308 18012 26314
rect 17960 26250 18012 26256
rect 17224 26036 17276 26042
rect 17224 25978 17276 25984
rect 17868 26036 17920 26042
rect 17868 25978 17920 25984
rect 17972 25906 18000 26250
rect 17960 25900 18012 25906
rect 17960 25842 18012 25848
rect 18248 25498 18276 26454
rect 18432 26314 18460 26998
rect 18616 26994 18644 27406
rect 18800 27130 18828 37198
rect 19996 37126 20024 39200
rect 21284 37126 21312 39200
rect 23216 39114 23244 39200
rect 23308 39114 23336 39222
rect 23216 39086 23336 39114
rect 23492 37262 23520 39222
rect 25134 39200 25190 39800
rect 26422 39200 26478 39800
rect 28354 39200 28410 39800
rect 30286 39200 30342 39800
rect 31574 39200 31630 39800
rect 33506 39200 33562 39800
rect 35438 39200 35494 39800
rect 36726 39200 36782 39800
rect 25148 37466 25176 39200
rect 25136 37460 25188 37466
rect 25136 37402 25188 37408
rect 25148 37262 25176 37402
rect 22008 37256 22060 37262
rect 22008 37198 22060 37204
rect 23480 37256 23532 37262
rect 23480 37198 23532 37204
rect 25136 37256 25188 37262
rect 25136 37198 25188 37204
rect 21824 37188 21876 37194
rect 21824 37130 21876 37136
rect 19984 37120 20036 37126
rect 19984 37062 20036 37068
rect 21272 37120 21324 37126
rect 21272 37062 21324 37068
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19432 31816 19484 31822
rect 19432 31758 19484 31764
rect 19444 31414 19472 31758
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19432 31408 19484 31414
rect 19432 31350 19484 31356
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19340 30388 19392 30394
rect 19340 30330 19392 30336
rect 19248 27872 19300 27878
rect 19248 27814 19300 27820
rect 19156 27532 19208 27538
rect 19156 27474 19208 27480
rect 19168 27334 19196 27474
rect 19156 27328 19208 27334
rect 19156 27270 19208 27276
rect 18788 27124 18840 27130
rect 18788 27066 18840 27072
rect 19260 26994 19288 27814
rect 18604 26988 18656 26994
rect 18604 26930 18656 26936
rect 19248 26988 19300 26994
rect 19248 26930 19300 26936
rect 19260 26790 19288 26930
rect 19248 26784 19300 26790
rect 19248 26726 19300 26732
rect 19260 26382 19288 26726
rect 19248 26376 19300 26382
rect 19248 26318 19300 26324
rect 18420 26308 18472 26314
rect 18420 26250 18472 26256
rect 18236 25492 18288 25498
rect 18236 25434 18288 25440
rect 17868 25356 17920 25362
rect 17868 25298 17920 25304
rect 17500 25220 17552 25226
rect 17500 25162 17552 25168
rect 17512 24750 17540 25162
rect 17880 24818 17908 25298
rect 18328 25288 18380 25294
rect 18328 25230 18380 25236
rect 17868 24812 17920 24818
rect 17868 24754 17920 24760
rect 17500 24744 17552 24750
rect 17500 24686 17552 24692
rect 17868 24608 17920 24614
rect 17868 24550 17920 24556
rect 17880 24410 17908 24550
rect 17868 24404 17920 24410
rect 17868 24346 17920 24352
rect 17500 24200 17552 24206
rect 17500 24142 17552 24148
rect 17512 23866 17540 24142
rect 17500 23860 17552 23866
rect 17500 23802 17552 23808
rect 18340 22642 18368 25230
rect 18328 22636 18380 22642
rect 18328 22578 18380 22584
rect 17684 18624 17736 18630
rect 17684 18566 17736 18572
rect 17696 14346 17724 18566
rect 17684 14340 17736 14346
rect 17684 14282 17736 14288
rect 17132 3120 17184 3126
rect 17132 3062 17184 3068
rect 19352 3058 19380 30330
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19984 26240 20036 26246
rect 19984 26182 20036 26188
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19996 25906 20024 26182
rect 19984 25900 20036 25906
rect 19984 25842 20036 25848
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 21836 20058 21864 37130
rect 22020 36582 22048 37198
rect 26436 37126 26464 39200
rect 28368 37126 28396 39200
rect 30300 37330 30328 39200
rect 31588 37346 31616 39200
rect 30288 37324 30340 37330
rect 31588 37318 31708 37346
rect 30288 37266 30340 37272
rect 28448 37256 28500 37262
rect 28448 37198 28500 37204
rect 31484 37256 31536 37262
rect 31484 37198 31536 37204
rect 31680 37210 31708 37318
rect 25320 37120 25372 37126
rect 25320 37062 25372 37068
rect 26424 37120 26476 37126
rect 26424 37062 26476 37068
rect 28356 37120 28408 37126
rect 28356 37062 28408 37068
rect 22008 36576 22060 36582
rect 22008 36518 22060 36524
rect 24860 27328 24912 27334
rect 24860 27270 24912 27276
rect 22192 24676 22244 24682
rect 22192 24618 22244 24624
rect 22204 23730 22232 24618
rect 24492 24608 24544 24614
rect 24492 24550 24544 24556
rect 22192 23724 22244 23730
rect 22192 23666 22244 23672
rect 22204 23118 22232 23666
rect 22192 23112 22244 23118
rect 22192 23054 22244 23060
rect 21824 20052 21876 20058
rect 21824 19994 21876 20000
rect 21836 19854 21864 19994
rect 21824 19848 21876 19854
rect 21824 19790 21876 19796
rect 20812 19712 20864 19718
rect 20812 19654 20864 19660
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 15844 3052 15896 3058
rect 15844 2994 15896 3000
rect 19340 3052 19392 3058
rect 19340 2994 19392 3000
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 15212 2446 15240 2790
rect 15856 2650 15884 2994
rect 20824 2650 20852 19654
rect 22008 2848 22060 2854
rect 22008 2790 22060 2796
rect 15844 2644 15896 2650
rect 15844 2586 15896 2592
rect 20812 2644 20864 2650
rect 20812 2586 20864 2592
rect 20824 2446 20852 2586
rect 22020 2582 22048 2790
rect 22204 2650 22232 23054
rect 24504 8634 24532 24550
rect 24872 14414 24900 27270
rect 25332 24274 25360 37062
rect 28460 35290 28488 37198
rect 30564 37120 30616 37126
rect 30564 37062 30616 37068
rect 30576 36310 30604 37062
rect 30564 36304 30616 36310
rect 30564 36246 30616 36252
rect 28448 35284 28500 35290
rect 28448 35226 28500 35232
rect 27896 35080 27948 35086
rect 27896 35022 27948 35028
rect 27908 31822 27936 35022
rect 31496 33658 31524 37198
rect 31680 37182 31800 37210
rect 31772 37126 31800 37182
rect 31852 37188 31904 37194
rect 31852 37130 31904 37136
rect 31760 37120 31812 37126
rect 31760 37062 31812 37068
rect 31484 33652 31536 33658
rect 31484 33594 31536 33600
rect 27896 31816 27948 31822
rect 27896 31758 27948 31764
rect 25872 30048 25924 30054
rect 25872 29990 25924 29996
rect 25884 24818 25912 29990
rect 26148 27056 26200 27062
rect 26148 26998 26200 27004
rect 25872 24812 25924 24818
rect 25872 24754 25924 24760
rect 26160 24410 26188 26998
rect 31864 26234 31892 37130
rect 33520 37126 33548 39200
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 35452 37466 35480 39200
rect 35806 38856 35862 38865
rect 35806 38791 35862 38800
rect 35622 37496 35678 37505
rect 35440 37460 35492 37466
rect 35622 37431 35678 37440
rect 35440 37402 35492 37408
rect 35452 37262 35480 37402
rect 33600 37256 33652 37262
rect 33600 37198 33652 37204
rect 35440 37256 35492 37262
rect 35440 37198 35492 37204
rect 33508 37120 33560 37126
rect 33508 37062 33560 37068
rect 32404 26376 32456 26382
rect 32404 26318 32456 26324
rect 31772 26206 31892 26234
rect 26148 24404 26200 24410
rect 26148 24346 26200 24352
rect 25320 24268 25372 24274
rect 25320 24210 25372 24216
rect 30564 21956 30616 21962
rect 30564 21898 30616 21904
rect 27160 21684 27212 21690
rect 27160 21626 27212 21632
rect 25412 21140 25464 21146
rect 25412 21082 25464 21088
rect 25424 16114 25452 21082
rect 27172 17202 27200 21626
rect 30576 21146 30604 21898
rect 31772 21894 31800 26206
rect 31760 21888 31812 21894
rect 31760 21830 31812 21836
rect 30564 21140 30616 21146
rect 30564 21082 30616 21088
rect 27160 17196 27212 17202
rect 27160 17138 27212 17144
rect 25412 16108 25464 16114
rect 25412 16050 25464 16056
rect 25596 15904 25648 15910
rect 25596 15846 25648 15852
rect 25608 15706 25636 15846
rect 25596 15700 25648 15706
rect 25596 15642 25648 15648
rect 24860 14408 24912 14414
rect 24860 14350 24912 14356
rect 25044 14272 25096 14278
rect 25044 14214 25096 14220
rect 24492 8628 24544 8634
rect 24492 8570 24544 8576
rect 24676 2984 24728 2990
rect 24676 2926 24728 2932
rect 22192 2644 22244 2650
rect 22192 2586 22244 2592
rect 22008 2576 22060 2582
rect 22008 2518 22060 2524
rect 15200 2440 15252 2446
rect 15200 2382 15252 2388
rect 20812 2440 20864 2446
rect 20812 2382 20864 2388
rect 24688 2378 24716 2926
rect 25056 2650 25084 14214
rect 30012 8492 30064 8498
rect 30012 8434 30064 8440
rect 30024 3058 30052 8434
rect 30012 3052 30064 3058
rect 30012 2994 30064 3000
rect 25044 2644 25096 2650
rect 25044 2586 25096 2592
rect 30024 2514 30052 2994
rect 32220 2848 32272 2854
rect 32220 2790 32272 2796
rect 30012 2508 30064 2514
rect 30012 2450 30064 2456
rect 32232 2378 32260 2790
rect 32416 2650 32444 26318
rect 33416 24812 33468 24818
rect 33416 24754 33468 24760
rect 33428 24206 33456 24754
rect 33612 24682 33640 37198
rect 35532 37188 35584 37194
rect 35532 37130 35584 37136
rect 35544 36650 35572 37130
rect 35636 36922 35664 37431
rect 35820 36922 35848 38791
rect 35624 36916 35676 36922
rect 35624 36858 35676 36864
rect 35808 36916 35860 36922
rect 35808 36858 35860 36864
rect 35624 36780 35676 36786
rect 35624 36722 35676 36728
rect 36176 36780 36228 36786
rect 36176 36722 36228 36728
rect 35532 36644 35584 36650
rect 35532 36586 35584 36592
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35348 36032 35400 36038
rect 35348 35974 35400 35980
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34796 34400 34848 34406
rect 34796 34342 34848 34348
rect 34808 33998 34836 34342
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34796 33992 34848 33998
rect 34796 33934 34848 33940
rect 34980 33856 35032 33862
rect 34980 33798 35032 33804
rect 34992 33522 35020 33798
rect 34980 33516 35032 33522
rect 34980 33458 35032 33464
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 33600 24676 33652 24682
rect 33600 24618 33652 24624
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 33416 24200 33468 24206
rect 33416 24142 33468 24148
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 35360 22982 35388 35974
rect 35440 35488 35492 35494
rect 35440 35430 35492 35436
rect 35452 23526 35480 35430
rect 35636 32026 35664 36722
rect 35900 35080 35952 35086
rect 35900 35022 35952 35028
rect 35624 32020 35676 32026
rect 35624 31962 35676 31968
rect 35912 30258 35940 35022
rect 36084 32360 36136 32366
rect 36084 32302 36136 32308
rect 35992 31816 36044 31822
rect 35992 31758 36044 31764
rect 35900 30252 35952 30258
rect 35900 30194 35952 30200
rect 36004 28558 36032 31758
rect 36096 31482 36124 32302
rect 36084 31476 36136 31482
rect 36084 31418 36136 31424
rect 35992 28552 36044 28558
rect 35992 28494 36044 28500
rect 36004 27130 36032 28494
rect 35992 27124 36044 27130
rect 35992 27066 36044 27072
rect 35532 26308 35584 26314
rect 35532 26250 35584 26256
rect 35544 24818 35572 26250
rect 35532 24812 35584 24818
rect 35532 24754 35584 24760
rect 36084 24676 36136 24682
rect 36084 24618 36136 24624
rect 35992 24608 36044 24614
rect 35992 24550 36044 24556
rect 35900 23724 35952 23730
rect 35900 23666 35952 23672
rect 35440 23520 35492 23526
rect 35440 23462 35492 23468
rect 35912 23118 35940 23666
rect 35900 23112 35952 23118
rect 35900 23054 35952 23060
rect 35348 22976 35400 22982
rect 35348 22918 35400 22924
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 35900 21888 35952 21894
rect 35900 21830 35952 21836
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 35716 20936 35768 20942
rect 35716 20878 35768 20884
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34152 15972 34204 15978
rect 34152 15914 34204 15920
rect 33140 3392 33192 3398
rect 33140 3334 33192 3340
rect 33152 2922 33180 3334
rect 33140 2916 33192 2922
rect 33140 2858 33192 2864
rect 34164 2650 34192 15914
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34520 15700 34572 15706
rect 34520 15642 34572 15648
rect 34532 13938 34560 15642
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34520 13932 34572 13938
rect 34520 13874 34572 13880
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34888 3460 34940 3466
rect 34888 3402 34940 3408
rect 34900 3058 34928 3402
rect 34888 3052 34940 3058
rect 34888 2994 34940 3000
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 32404 2644 32456 2650
rect 32404 2586 32456 2592
rect 34152 2644 34204 2650
rect 34152 2586 34204 2592
rect 35728 2514 35756 20878
rect 35912 6458 35940 21830
rect 36004 21554 36032 24550
rect 36096 23746 36124 24618
rect 36188 23866 36216 36722
rect 36740 36378 36768 39200
rect 36728 36372 36780 36378
rect 36728 36314 36780 36320
rect 36268 35488 36320 35494
rect 36266 35456 36268 35465
rect 36320 35456 36322 35465
rect 36266 35391 36322 35400
rect 36452 33448 36504 33454
rect 36266 33416 36322 33425
rect 36452 33390 36504 33396
rect 36266 33351 36268 33360
rect 36320 33351 36322 33360
rect 36268 33322 36320 33328
rect 36360 32768 36412 32774
rect 36360 32710 36412 32716
rect 36372 32366 36400 32710
rect 36360 32360 36412 32366
rect 36360 32302 36412 32308
rect 36372 32065 36400 32302
rect 36358 32056 36414 32065
rect 36358 31991 36414 32000
rect 36360 30184 36412 30190
rect 36360 30126 36412 30132
rect 36372 30025 36400 30126
rect 36358 30016 36414 30025
rect 36358 29951 36414 29960
rect 36372 29850 36400 29951
rect 36360 29844 36412 29850
rect 36360 29786 36412 29792
rect 36464 28082 36492 33390
rect 36452 28076 36504 28082
rect 36452 28018 36504 28024
rect 36360 28008 36412 28014
rect 36358 27976 36360 27985
rect 36412 27976 36414 27985
rect 36358 27911 36414 27920
rect 36372 27674 36400 27911
rect 36360 27668 36412 27674
rect 36360 27610 36412 27616
rect 36464 27470 36492 28018
rect 36452 27464 36504 27470
rect 36452 27406 36504 27412
rect 36360 26988 36412 26994
rect 36360 26930 36412 26936
rect 36372 26625 36400 26930
rect 36358 26616 36414 26625
rect 36358 26551 36414 26560
rect 36268 24608 36320 24614
rect 36266 24576 36268 24585
rect 36320 24576 36322 24585
rect 36266 24511 36322 24520
rect 36176 23860 36228 23866
rect 36176 23802 36228 23808
rect 36096 23718 36216 23746
rect 36084 22636 36136 22642
rect 36084 22578 36136 22584
rect 35992 21548 36044 21554
rect 35992 21490 36044 21496
rect 36096 21146 36124 22578
rect 36084 21140 36136 21146
rect 36084 21082 36136 21088
rect 36188 16114 36216 23718
rect 36452 23112 36504 23118
rect 36452 23054 36504 23060
rect 36266 22536 36322 22545
rect 36266 22471 36268 22480
rect 36320 22471 36322 22480
rect 36268 22442 36320 22448
rect 36268 21344 36320 21350
rect 36268 21286 36320 21292
rect 36280 21185 36308 21286
rect 36266 21176 36322 21185
rect 36266 21111 36322 21120
rect 36266 17096 36322 17105
rect 36266 17031 36268 17040
rect 36320 17031 36322 17040
rect 36268 17002 36320 17008
rect 36176 16108 36228 16114
rect 36176 16050 36228 16056
rect 36360 16040 36412 16046
rect 36360 15982 36412 15988
rect 36372 15745 36400 15982
rect 36358 15736 36414 15745
rect 36358 15671 36360 15680
rect 36412 15671 36414 15680
rect 36360 15642 36412 15648
rect 36176 14408 36228 14414
rect 36176 14350 36228 14356
rect 36188 11558 36216 14350
rect 36268 13728 36320 13734
rect 36266 13696 36268 13705
rect 36320 13696 36322 13705
rect 36266 13631 36322 13640
rect 36360 11756 36412 11762
rect 36360 11698 36412 11704
rect 36372 11665 36400 11698
rect 36358 11656 36414 11665
rect 36358 11591 36414 11600
rect 36176 11552 36228 11558
rect 36176 11494 36228 11500
rect 36084 9376 36136 9382
rect 36084 9318 36136 9324
rect 36096 8498 36124 9318
rect 36188 8566 36216 11494
rect 36464 10674 36492 23054
rect 36452 10668 36504 10674
rect 36452 10610 36504 10616
rect 36360 10600 36412 10606
rect 36360 10542 36412 10548
rect 36372 10305 36400 10542
rect 36358 10296 36414 10305
rect 36358 10231 36360 10240
rect 36412 10231 36414 10240
rect 36360 10202 36412 10208
rect 36176 8560 36228 8566
rect 36176 8502 36228 8508
rect 36084 8492 36136 8498
rect 36084 8434 36136 8440
rect 36084 8356 36136 8362
rect 36084 8298 36136 8304
rect 36268 8356 36320 8362
rect 36268 8298 36320 8304
rect 35900 6452 35952 6458
rect 35900 6394 35952 6400
rect 36096 5234 36124 8298
rect 36280 8265 36308 8298
rect 36266 8256 36322 8265
rect 36266 8191 36322 8200
rect 36360 6316 36412 6322
rect 36360 6258 36412 6264
rect 36372 6225 36400 6258
rect 36358 6216 36414 6225
rect 36358 6151 36414 6160
rect 36084 5228 36136 5234
rect 36084 5170 36136 5176
rect 36268 5024 36320 5030
rect 36268 4966 36320 4972
rect 36280 4865 36308 4966
rect 36266 4856 36322 4865
rect 36266 4791 36322 4800
rect 36360 3936 36412 3942
rect 36360 3878 36412 3884
rect 36268 3392 36320 3398
rect 36268 3334 36320 3340
rect 36280 2825 36308 3334
rect 36372 2990 36400 3878
rect 36360 2984 36412 2990
rect 36360 2926 36412 2932
rect 37372 2984 37424 2990
rect 37372 2926 37424 2932
rect 36544 2848 36596 2854
rect 36266 2816 36322 2825
rect 36544 2790 36596 2796
rect 36266 2751 36322 2760
rect 35716 2508 35768 2514
rect 35716 2450 35768 2456
rect 35440 2440 35492 2446
rect 35440 2382 35492 2388
rect 3240 2372 3292 2378
rect 3240 2314 3292 2320
rect 9680 2372 9732 2378
rect 9680 2314 9732 2320
rect 10232 2372 10284 2378
rect 10232 2314 10284 2320
rect 13544 2372 13596 2378
rect 13544 2314 13596 2320
rect 15108 2372 15160 2378
rect 15108 2314 15160 2320
rect 21916 2372 21968 2378
rect 21916 2314 21968 2320
rect 24676 2372 24728 2378
rect 24676 2314 24728 2320
rect 32220 2372 32272 2378
rect 32220 2314 32272 2320
rect 34152 2372 34204 2378
rect 34152 2314 34204 2320
rect 2320 1352 2372 1358
rect 2320 1294 2372 1300
rect 3252 800 3280 2314
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 4540 800 4568 2246
rect 6472 800 6500 2246
rect 8404 800 8432 2246
rect 9692 800 9720 2314
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 11624 800 11652 2246
rect 13556 800 13584 2314
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 18696 2304 18748 2310
rect 18696 2246 18748 2252
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 14844 800 14872 2246
rect 16776 800 16804 2246
rect 18708 800 18736 2246
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19996 800 20024 2246
rect 21928 800 21956 2314
rect 23848 2304 23900 2310
rect 23848 2246 23900 2252
rect 25136 2304 25188 2310
rect 25136 2246 25188 2252
rect 27068 2304 27120 2310
rect 27068 2246 27120 2252
rect 29000 2304 29052 2310
rect 29000 2246 29052 2252
rect 30288 2304 30340 2310
rect 30288 2246 30340 2252
rect 23860 800 23888 2246
rect 25148 800 25176 2246
rect 27080 800 27108 2246
rect 29012 800 29040 2246
rect 30300 800 30328 2246
rect 32232 800 32260 2314
rect 34164 800 34192 2314
rect 35452 800 35480 2382
rect 18 200 74 800
rect 1306 200 1362 800
rect 3238 200 3294 800
rect 4526 200 4582 800
rect 6458 200 6514 800
rect 8390 200 8446 800
rect 9678 200 9734 800
rect 11610 200 11666 800
rect 13542 200 13598 800
rect 14830 200 14886 800
rect 16762 200 16818 800
rect 18694 200 18750 800
rect 19982 200 20038 800
rect 21914 200 21970 800
rect 23846 200 23902 800
rect 25134 200 25190 800
rect 27066 200 27122 800
rect 28998 200 29054 800
rect 30286 200 30342 800
rect 32218 200 32274 800
rect 34150 200 34206 800
rect 35438 200 35494 800
rect 36556 785 36584 2790
rect 37384 800 37412 2926
rect 36542 776 36598 785
rect 36542 711 36598 720
rect 37370 200 37426 800
<< via2 >>
rect 3422 39480 3478 39536
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4066 36080 4122 36136
rect 1490 30660 1546 30696
rect 1490 30640 1492 30660
rect 1492 30640 1544 30660
rect 1544 30640 1546 30660
rect 2226 32000 2282 32056
rect 1582 28600 1638 28656
rect 1766 26560 1822 26616
rect 1582 25236 1584 25256
rect 1584 25236 1636 25256
rect 1636 25236 1638 25256
rect 1582 25200 1638 25236
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 3790 31864 3846 31920
rect 3974 31456 4030 31512
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 5538 37304 5594 37360
rect 4986 36252 4988 36272
rect 4988 36252 5040 36272
rect 5040 36252 5042 36272
rect 4986 36216 5042 36252
rect 4894 32428 4950 32464
rect 4894 32408 4896 32428
rect 4896 32408 4948 32428
rect 4948 32408 4950 32428
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 5538 34604 5594 34640
rect 5538 34584 5540 34604
rect 5540 34584 5592 34604
rect 5592 34584 5594 34604
rect 5446 32852 5448 32872
rect 5448 32852 5500 32872
rect 5500 32852 5502 32872
rect 5446 32816 5502 32852
rect 5446 32408 5502 32464
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 1674 23160 1730 23216
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 1674 21120 1730 21176
rect 1674 19760 1730 19816
rect 1582 17756 1584 17776
rect 1584 17756 1636 17776
rect 1636 17756 1638 17776
rect 1582 17720 1638 17756
rect 1674 15680 1730 15736
rect 1674 14340 1730 14376
rect 1674 14320 1676 14340
rect 1676 14320 1728 14340
rect 1728 14320 1730 14340
rect 1674 12280 1730 12336
rect 1674 10240 1730 10296
rect 1582 8916 1584 8936
rect 1584 8916 1636 8936
rect 1636 8916 1638 8936
rect 1582 8880 1638 8916
rect 1674 6840 1730 6896
rect 1582 4800 1638 4856
rect 1674 3440 1730 3496
rect 2502 18828 2558 18864
rect 2502 18808 2504 18828
rect 2504 18808 2556 18828
rect 2556 18808 2558 18828
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 6550 35944 6606 36000
rect 6642 35264 6698 35320
rect 6550 31900 6552 31920
rect 6552 31900 6604 31920
rect 6604 31900 6606 31920
rect 6550 31864 6606 31900
rect 7378 35284 7434 35320
rect 7378 35264 7380 35284
rect 7380 35264 7432 35284
rect 7432 35264 7434 35284
rect 8482 36216 8538 36272
rect 7746 32816 7802 32872
rect 7378 29144 7434 29200
rect 5906 21936 5962 21992
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 9586 34584 9642 34640
rect 10506 35264 10562 35320
rect 10690 34992 10746 35048
rect 9218 31456 9274 31512
rect 10414 34584 10470 34640
rect 10046 29008 10102 29064
rect 10322 29144 10378 29200
rect 12622 35264 12678 35320
rect 11334 28484 11390 28520
rect 11334 28464 11336 28484
rect 11336 28464 11388 28484
rect 11388 28464 11390 28484
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 1674 1400 1730 1456
rect 11886 29008 11942 29064
rect 12254 28600 12310 28656
rect 13266 34992 13322 35048
rect 14646 28600 14702 28656
rect 14738 28056 14794 28112
rect 15290 28464 15346 28520
rect 18050 29008 18106 29064
rect 18694 28076 18750 28112
rect 18694 28056 18696 28076
rect 18696 28056 18748 28076
rect 18748 28056 18750 28076
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 35806 38800 35862 38856
rect 35622 37440 35678 37496
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 36266 35436 36268 35456
rect 36268 35436 36320 35456
rect 36320 35436 36322 35456
rect 36266 35400 36322 35436
rect 36266 33380 36322 33416
rect 36266 33360 36268 33380
rect 36268 33360 36320 33380
rect 36320 33360 36322 33380
rect 36358 32000 36414 32056
rect 36358 29960 36414 30016
rect 36358 27956 36360 27976
rect 36360 27956 36412 27976
rect 36412 27956 36414 27976
rect 36358 27920 36414 27956
rect 36358 26560 36414 26616
rect 36266 24556 36268 24576
rect 36268 24556 36320 24576
rect 36320 24556 36322 24576
rect 36266 24520 36322 24556
rect 36266 22500 36322 22536
rect 36266 22480 36268 22500
rect 36268 22480 36320 22500
rect 36320 22480 36322 22500
rect 36266 21120 36322 21176
rect 36266 17060 36322 17096
rect 36266 17040 36268 17060
rect 36268 17040 36320 17060
rect 36320 17040 36322 17060
rect 36358 15700 36414 15736
rect 36358 15680 36360 15700
rect 36360 15680 36412 15700
rect 36412 15680 36414 15700
rect 36266 13676 36268 13696
rect 36268 13676 36320 13696
rect 36320 13676 36322 13696
rect 36266 13640 36322 13676
rect 36358 11600 36414 11656
rect 36358 10260 36414 10296
rect 36358 10240 36360 10260
rect 36360 10240 36412 10260
rect 36412 10240 36414 10260
rect 36266 8200 36322 8256
rect 36358 6160 36414 6216
rect 36266 4800 36322 4856
rect 36266 2760 36322 2816
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 36542 720 36598 776
<< metal3 >>
rect 200 39538 800 39568
rect 3417 39538 3483 39541
rect 200 39536 3483 39538
rect 200 39480 3422 39536
rect 3478 39480 3483 39536
rect 200 39478 3483 39480
rect 200 39448 800 39478
rect 3417 39475 3483 39478
rect 35801 38858 35867 38861
rect 37200 38858 37800 38888
rect 35801 38856 37800 38858
rect 35801 38800 35806 38856
rect 35862 38800 37800 38856
rect 35801 38798 37800 38800
rect 35801 38795 35867 38798
rect 37200 38768 37800 38798
rect 4210 37568 4526 37569
rect 200 37498 800 37528
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 35617 37498 35683 37501
rect 37200 37498 37800 37528
rect 200 37438 4124 37498
rect 200 37408 800 37438
rect 4064 37362 4124 37438
rect 35617 37496 37800 37498
rect 35617 37440 35622 37496
rect 35678 37440 37800 37496
rect 35617 37438 37800 37440
rect 35617 37435 35683 37438
rect 37200 37408 37800 37438
rect 5533 37362 5599 37365
rect 4064 37360 5599 37362
rect 4064 37304 5538 37360
rect 5594 37304 5599 37360
rect 4064 37302 5599 37304
rect 5533 37299 5599 37302
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 4981 36274 5047 36277
rect 8477 36274 8543 36277
rect 4981 36272 8543 36274
rect 4981 36216 4986 36272
rect 5042 36216 8482 36272
rect 8538 36216 8543 36272
rect 4981 36214 8543 36216
rect 4981 36211 5047 36214
rect 8477 36211 8543 36214
rect 200 36138 800 36168
rect 4061 36138 4127 36141
rect 200 36136 4127 36138
rect 200 36080 4066 36136
rect 4122 36080 4127 36136
rect 200 36078 4127 36080
rect 200 36048 800 36078
rect 4061 36075 4127 36078
rect 5942 35940 5948 36004
rect 6012 36002 6018 36004
rect 6545 36002 6611 36005
rect 6012 36000 6611 36002
rect 6012 35944 6550 36000
rect 6606 35944 6611 36000
rect 6012 35942 6611 35944
rect 6012 35940 6018 35942
rect 6545 35939 6611 35942
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 36261 35458 36327 35461
rect 37200 35458 37800 35488
rect 36261 35456 37800 35458
rect 36261 35400 36266 35456
rect 36322 35400 37800 35456
rect 36261 35398 37800 35400
rect 36261 35395 36327 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 37200 35368 37800 35398
rect 34930 35327 35246 35328
rect 6637 35322 6703 35325
rect 7373 35322 7439 35325
rect 6637 35320 7439 35322
rect 6637 35264 6642 35320
rect 6698 35264 7378 35320
rect 7434 35264 7439 35320
rect 6637 35262 7439 35264
rect 6637 35259 6703 35262
rect 7373 35259 7439 35262
rect 10501 35322 10567 35325
rect 12617 35322 12683 35325
rect 10501 35320 12683 35322
rect 10501 35264 10506 35320
rect 10562 35264 12622 35320
rect 12678 35264 12683 35320
rect 10501 35262 12683 35264
rect 10501 35259 10567 35262
rect 12617 35259 12683 35262
rect 10685 35050 10751 35053
rect 13261 35050 13327 35053
rect 10685 35048 13327 35050
rect 10685 34992 10690 35048
rect 10746 34992 13266 35048
rect 13322 34992 13327 35048
rect 10685 34990 13327 34992
rect 10685 34987 10751 34990
rect 13261 34987 13327 34990
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 5533 34642 5599 34645
rect 9581 34642 9647 34645
rect 5533 34640 9647 34642
rect 5533 34584 5538 34640
rect 5594 34584 9586 34640
rect 9642 34584 9647 34640
rect 5533 34582 9647 34584
rect 5533 34579 5599 34582
rect 9581 34579 9647 34582
rect 10409 34642 10475 34645
rect 10542 34642 10548 34644
rect 10409 34640 10548 34642
rect 10409 34584 10414 34640
rect 10470 34584 10548 34640
rect 10409 34582 10548 34584
rect 10409 34579 10475 34582
rect 10542 34580 10548 34582
rect 10612 34580 10618 34644
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 200 34008 800 34128
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 36261 33418 36327 33421
rect 37200 33418 37800 33448
rect 36261 33416 37800 33418
rect 36261 33360 36266 33416
rect 36322 33360 37800 33416
rect 36261 33358 37800 33360
rect 36261 33355 36327 33358
rect 37200 33328 37800 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 5441 32874 5507 32877
rect 7741 32874 7807 32877
rect 5441 32872 7807 32874
rect 5441 32816 5446 32872
rect 5502 32816 7746 32872
rect 7802 32816 7807 32872
rect 5441 32814 7807 32816
rect 5441 32811 5507 32814
rect 7741 32811 7807 32814
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4889 32466 4955 32469
rect 5441 32466 5507 32469
rect 4889 32464 5507 32466
rect 4889 32408 4894 32464
rect 4950 32408 5446 32464
rect 5502 32408 5507 32464
rect 4889 32406 5507 32408
rect 4889 32403 4955 32406
rect 5441 32403 5507 32406
rect 4210 32128 4526 32129
rect 200 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 2221 32058 2287 32061
rect 200 32056 2287 32058
rect 200 32000 2226 32056
rect 2282 32000 2287 32056
rect 200 31998 2287 32000
rect 200 31968 800 31998
rect 2221 31995 2287 31998
rect 36353 32058 36419 32061
rect 37200 32058 37800 32088
rect 36353 32056 37800 32058
rect 36353 32000 36358 32056
rect 36414 32000 37800 32056
rect 36353 31998 37800 32000
rect 36353 31995 36419 31998
rect 37200 31968 37800 31998
rect 3785 31922 3851 31925
rect 6545 31922 6611 31925
rect 3785 31920 6611 31922
rect 3785 31864 3790 31920
rect 3846 31864 6550 31920
rect 6606 31864 6611 31920
rect 3785 31862 6611 31864
rect 3785 31859 3851 31862
rect 6545 31859 6611 31862
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 3969 31514 4035 31517
rect 9213 31514 9279 31517
rect 3969 31512 9279 31514
rect 3969 31456 3974 31512
rect 4030 31456 9218 31512
rect 9274 31456 9279 31512
rect 3969 31454 9279 31456
rect 3969 31451 4035 31454
rect 9213 31451 9279 31454
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 200 30698 800 30728
rect 1485 30698 1551 30701
rect 200 30696 1551 30698
rect 200 30640 1490 30696
rect 1546 30640 1551 30696
rect 200 30638 1551 30640
rect 200 30608 800 30638
rect 1485 30635 1551 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 36353 30018 36419 30021
rect 37200 30018 37800 30048
rect 36353 30016 37800 30018
rect 36353 29960 36358 30016
rect 36414 29960 37800 30016
rect 36353 29958 37800 29960
rect 36353 29955 36419 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 37200 29928 37800 29958
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 7373 29202 7439 29205
rect 10317 29202 10383 29205
rect 7373 29200 10383 29202
rect 7373 29144 7378 29200
rect 7434 29144 10322 29200
rect 10378 29144 10383 29200
rect 7373 29142 10383 29144
rect 7373 29139 7439 29142
rect 10317 29139 10383 29142
rect 10041 29066 10107 29069
rect 11881 29066 11947 29069
rect 18045 29066 18111 29069
rect 10041 29064 18111 29066
rect 10041 29008 10046 29064
rect 10102 29008 11886 29064
rect 11942 29008 18050 29064
rect 18106 29008 18111 29064
rect 10041 29006 18111 29008
rect 10041 29003 10107 29006
rect 11881 29003 11947 29006
rect 18045 29003 18111 29006
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 200 28658 800 28688
rect 1577 28658 1643 28661
rect 200 28656 1643 28658
rect 200 28600 1582 28656
rect 1638 28600 1643 28656
rect 200 28598 1643 28600
rect 200 28568 800 28598
rect 1577 28595 1643 28598
rect 12249 28658 12315 28661
rect 14641 28658 14707 28661
rect 12249 28656 14707 28658
rect 12249 28600 12254 28656
rect 12310 28600 14646 28656
rect 14702 28600 14707 28656
rect 12249 28598 14707 28600
rect 12249 28595 12315 28598
rect 14641 28595 14707 28598
rect 11329 28522 11395 28525
rect 15285 28522 15351 28525
rect 11329 28520 15351 28522
rect 11329 28464 11334 28520
rect 11390 28464 15290 28520
rect 15346 28464 15351 28520
rect 11329 28462 15351 28464
rect 11329 28459 11395 28462
rect 15285 28459 15351 28462
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 14733 28114 14799 28117
rect 18689 28114 18755 28117
rect 14733 28112 18755 28114
rect 14733 28056 14738 28112
rect 14794 28056 18694 28112
rect 18750 28056 18755 28112
rect 14733 28054 18755 28056
rect 14733 28051 14799 28054
rect 18689 28051 18755 28054
rect 36353 27978 36419 27981
rect 37200 27978 37800 28008
rect 36353 27976 37800 27978
rect 36353 27920 36358 27976
rect 36414 27920 37800 27976
rect 36353 27918 37800 27920
rect 36353 27915 36419 27918
rect 37200 27888 37800 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 200 26618 800 26648
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 1761 26618 1827 26621
rect 200 26616 1827 26618
rect 200 26560 1766 26616
rect 1822 26560 1827 26616
rect 200 26558 1827 26560
rect 200 26528 800 26558
rect 1761 26555 1827 26558
rect 36353 26618 36419 26621
rect 37200 26618 37800 26648
rect 36353 26616 37800 26618
rect 36353 26560 36358 26616
rect 36414 26560 37800 26616
rect 36353 26558 37800 26560
rect 36353 26555 36419 26558
rect 37200 26528 37800 26558
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 200 25258 800 25288
rect 1577 25258 1643 25261
rect 200 25256 1643 25258
rect 200 25200 1582 25256
rect 1638 25200 1643 25256
rect 200 25198 1643 25200
rect 200 25168 800 25198
rect 1577 25195 1643 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 36261 24578 36327 24581
rect 37200 24578 37800 24608
rect 36261 24576 37800 24578
rect 36261 24520 36266 24576
rect 36322 24520 37800 24576
rect 36261 24518 37800 24520
rect 36261 24515 36327 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 37200 24488 37800 24518
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 200 23218 800 23248
rect 1669 23218 1735 23221
rect 200 23216 1735 23218
rect 200 23160 1674 23216
rect 1730 23160 1735 23216
rect 200 23158 1735 23160
rect 200 23128 800 23158
rect 1669 23155 1735 23158
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 36261 22538 36327 22541
rect 37200 22538 37800 22568
rect 36261 22536 37800 22538
rect 36261 22480 36266 22536
rect 36322 22480 37800 22536
rect 36261 22478 37800 22480
rect 36261 22475 36327 22478
rect 37200 22448 37800 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 5901 21996 5967 21997
rect 5901 21994 5948 21996
rect 5856 21992 5948 21994
rect 5856 21936 5906 21992
rect 5856 21934 5948 21936
rect 5901 21932 5948 21934
rect 6012 21932 6018 21996
rect 5901 21931 5967 21932
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 200 21178 800 21208
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 1669 21178 1735 21181
rect 200 21176 1735 21178
rect 200 21120 1674 21176
rect 1730 21120 1735 21176
rect 200 21118 1735 21120
rect 200 21088 800 21118
rect 1669 21115 1735 21118
rect 36261 21178 36327 21181
rect 37200 21178 37800 21208
rect 36261 21176 37800 21178
rect 36261 21120 36266 21176
rect 36322 21120 37800 21176
rect 36261 21118 37800 21120
rect 36261 21115 36327 21118
rect 37200 21088 37800 21118
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 200 19818 800 19848
rect 1669 19818 1735 19821
rect 200 19816 1735 19818
rect 200 19760 1674 19816
rect 1730 19760 1735 19816
rect 200 19758 1735 19760
rect 200 19728 800 19758
rect 1669 19755 1735 19758
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 37200 19048 37800 19168
rect 34930 19007 35246 19008
rect 2497 18866 2563 18869
rect 10542 18866 10548 18868
rect 2497 18864 10548 18866
rect 2497 18808 2502 18864
rect 2558 18808 10548 18864
rect 2497 18806 10548 18808
rect 2497 18803 2563 18806
rect 10542 18804 10548 18806
rect 10612 18804 10618 18868
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 200 17778 800 17808
rect 1577 17778 1643 17781
rect 200 17776 1643 17778
rect 200 17720 1582 17776
rect 1638 17720 1643 17776
rect 200 17718 1643 17720
rect 200 17688 800 17718
rect 1577 17715 1643 17718
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 36261 17098 36327 17101
rect 37200 17098 37800 17128
rect 36261 17096 37800 17098
rect 36261 17040 36266 17096
rect 36322 17040 37800 17096
rect 36261 17038 37800 17040
rect 36261 17035 36327 17038
rect 37200 17008 37800 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 200 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 1669 15738 1735 15741
rect 200 15736 1735 15738
rect 200 15680 1674 15736
rect 1730 15680 1735 15736
rect 200 15678 1735 15680
rect 200 15648 800 15678
rect 1669 15675 1735 15678
rect 36353 15738 36419 15741
rect 37200 15738 37800 15768
rect 36353 15736 37800 15738
rect 36353 15680 36358 15736
rect 36414 15680 37800 15736
rect 36353 15678 37800 15680
rect 36353 15675 36419 15678
rect 37200 15648 37800 15678
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 200 14378 800 14408
rect 1669 14378 1735 14381
rect 200 14376 1735 14378
rect 200 14320 1674 14376
rect 1730 14320 1735 14376
rect 200 14318 1735 14320
rect 200 14288 800 14318
rect 1669 14315 1735 14318
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 36261 13698 36327 13701
rect 37200 13698 37800 13728
rect 36261 13696 37800 13698
rect 36261 13640 36266 13696
rect 36322 13640 37800 13696
rect 36261 13638 37800 13640
rect 36261 13635 36327 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 37200 13608 37800 13638
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 200 12338 800 12368
rect 1669 12338 1735 12341
rect 200 12336 1735 12338
rect 200 12280 1674 12336
rect 1730 12280 1735 12336
rect 200 12278 1735 12280
rect 200 12248 800 12278
rect 1669 12275 1735 12278
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 36353 11658 36419 11661
rect 37200 11658 37800 11688
rect 36353 11656 37800 11658
rect 36353 11600 36358 11656
rect 36414 11600 37800 11656
rect 36353 11598 37800 11600
rect 36353 11595 36419 11598
rect 37200 11568 37800 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 200 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 1669 10298 1735 10301
rect 200 10296 1735 10298
rect 200 10240 1674 10296
rect 1730 10240 1735 10296
rect 200 10238 1735 10240
rect 200 10208 800 10238
rect 1669 10235 1735 10238
rect 36353 10298 36419 10301
rect 37200 10298 37800 10328
rect 36353 10296 37800 10298
rect 36353 10240 36358 10296
rect 36414 10240 37800 10296
rect 36353 10238 37800 10240
rect 36353 10235 36419 10238
rect 37200 10208 37800 10238
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 200 8938 800 8968
rect 1577 8938 1643 8941
rect 200 8936 1643 8938
rect 200 8880 1582 8936
rect 1638 8880 1643 8936
rect 200 8878 1643 8880
rect 200 8848 800 8878
rect 1577 8875 1643 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 36261 8258 36327 8261
rect 37200 8258 37800 8288
rect 36261 8256 37800 8258
rect 36261 8200 36266 8256
rect 36322 8200 37800 8256
rect 36261 8198 37800 8200
rect 36261 8195 36327 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 37200 8168 37800 8198
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 200 6898 800 6928
rect 1669 6898 1735 6901
rect 200 6896 1735 6898
rect 200 6840 1674 6896
rect 1730 6840 1735 6896
rect 200 6838 1735 6840
rect 200 6808 800 6838
rect 1669 6835 1735 6838
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 36353 6218 36419 6221
rect 37200 6218 37800 6248
rect 36353 6216 37800 6218
rect 36353 6160 36358 6216
rect 36414 6160 37800 6216
rect 36353 6158 37800 6160
rect 36353 6155 36419 6158
rect 37200 6128 37800 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 200 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 1577 4858 1643 4861
rect 200 4856 1643 4858
rect 200 4800 1582 4856
rect 1638 4800 1643 4856
rect 200 4798 1643 4800
rect 200 4768 800 4798
rect 1577 4795 1643 4798
rect 36261 4858 36327 4861
rect 37200 4858 37800 4888
rect 36261 4856 37800 4858
rect 36261 4800 36266 4856
rect 36322 4800 37800 4856
rect 36261 4798 37800 4800
rect 36261 4795 36327 4798
rect 37200 4768 37800 4798
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 200 3498 800 3528
rect 1669 3498 1735 3501
rect 200 3496 1735 3498
rect 200 3440 1674 3496
rect 1730 3440 1735 3496
rect 200 3438 1735 3440
rect 200 3408 800 3438
rect 1669 3435 1735 3438
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 36261 2818 36327 2821
rect 37200 2818 37800 2848
rect 36261 2816 37800 2818
rect 36261 2760 36266 2816
rect 36322 2760 37800 2816
rect 36261 2758 37800 2760
rect 36261 2755 36327 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 37200 2728 37800 2758
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 200 1458 800 1488
rect 1669 1458 1735 1461
rect 200 1456 1735 1458
rect 200 1400 1674 1456
rect 1730 1400 1735 1456
rect 200 1398 1735 1400
rect 200 1368 800 1398
rect 1669 1395 1735 1398
rect 36537 778 36603 781
rect 37200 778 37800 808
rect 36537 776 37800 778
rect 36537 720 36542 776
rect 36598 720 37800 776
rect 36537 718 37800 720
rect 36537 715 36603 718
rect 37200 688 37800 718
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 5948 35940 6012 36004
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 10548 34580 10612 34644
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 5948 21992 6012 21996
rect 5948 21936 5962 21992
rect 5962 21936 6012 21992
rect 5948 21932 6012 21936
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 10548 18804 10612 18868
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 5947 36004 6013 36005
rect 5947 35940 5948 36004
rect 6012 35940 6013 36004
rect 5947 35939 6013 35940
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 5950 21997 6010 35939
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 10547 34644 10613 34645
rect 10547 34580 10548 34644
rect 10612 34580 10613 34644
rect 10547 34579 10613 34580
rect 5947 21996 6013 21997
rect 5947 21932 5948 21996
rect 6012 21932 6013 21996
rect 5947 21931 6013 21932
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 10550 18869 10610 34579
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 10547 18868 10613 18869
rect 10547 18804 10548 18868
rect 10612 18804 10613 18868
rect 10547 18803 10613 18804
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__137__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 19596 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1667941163
transform 1 0 11684 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__145__A
timestamp 1667941163
transform -1 0 19228 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__A
timestamp 1667941163
transform 1 0 19412 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__149__A
timestamp 1667941163
transform -1 0 20148 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__153__A
timestamp 1667941163
transform -1 0 19780 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__157__A
timestamp 1667941163
transform 1 0 9752 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__A
timestamp 1667941163
transform -1 0 12788 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__161__A
timestamp 1667941163
transform -1 0 12236 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__162__A
timestamp 1667941163
transform 1 0 16836 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__165__A
timestamp 1667941163
transform 1 0 10948 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__166__A
timestamp 1667941163
transform -1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__A
timestamp 1667941163
transform 1 0 16100 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__A
timestamp 1667941163
transform -1 0 18860 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__A
timestamp 1667941163
transform 1 0 9108 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__A
timestamp 1667941163
transform 1 0 14260 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__185__A
timestamp 1667941163
transform 1 0 14996 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__A
timestamp 1667941163
transform 1 0 18492 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__188__A
timestamp 1667941163
transform -1 0 17664 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__A
timestamp 1667941163
transform 1 0 9660 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A
timestamp 1667941163
transform -1 0 20332 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__A
timestamp 1667941163
transform 1 0 8372 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A
timestamp 1667941163
transform 1 0 8464 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__A
timestamp 1667941163
transform 1 0 10212 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__A
timestamp 1667941163
transform 1 0 8096 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__A
timestamp 1667941163
transform -1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__198__A
timestamp 1667941163
transform -1 0 15088 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__200__A
timestamp 1667941163
transform 1 0 11684 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__201__A
timestamp 1667941163
transform -1 0 16836 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__202__A
timestamp 1667941163
transform 1 0 13616 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__A
timestamp 1667941163
transform 1 0 18676 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__A
timestamp 1667941163
transform -1 0 19872 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__A
timestamp 1667941163
transform -1 0 8648 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__215__A
timestamp 1667941163
transform -1 0 19320 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__217__A
timestamp 1667941163
transform -1 0 20148 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A
timestamp 1667941163
transform -1 0 7728 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__221__A
timestamp 1667941163
transform -1 0 14444 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__A
timestamp 1667941163
transform 1 0 19412 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__A
timestamp 1667941163
transform -1 0 31280 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__232__A
timestamp 1667941163
transform -1 0 17756 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__233__A
timestamp 1667941163
transform 1 0 18860 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__A
timestamp 1667941163
transform 1 0 16836 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__A
timestamp 1667941163
transform 1 0 15732 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__238__A
timestamp 1667941163
transform -1 0 35696 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__A
timestamp 1667941163
transform 1 0 23276 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A
timestamp 1667941163
transform -1 0 7360 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__242__A
timestamp 1667941163
transform 1 0 12972 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A
timestamp 1667941163
transform -1 0 9936 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__A
timestamp 1667941163
transform 1 0 5244 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__A
timestamp 1667941163
transform -1 0 35604 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__248__A
timestamp 1667941163
transform -1 0 11868 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__249__A
timestamp 1667941163
transform 1 0 15548 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__250__A
timestamp 1667941163
transform -1 0 23828 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__254__A
timestamp 1667941163
transform 1 0 14260 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__A
timestamp 1667941163
transform 1 0 12052 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__A
timestamp 1667941163
transform 1 0 14812 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__A
timestamp 1667941163
transform 1 0 16468 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__A
timestamp 1667941163
transform 1 0 13524 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__A
timestamp 1667941163
transform -1 0 14720 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__300__A
timestamp 1667941163
transform 1 0 12328 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__301__A
timestamp 1667941163
transform 1 0 14812 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__302__CLK
timestamp 1667941163
transform 1 0 9108 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__303__CLK
timestamp 1667941163
transform 1 0 4048 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__304__CLK
timestamp 1667941163
transform 1 0 3496 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__304__D
timestamp 1667941163
transform 1 0 4784 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__305__CLK
timestamp 1667941163
transform 1 0 10764 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__306__CLK
timestamp 1667941163
transform 1 0 9108 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__307__CLK
timestamp 1667941163
transform 1 0 4508 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__307__D
timestamp 1667941163
transform -1 0 5520 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__308__CLK
timestamp 1667941163
transform 1 0 15088 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__309__CLK
timestamp 1667941163
transform 1 0 15272 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__310__CLK
timestamp 1667941163
transform 1 0 15364 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__310__D
timestamp 1667941163
transform -1 0 16100 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__311__CLK
timestamp 1667941163
transform 1 0 14260 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__311__D
timestamp 1667941163
transform 1 0 12972 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__312__CLK
timestamp 1667941163
transform 1 0 13524 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__312__D
timestamp 1667941163
transform 1 0 10764 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__313__CLK
timestamp 1667941163
transform 1 0 11408 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__314__CLK
timestamp 1667941163
transform -1 0 3956 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__315__CLK
timestamp 1667941163
transform -1 0 4508 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__316__CLK
timestamp 1667941163
transform 1 0 5060 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__316__D
timestamp 1667941163
transform 1 0 14260 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__317__CLK
timestamp 1667941163
transform 1 0 14812 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__317__D
timestamp 1667941163
transform -1 0 6072 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__318__CLK
timestamp 1667941163
transform 1 0 15180 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__318__D
timestamp 1667941163
transform 1 0 14076 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__319__CLK
timestamp 1667941163
transform 1 0 15916 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__320__CLK
timestamp 1667941163
transform 1 0 14720 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__321__CLK
timestamp 1667941163
transform -1 0 16284 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__322__CLK
timestamp 1667941163
transform 1 0 14260 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__323__CLK
timestamp 1667941163
transform 1 0 12972 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__324__CLK
timestamp 1667941163
transform 1 0 5244 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__325__CLK
timestamp 1667941163
transform 1 0 4048 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__326__CLK
timestamp 1667941163
transform 1 0 5796 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__327__CLK
timestamp 1667941163
transform 1 0 5336 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__328__CLK
timestamp 1667941163
transform 1 0 3956 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__328__D
timestamp 1667941163
transform 1 0 5888 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__329__CLK
timestamp 1667941163
transform 1 0 14260 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__329__D
timestamp 1667941163
transform 1 0 13524 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__330__CLK
timestamp 1667941163
transform 1 0 13524 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__331__CLK
timestamp 1667941163
transform 1 0 11960 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__332__CLK
timestamp 1667941163
transform 1 0 4692 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__333__CLK
timestamp 1667941163
transform 1 0 10580 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__334__CLK
timestamp 1667941163
transform 1 0 5888 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__334__D
timestamp 1667941163
transform -1 0 6072 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__CLK
timestamp 1667941163
transform 1 0 3956 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__336__CLK
timestamp 1667941163
transform 1 0 9660 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__337__CLK
timestamp 1667941163
transform 1 0 6532 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__338__CLK
timestamp 1667941163
transform 1 0 15732 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__CLK
timestamp 1667941163
transform 1 0 15824 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__340__CLK
timestamp 1667941163
transform 1 0 14628 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__CLK
timestamp 1667941163
transform 1 0 14720 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__D
timestamp 1667941163
transform 1 0 12512 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__CLK
timestamp 1667941163
transform 1 0 10212 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__CLK
timestamp 1667941163
transform 1 0 15272 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__352__A
timestamp 1667941163
transform 1 0 15548 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__353__A
timestamp 1667941163
transform 1 0 2944 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__354__A
timestamp 1667941163
transform 1 0 12328 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__A
timestamp 1667941163
transform -1 0 32568 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__357__A
timestamp 1667941163
transform 1 0 19228 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__358__A
timestamp 1667941163
transform -1 0 27968 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__359__A
timestamp 1667941163
transform 1 0 2576 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__360__A
timestamp 1667941163
transform 1 0 22080 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__363__A
timestamp 1667941163
transform -1 0 25668 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__365__A
timestamp 1667941163
transform -1 0 26220 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__369__A
timestamp 1667941163
transform -1 0 6532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__372__A
timestamp 1667941163
transform -1 0 28704 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__373__A
timestamp 1667941163
transform -1 0 17204 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__374__A
timestamp 1667941163
transform 1 0 2392 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__380__A
timestamp 1667941163
transform 1 0 21804 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__381__A
timestamp 1667941163
transform -1 0 35512 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__382__A
timestamp 1667941163
transform 1 0 14260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__383__A
timestamp 1667941163
transform -1 0 13984 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__A
timestamp 1667941163
transform 1 0 6992 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__385__A
timestamp 1667941163
transform -1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__386__A
timestamp 1667941163
transform 1 0 11408 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__403__A
timestamp 1667941163
transform -1 0 17756 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__423__A
timestamp 1667941163
transform 1 0 19412 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__431__A
timestamp 1667941163
transform 1 0 17940 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1667941163
transform -1 0 36432 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1667941163
transform -1 0 17664 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1667941163
transform -1 0 15732 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1667941163
transform -1 0 36432 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1667941163
transform -1 0 15548 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1667941163
transform -1 0 2392 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1667941163
transform -1 0 11224 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1667941163
transform -1 0 14444 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1667941163
transform -1 0 36432 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1667941163
transform -1 0 1748 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1667941163
transform -1 0 35788 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1667941163
transform -1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1667941163
transform -1 0 35144 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1667941163
transform -1 0 1748 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1667941163
transform -1 0 1748 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1667941163
transform -1 0 24840 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1667941163
transform -1 0 35052 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1667941163
transform -1 0 33672 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1667941163
transform -1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1667941163
transform -1 0 36432 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1667941163
transform -1 0 1748 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1667941163
transform -1 0 4140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1667941163
transform -1 0 10396 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1667941163
transform -1 0 32476 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1667941163
transform -1 0 35788 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1667941163
transform -1 0 35788 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1667941163
transform -1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1667941163
transform -1 0 14168 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1667941163
transform -1 0 36432 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1667941163
transform -1 0 8648 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1667941163
transform -1 0 36432 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1667941163
transform -1 0 2392 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1667941163
transform -1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1667941163
transform -1 0 1748 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1667941163
transform -1 0 2300 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1667941163
transform -1 0 12604 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1667941163
transform -1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1667941163
transform -1 0 2484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1667941163
transform -1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1667941163
transform -1 0 29992 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output45_A
timestamp 1667941163
transform -1 0 35696 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output51_A
timestamp 1667941163
transform -1 0 28060 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output64_A
timestamp 1667941163
transform 1 0 35512 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output71_A
timestamp 1667941163
transform -1 0 35696 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output73_A
timestamp 1667941163
transform 1 0 16192 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output75_A
timestamp 1667941163
transform -1 0 35696 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output82_A
timestamp 1667941163
transform 1 0 20792 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2576 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1667941163
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33
timestamp 1667941163
transform 1 0 4140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4968 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1667941163
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63
timestamp 1667941163
transform 1 0 6900 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75
timestamp 1667941163
transform 1 0 8004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79
timestamp 1667941163
transform 1 0 8372 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1667941163
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97
timestamp 1667941163
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105
timestamp 1667941163
transform 1 0 10764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1667941163
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119
timestamp 1667941163
transform 1 0 12052 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_131 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 13156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1667941163
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_145
timestamp 1667941163
transform 1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_149
timestamp 1667941163
transform 1 0 14812 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_154 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 15272 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_162
timestamp 1667941163
transform 1 0 16008 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1667941163
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_175
timestamp 1667941163
transform 1 0 17204 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1667941163
transform 1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_191
timestamp 1667941163
transform 1 0 18676 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1667941163
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_202
timestamp 1667941163
transform 1 0 19688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_210
timestamp 1667941163
transform 1 0 20424 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_216
timestamp 1667941163
transform 1 0 20976 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1667941163
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_231
timestamp 1667941163
transform 1 0 22356 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_243
timestamp 1667941163
transform 1 0 23460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_247
timestamp 1667941163
transform 1 0 23828 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1667941163
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_265
timestamp 1667941163
transform 1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273
timestamp 1667941163
transform 1 0 26220 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1667941163
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_287
timestamp 1667941163
transform 1 0 27508 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_299
timestamp 1667941163
transform 1 0 28612 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_303
timestamp 1667941163
transform 1 0 28980 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1667941163
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_321
timestamp 1667941163
transform 1 0 30636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_329
timestamp 1667941163
transform 1 0 31372 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1667941163
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_343
timestamp 1667941163
transform 1 0 32660 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_351
timestamp 1667941163
transform 1 0 33396 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_354
timestamp 1667941163
transform 1 0 33672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_362
timestamp 1667941163
transform 1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_369
timestamp 1667941163
transform 1 0 35052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_373
timestamp 1667941163
transform 1 0 35420 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_384
timestamp 1667941163
transform 1 0 36432 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1667941163
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1667941163
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1667941163
transform 1 0 3588 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_34
timestamp 1667941163
transform 1 0 4232 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_46
timestamp 1667941163
transform 1 0 5336 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1667941163
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1667941163
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1667941163
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_93
timestamp 1667941163
transform 1 0 9660 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_101
timestamp 1667941163
transform 1 0 10396 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_109
timestamp 1667941163
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_118
timestamp 1667941163
transform 1 0 11960 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_124
timestamp 1667941163
transform 1 0 12512 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_136
timestamp 1667941163
transform 1 0 13616 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_148
timestamp 1667941163
transform 1 0 14720 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_156
timestamp 1667941163
transform 1 0 15456 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1667941163
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1667941163
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1667941163
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_193
timestamp 1667941163
transform 1 0 18860 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_197
timestamp 1667941163
transform 1 0 19228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_201
timestamp 1667941163
transform 1 0 19596 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_207
timestamp 1667941163
transform 1 0 20148 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_219
timestamp 1667941163
transform 1 0 21252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1667941163
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_237
timestamp 1667941163
transform 1 0 22908 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_241
timestamp 1667941163
transform 1 0 23276 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_247
timestamp 1667941163
transform 1 0 23828 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_259
timestamp 1667941163
transform 1 0 24932 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_271
timestamp 1667941163
transform 1 0 26036 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1667941163
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1667941163
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1667941163
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1667941163
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1667941163
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1667941163
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_341
timestamp 1667941163
transform 1 0 32476 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_350
timestamp 1667941163
transform 1 0 33304 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_362
timestamp 1667941163
transform 1 0 34408 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_370
timestamp 1667941163
transform 1 0 35144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_384
timestamp 1667941163
transform 1 0 36432 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_9
timestamp 1667941163
transform 1 0 1932 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_16
timestamp 1667941163
transform 1 0 2576 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1667941163
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1667941163
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1667941163
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1667941163
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1667941163
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1667941163
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1667941163
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1667941163
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1667941163
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_149
timestamp 1667941163
transform 1 0 14812 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_153
timestamp 1667941163
transform 1 0 15180 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_159
timestamp 1667941163
transform 1 0 15732 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_171
timestamp 1667941163
transform 1 0 16836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_183
timestamp 1667941163
transform 1 0 17940 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1667941163
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1667941163
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1667941163
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1667941163
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1667941163
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1667941163
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1667941163
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1667941163
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1667941163
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1667941163
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1667941163
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1667941163
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1667941163
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1667941163
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1667941163
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1667941163
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_373
timestamp 1667941163
transform 1 0 35420 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_376
timestamp 1667941163
transform 1 0 35696 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_384
timestamp 1667941163
transform 1 0 36432 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1667941163
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1667941163
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1667941163
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1667941163
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1667941163
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1667941163
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1667941163
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1667941163
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1667941163
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1667941163
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1667941163
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1667941163
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1667941163
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1667941163
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1667941163
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1667941163
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1667941163
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1667941163
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1667941163
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1667941163
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1667941163
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1667941163
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1667941163
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1667941163
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1667941163
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1667941163
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1667941163
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1667941163
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1667941163
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1667941163
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1667941163
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_373
timestamp 1667941163
transform 1 0 35420 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_381
timestamp 1667941163
transform 1 0 36156 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_384
timestamp 1667941163
transform 1 0 36432 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1667941163
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1667941163
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1667941163
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1667941163
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1667941163
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1667941163
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1667941163
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1667941163
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1667941163
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1667941163
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1667941163
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1667941163
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1667941163
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1667941163
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1667941163
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1667941163
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1667941163
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1667941163
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1667941163
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1667941163
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1667941163
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1667941163
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1667941163
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1667941163
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1667941163
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1667941163
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1667941163
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1667941163
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1667941163
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1667941163
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1667941163
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_385
timestamp 1667941163
transform 1 0 36524 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_8
timestamp 1667941163
transform 1 0 1840 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_14
timestamp 1667941163
transform 1 0 2392 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_26
timestamp 1667941163
transform 1 0 3496 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_38
timestamp 1667941163
transform 1 0 4600 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_50
timestamp 1667941163
transform 1 0 5704 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1667941163
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1667941163
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1667941163
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1667941163
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1667941163
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1667941163
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1667941163
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1667941163
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1667941163
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1667941163
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1667941163
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1667941163
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1667941163
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1667941163
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1667941163
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1667941163
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1667941163
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1667941163
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1667941163
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1667941163
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1667941163
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1667941163
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1667941163
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1667941163
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1667941163
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1667941163
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1667941163
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_373
timestamp 1667941163
transform 1 0 35420 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_379
timestamp 1667941163
transform 1 0 35972 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_384
timestamp 1667941163
transform 1 0 36432 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1667941163
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1667941163
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1667941163
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1667941163
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1667941163
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1667941163
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1667941163
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1667941163
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1667941163
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1667941163
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1667941163
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1667941163
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1667941163
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1667941163
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1667941163
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1667941163
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1667941163
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1667941163
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1667941163
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1667941163
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1667941163
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1667941163
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1667941163
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1667941163
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1667941163
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1667941163
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1667941163
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1667941163
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1667941163
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1667941163
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1667941163
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1667941163
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_377
timestamp 1667941163
transform 1 0 35788 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_385
timestamp 1667941163
transform 1 0 36524 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1667941163
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1667941163
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1667941163
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1667941163
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1667941163
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1667941163
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1667941163
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1667941163
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1667941163
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1667941163
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1667941163
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1667941163
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_149
timestamp 1667941163
transform 1 0 14812 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_153
timestamp 1667941163
transform 1 0 15180 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_159
timestamp 1667941163
transform 1 0 15732 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1667941163
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1667941163
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1667941163
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1667941163
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1667941163
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1667941163
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1667941163
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1667941163
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1667941163
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1667941163
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1667941163
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1667941163
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1667941163
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1667941163
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1667941163
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1667941163
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1667941163
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1667941163
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_373
timestamp 1667941163
transform 1 0 35420 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_377
timestamp 1667941163
transform 1 0 35788 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_384
timestamp 1667941163
transform 1 0 36432 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1667941163
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1667941163
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1667941163
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_53
timestamp 1667941163
transform 1 0 5980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_60
timestamp 1667941163
transform 1 0 6624 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_66
timestamp 1667941163
transform 1 0 7176 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_78
timestamp 1667941163
transform 1 0 8280 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1667941163
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1667941163
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1667941163
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1667941163
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1667941163
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1667941163
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1667941163
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1667941163
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1667941163
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1667941163
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1667941163
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1667941163
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1667941163
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1667941163
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1667941163
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1667941163
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1667941163
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1667941163
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1667941163
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1667941163
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1667941163
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1667941163
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1667941163
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1667941163
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1667941163
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_385
timestamp 1667941163
transform 1 0 36524 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_9
timestamp 1667941163
transform 1 0 1932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_21
timestamp 1667941163
transform 1 0 3036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_33
timestamp 1667941163
transform 1 0 4140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_45
timestamp 1667941163
transform 1 0 5244 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1667941163
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1667941163
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1667941163
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1667941163
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1667941163
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1667941163
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1667941163
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1667941163
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1667941163
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1667941163
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1667941163
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1667941163
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1667941163
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1667941163
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1667941163
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1667941163
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1667941163
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1667941163
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1667941163
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1667941163
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1667941163
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1667941163
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1667941163
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1667941163
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1667941163
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1667941163
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1667941163
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1667941163
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_385
timestamp 1667941163
transform 1 0 36524 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1667941163
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1667941163
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1667941163
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1667941163
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1667941163
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1667941163
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1667941163
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1667941163
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1667941163
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1667941163
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1667941163
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1667941163
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_153
timestamp 1667941163
transform 1 0 15180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_157
timestamp 1667941163
transform 1 0 15548 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_161
timestamp 1667941163
transform 1 0 15916 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_173
timestamp 1667941163
transform 1 0 17020 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_185
timestamp 1667941163
transform 1 0 18124 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1667941163
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1667941163
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1667941163
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1667941163
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1667941163
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1667941163
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1667941163
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1667941163
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1667941163
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1667941163
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1667941163
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1667941163
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1667941163
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1667941163
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1667941163
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1667941163
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_385
timestamp 1667941163
transform 1 0 36524 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_7
timestamp 1667941163
transform 1 0 1748 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_19
timestamp 1667941163
transform 1 0 2852 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_31
timestamp 1667941163
transform 1 0 3956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_43
timestamp 1667941163
transform 1 0 5060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1667941163
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1667941163
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1667941163
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp 1667941163
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1667941163
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1667941163
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_149
timestamp 1667941163
transform 1 0 14812 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_155
timestamp 1667941163
transform 1 0 15364 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1667941163
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1667941163
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1667941163
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1667941163
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1667941163
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1667941163
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1667941163
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1667941163
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_249
timestamp 1667941163
transform 1 0 24012 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_256
timestamp 1667941163
transform 1 0 24656 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_268
timestamp 1667941163
transform 1 0 25760 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1667941163
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1667941163
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1667941163
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1667941163
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1667941163
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1667941163
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_376
timestamp 1667941163
transform 1 0 35696 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_384
timestamp 1667941163
transform 1 0 36432 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1667941163
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1667941163
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1667941163
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1667941163
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1667941163
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1667941163
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1667941163
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1667941163
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1667941163
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1667941163
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1667941163
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1667941163
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1667941163
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1667941163
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1667941163
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1667941163
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1667941163
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1667941163
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1667941163
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1667941163
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1667941163
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1667941163
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1667941163
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1667941163
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1667941163
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1667941163
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1667941163
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1667941163
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1667941163
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1667941163
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1667941163
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1667941163
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_385
timestamp 1667941163
transform 1 0 36524 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1667941163
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1667941163
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_39
timestamp 1667941163
transform 1 0 4692 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_48
timestamp 1667941163
transform 1 0 5520 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1667941163
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1667941163
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1667941163
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1667941163
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1667941163
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1667941163
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1667941163
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1667941163
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1667941163
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1667941163
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1667941163
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1667941163
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1667941163
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1667941163
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1667941163
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1667941163
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1667941163
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1667941163
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1667941163
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1667941163
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1667941163
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1667941163
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1667941163
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1667941163
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1667941163
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_375
timestamp 1667941163
transform 1 0 35604 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_382
timestamp 1667941163
transform 1 0 36248 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1667941163
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1667941163
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1667941163
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1667941163
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1667941163
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1667941163
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1667941163
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1667941163
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1667941163
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1667941163
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1667941163
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1667941163
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1667941163
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1667941163
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1667941163
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1667941163
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1667941163
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1667941163
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1667941163
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1667941163
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1667941163
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1667941163
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1667941163
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1667941163
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1667941163
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1667941163
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1667941163
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1667941163
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1667941163
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1667941163
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1667941163
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1667941163
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_381
timestamp 1667941163
transform 1 0 36156 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_384
timestamp 1667941163
transform 1 0 36432 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_9
timestamp 1667941163
transform 1 0 1932 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_21
timestamp 1667941163
transform 1 0 3036 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_33
timestamp 1667941163
transform 1 0 4140 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_45
timestamp 1667941163
transform 1 0 5244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1667941163
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1667941163
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1667941163
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1667941163
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1667941163
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1667941163
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1667941163
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1667941163
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1667941163
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1667941163
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1667941163
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1667941163
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1667941163
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1667941163
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1667941163
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1667941163
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1667941163
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1667941163
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1667941163
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1667941163
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1667941163
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1667941163
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1667941163
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1667941163
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1667941163
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1667941163
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1667941163
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_373
timestamp 1667941163
transform 1 0 35420 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_384
timestamp 1667941163
transform 1 0 36432 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1667941163
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1667941163
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1667941163
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1667941163
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1667941163
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1667941163
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1667941163
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1667941163
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1667941163
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1667941163
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1667941163
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1667941163
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1667941163
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1667941163
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1667941163
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1667941163
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1667941163
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1667941163
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1667941163
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1667941163
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1667941163
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1667941163
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1667941163
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1667941163
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1667941163
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1667941163
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1667941163
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1667941163
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1667941163
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1667941163
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1667941163
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_385
timestamp 1667941163
transform 1 0 36524 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1667941163
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1667941163
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1667941163
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1667941163
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1667941163
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1667941163
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1667941163
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1667941163
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1667941163
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1667941163
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1667941163
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1667941163
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1667941163
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1667941163
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1667941163
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1667941163
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1667941163
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1667941163
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1667941163
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1667941163
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1667941163
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1667941163
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1667941163
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1667941163
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1667941163
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1667941163
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1667941163
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1667941163
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1667941163
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1667941163
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1667941163
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1667941163
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_373
timestamp 1667941163
transform 1 0 35420 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_377
timestamp 1667941163
transform 1 0 35788 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_384
timestamp 1667941163
transform 1 0 36432 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1667941163
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1667941163
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1667941163
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1667941163
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1667941163
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1667941163
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1667941163
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1667941163
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1667941163
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1667941163
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1667941163
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1667941163
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1667941163
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1667941163
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1667941163
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1667941163
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1667941163
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1667941163
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1667941163
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1667941163
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1667941163
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1667941163
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1667941163
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1667941163
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1667941163
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1667941163
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1667941163
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1667941163
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1667941163
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1667941163
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1667941163
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1667941163
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_377
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_385
timestamp 1667941163
transform 1 0 36524 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_9
timestamp 1667941163
transform 1 0 1932 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_21
timestamp 1667941163
transform 1 0 3036 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_33
timestamp 1667941163
transform 1 0 4140 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_45
timestamp 1667941163
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1667941163
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1667941163
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1667941163
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1667941163
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1667941163
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1667941163
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1667941163
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1667941163
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1667941163
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1667941163
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1667941163
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1667941163
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1667941163
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1667941163
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1667941163
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1667941163
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1667941163
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1667941163
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1667941163
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1667941163
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1667941163
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1667941163
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1667941163
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1667941163
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1667941163
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1667941163
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1667941163
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1667941163
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_385
timestamp 1667941163
transform 1 0 36524 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_10
timestamp 1667941163
transform 1 0 2024 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_22
timestamp 1667941163
transform 1 0 3128 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1667941163
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1667941163
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1667941163
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1667941163
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1667941163
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1667941163
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1667941163
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1667941163
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1667941163
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1667941163
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1667941163
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1667941163
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1667941163
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1667941163
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1667941163
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1667941163
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1667941163
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1667941163
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1667941163
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1667941163
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1667941163
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1667941163
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1667941163
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1667941163
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1667941163
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1667941163
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1667941163
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1667941163
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1667941163
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1667941163
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_385
timestamp 1667941163
transform 1 0 36524 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_7
timestamp 1667941163
transform 1 0 1748 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_19
timestamp 1667941163
transform 1 0 2852 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_31
timestamp 1667941163
transform 1 0 3956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_43
timestamp 1667941163
transform 1 0 5060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1667941163
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1667941163
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1667941163
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1667941163
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1667941163
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_125
timestamp 1667941163
transform 1 0 12604 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_134
timestamp 1667941163
transform 1 0 13432 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_140
timestamp 1667941163
transform 1 0 13984 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_152
timestamp 1667941163
transform 1 0 15088 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1667941163
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1667941163
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1667941163
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1667941163
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1667941163
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1667941163
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1667941163
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1667941163
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1667941163
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1667941163
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1667941163
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1667941163
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1667941163
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1667941163
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1667941163
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1667941163
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_373
timestamp 1667941163
transform 1 0 35420 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_379
timestamp 1667941163
transform 1 0 35972 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_384
timestamp 1667941163
transform 1 0 36432 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_9
timestamp 1667941163
transform 1 0 1932 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_21
timestamp 1667941163
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1667941163
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1667941163
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1667941163
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1667941163
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1667941163
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1667941163
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1667941163
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1667941163
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1667941163
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1667941163
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1667941163
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1667941163
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1667941163
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1667941163
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1667941163
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1667941163
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1667941163
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1667941163
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1667941163
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1667941163
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1667941163
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_257
timestamp 1667941163
transform 1 0 24748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_261
timestamp 1667941163
transform 1 0 25116 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_267
timestamp 1667941163
transform 1 0 25668 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_279
timestamp 1667941163
transform 1 0 26772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_291
timestamp 1667941163
transform 1 0 27876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_303
timestamp 1667941163
transform 1 0 28980 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1667941163
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_321
timestamp 1667941163
transform 1 0 30636 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_330
timestamp 1667941163
transform 1 0 31464 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_342
timestamp 1667941163
transform 1 0 32568 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_354
timestamp 1667941163
transform 1 0 33672 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_362
timestamp 1667941163
transform 1 0 34408 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_377
timestamp 1667941163
transform 1 0 35788 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_385
timestamp 1667941163
transform 1 0 36524 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1667941163
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1667941163
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1667941163
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1667941163
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1667941163
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1667941163
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1667941163
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1667941163
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1667941163
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1667941163
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1667941163
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1667941163
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1667941163
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1667941163
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1667941163
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1667941163
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1667941163
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1667941163
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1667941163
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1667941163
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1667941163
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1667941163
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1667941163
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1667941163
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1667941163
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1667941163
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1667941163
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1667941163
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1667941163
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1667941163
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1667941163
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1667941163
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_385
timestamp 1667941163
transform 1 0 36524 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1667941163
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1667941163
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1667941163
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1667941163
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1667941163
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1667941163
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1667941163
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1667941163
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1667941163
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1667941163
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1667941163
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1667941163
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1667941163
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1667941163
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1667941163
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1667941163
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1667941163
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1667941163
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1667941163
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1667941163
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1667941163
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1667941163
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1667941163
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1667941163
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1667941163
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1667941163
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1667941163
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1667941163
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1667941163
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1667941163
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1667941163
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1667941163
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_381
timestamp 1667941163
transform 1 0 36156 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_384
timestamp 1667941163
transform 1 0 36432 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_9
timestamp 1667941163
transform 1 0 1932 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_21
timestamp 1667941163
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_33
timestamp 1667941163
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1667941163
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1667941163
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1667941163
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1667941163
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1667941163
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1667941163
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1667941163
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_125
timestamp 1667941163
transform 1 0 12604 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_133
timestamp 1667941163
transform 1 0 13340 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_139
timestamp 1667941163
transform 1 0 13892 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_145
timestamp 1667941163
transform 1 0 14444 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_157
timestamp 1667941163
transform 1 0 15548 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_165
timestamp 1667941163
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1667941163
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1667941163
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1667941163
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1667941163
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1667941163
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1667941163
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1667941163
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_261
timestamp 1667941163
transform 1 0 25116 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_267
timestamp 1667941163
transform 1 0 25668 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1667941163
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1667941163
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1667941163
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1667941163
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1667941163
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1667941163
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1667941163
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1667941163
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_373
timestamp 1667941163
transform 1 0 35420 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_384
timestamp 1667941163
transform 1 0 36432 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1667941163
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1667941163
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1667941163
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1667941163
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1667941163
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1667941163
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1667941163
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1667941163
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1667941163
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1667941163
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1667941163
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1667941163
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1667941163
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1667941163
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1667941163
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1667941163
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1667941163
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1667941163
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1667941163
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1667941163
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1667941163
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1667941163
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1667941163
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1667941163
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1667941163
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1667941163
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1667941163
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1667941163
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1667941163
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1667941163
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1667941163
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1667941163
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_385
timestamp 1667941163
transform 1 0 36524 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1667941163
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1667941163
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1667941163
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1667941163
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1667941163
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1667941163
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1667941163
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1667941163
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1667941163
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1667941163
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1667941163
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1667941163
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1667941163
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1667941163
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1667941163
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1667941163
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1667941163
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1667941163
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1667941163
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1667941163
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1667941163
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1667941163
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1667941163
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1667941163
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1667941163
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_286
timestamp 1667941163
transform 1 0 27416 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_292
timestamp 1667941163
transform 1 0 27968 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_304
timestamp 1667941163
transform 1 0 29072 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_316
timestamp 1667941163
transform 1 0 30176 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_328
timestamp 1667941163
transform 1 0 31280 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1667941163
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1667941163
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_373
timestamp 1667941163
transform 1 0 35420 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_379
timestamp 1667941163
transform 1 0 35972 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_384
timestamp 1667941163
transform 1 0 36432 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_7
timestamp 1667941163
transform 1 0 1748 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_19
timestamp 1667941163
transform 1 0 2852 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1667941163
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1667941163
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1667941163
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1667941163
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1667941163
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1667941163
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1667941163
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1667941163
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1667941163
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1667941163
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1667941163
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1667941163
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1667941163
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1667941163
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1667941163
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1667941163
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1667941163
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1667941163
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1667941163
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1667941163
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1667941163
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1667941163
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1667941163
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1667941163
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1667941163
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1667941163
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1667941163
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1667941163
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1667941163
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1667941163
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1667941163
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_385
timestamp 1667941163
transform 1 0 36524 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_9
timestamp 1667941163
transform 1 0 1932 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_21
timestamp 1667941163
transform 1 0 3036 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_33
timestamp 1667941163
transform 1 0 4140 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_45
timestamp 1667941163
transform 1 0 5244 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp 1667941163
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1667941163
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1667941163
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1667941163
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1667941163
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1667941163
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1667941163
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1667941163
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1667941163
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1667941163
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1667941163
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1667941163
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1667941163
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1667941163
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1667941163
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1667941163
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1667941163
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1667941163
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1667941163
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1667941163
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1667941163
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1667941163
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1667941163
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1667941163
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1667941163
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1667941163
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1667941163
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1667941163
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_385
timestamp 1667941163
transform 1 0 36524 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_10
timestamp 1667941163
transform 1 0 2024 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_16
timestamp 1667941163
transform 1 0 2576 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1667941163
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1667941163
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_65
timestamp 1667941163
transform 1 0 7084 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1667941163
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1667941163
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1667941163
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1667941163
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1667941163
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1667941163
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1667941163
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1667941163
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_165
timestamp 1667941163
transform 1 0 16284 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_175
timestamp 1667941163
transform 1 0 17204 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_181
timestamp 1667941163
transform 1 0 17756 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_193
timestamp 1667941163
transform 1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1667941163
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1667941163
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1667941163
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1667941163
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1667941163
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1667941163
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1667941163
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1667941163
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1667941163
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1667941163
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1667941163
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1667941163
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1667941163
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1667941163
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1667941163
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_377
timestamp 1667941163
transform 1 0 35788 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_385
timestamp 1667941163
transform 1 0 36524 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1667941163
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1667941163
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1667941163
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1667941163
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1667941163
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1667941163
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1667941163
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1667941163
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1667941163
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1667941163
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1667941163
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1667941163
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1667941163
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1667941163
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1667941163
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1667941163
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1667941163
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1667941163
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1667941163
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1667941163
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1667941163
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1667941163
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1667941163
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1667941163
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1667941163
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1667941163
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1667941163
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1667941163
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1667941163
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1667941163
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1667941163
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1667941163
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_385
timestamp 1667941163
transform 1 0 36524 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_9
timestamp 1667941163
transform 1 0 1932 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_16
timestamp 1667941163
transform 1 0 2576 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_22
timestamp 1667941163
transform 1 0 3128 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1667941163
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1667941163
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_65
timestamp 1667941163
transform 1 0 7084 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_72
timestamp 1667941163
transform 1 0 7728 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_78
timestamp 1667941163
transform 1 0 8280 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_90
timestamp 1667941163
transform 1 0 9384 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_96
timestamp 1667941163
transform 1 0 9936 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_108
timestamp 1667941163
transform 1 0 11040 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_120
timestamp 1667941163
transform 1 0 12144 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_132
timestamp 1667941163
transform 1 0 13248 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1667941163
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1667941163
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1667941163
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1667941163
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1667941163
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_209
timestamp 1667941163
transform 1 0 20332 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_217
timestamp 1667941163
transform 1 0 21068 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_221
timestamp 1667941163
transform 1 0 21436 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_227
timestamp 1667941163
transform 1 0 21988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_239
timestamp 1667941163
transform 1 0 23092 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1667941163
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1667941163
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1667941163
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1667941163
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1667941163
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1667941163
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1667941163
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1667941163
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1667941163
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1667941163
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1667941163
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_377
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_385
timestamp 1667941163
transform 1 0 36524 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1667941163
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1667941163
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1667941163
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1667941163
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1667941163
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1667941163
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1667941163
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1667941163
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1667941163
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1667941163
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1667941163
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_137
timestamp 1667941163
transform 1 0 13708 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_146
timestamp 1667941163
transform 1 0 14536 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_152
timestamp 1667941163
transform 1 0 15088 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_156
timestamp 1667941163
transform 1 0 15456 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_160
timestamp 1667941163
transform 1 0 15824 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1667941163
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1667941163
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1667941163
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1667941163
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1667941163
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1667941163
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1667941163
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1667941163
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1667941163
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1667941163
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1667941163
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1667941163
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1667941163
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1667941163
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1667941163
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1667941163
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1667941163
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1667941163
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_385
timestamp 1667941163
transform 1 0 36524 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1667941163
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1667941163
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1667941163
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1667941163
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1667941163
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1667941163
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1667941163
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1667941163
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_109
timestamp 1667941163
transform 1 0 11132 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_117
timestamp 1667941163
transform 1 0 11868 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_121
timestamp 1667941163
transform 1 0 12236 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_131
timestamp 1667941163
transform 1 0 13156 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_135
timestamp 1667941163
transform 1 0 13524 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1667941163
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_156
timestamp 1667941163
transform 1 0 15456 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_168
timestamp 1667941163
transform 1 0 16560 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_180
timestamp 1667941163
transform 1 0 17664 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_192
timestamp 1667941163
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1667941163
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1667941163
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1667941163
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1667941163
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1667941163
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1667941163
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1667941163
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1667941163
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1667941163
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1667941163
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_317
timestamp 1667941163
transform 1 0 30268 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_322
timestamp 1667941163
transform 1 0 30728 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_328
timestamp 1667941163
transform 1 0 31280 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_340
timestamp 1667941163
transform 1 0 32384 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_352
timestamp 1667941163
transform 1 0 33488 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_371
timestamp 1667941163
transform 1 0 35236 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_374
timestamp 1667941163
transform 1 0 35512 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_381
timestamp 1667941163
transform 1 0 36156 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_385
timestamp 1667941163
transform 1 0 36524 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_9
timestamp 1667941163
transform 1 0 1932 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_21
timestamp 1667941163
transform 1 0 3036 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_33
timestamp 1667941163
transform 1 0 4140 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_45
timestamp 1667941163
transform 1 0 5244 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1667941163
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_65
timestamp 1667941163
transform 1 0 7084 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_77
timestamp 1667941163
transform 1 0 8188 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_89
timestamp 1667941163
transform 1 0 9292 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_101
timestamp 1667941163
transform 1 0 10396 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_109
timestamp 1667941163
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_121
timestamp 1667941163
transform 1 0 12236 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_127
timestamp 1667941163
transform 1 0 12788 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_134
timestamp 1667941163
transform 1 0 13432 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_141
timestamp 1667941163
transform 1 0 14076 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_148
timestamp 1667941163
transform 1 0 14720 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1667941163
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1667941163
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1667941163
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1667941163
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1667941163
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1667941163
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1667941163
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1667941163
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1667941163
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1667941163
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1667941163
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1667941163
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1667941163
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1667941163
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1667941163
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1667941163
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1667941163
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1667941163
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1667941163
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_373
timestamp 1667941163
transform 1 0 35420 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_379
timestamp 1667941163
transform 1 0 35972 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_384
timestamp 1667941163
transform 1 0 36432 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1667941163
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1667941163
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_41
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_49
timestamp 1667941163
transform 1 0 5612 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_53
timestamp 1667941163
transform 1 0 5980 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_59
timestamp 1667941163
transform 1 0 6532 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_66
timestamp 1667941163
transform 1 0 7176 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_72
timestamp 1667941163
transform 1 0 7728 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1667941163
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_90
timestamp 1667941163
transform 1 0 9384 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_98
timestamp 1667941163
transform 1 0 10120 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_101
timestamp 1667941163
transform 1 0 10396 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_108
timestamp 1667941163
transform 1 0 11040 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_115
timestamp 1667941163
transform 1 0 11684 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_123
timestamp 1667941163
transform 1 0 12420 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_127
timestamp 1667941163
transform 1 0 12788 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1667941163
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_145
timestamp 1667941163
transform 1 0 14444 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_158
timestamp 1667941163
transform 1 0 15640 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_165
timestamp 1667941163
transform 1 0 16284 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_171
timestamp 1667941163
transform 1 0 16836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_183
timestamp 1667941163
transform 1 0 17940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1667941163
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1667941163
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1667941163
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1667941163
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1667941163
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1667941163
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1667941163
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1667941163
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1667941163
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1667941163
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1667941163
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1667941163
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_336
timestamp 1667941163
transform 1 0 32016 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_342
timestamp 1667941163
transform 1 0 32568 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_354
timestamp 1667941163
transform 1 0 33672 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_362
timestamp 1667941163
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_377
timestamp 1667941163
transform 1 0 35788 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_385
timestamp 1667941163
transform 1 0 36524 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_12
timestamp 1667941163
transform 1 0 2208 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_18
timestamp 1667941163
transform 1 0 2760 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_30
timestamp 1667941163
transform 1 0 3864 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_42
timestamp 1667941163
transform 1 0 4968 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1667941163
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_69
timestamp 1667941163
transform 1 0 7452 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_80
timestamp 1667941163
transform 1 0 8464 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_93
timestamp 1667941163
transform 1 0 9660 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1667941163
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_117
timestamp 1667941163
transform 1 0 11868 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_124
timestamp 1667941163
transform 1 0 12512 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_131
timestamp 1667941163
transform 1 0 13156 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_143
timestamp 1667941163
transform 1 0 14260 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_156
timestamp 1667941163
transform 1 0 15456 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_163
timestamp 1667941163
transform 1 0 16100 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1667941163
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_173
timestamp 1667941163
transform 1 0 17020 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_185
timestamp 1667941163
transform 1 0 18124 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_197
timestamp 1667941163
transform 1 0 19228 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_209
timestamp 1667941163
transform 1 0 20332 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_221
timestamp 1667941163
transform 1 0 21436 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1667941163
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1667941163
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1667941163
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1667941163
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1667941163
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1667941163
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1667941163
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1667941163
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1667941163
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1667941163
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1667941163
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_373
timestamp 1667941163
transform 1 0 35420 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_379
timestamp 1667941163
transform 1 0 35972 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_384
timestamp 1667941163
transform 1 0 36432 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1667941163
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1667941163
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_41
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_49
timestamp 1667941163
transform 1 0 5612 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_55
timestamp 1667941163
transform 1 0 6164 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_67
timestamp 1667941163
transform 1 0 7268 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_79
timestamp 1667941163
transform 1 0 8372 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1667941163
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_97
timestamp 1667941163
transform 1 0 10028 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_104
timestamp 1667941163
transform 1 0 10672 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_117
timestamp 1667941163
transform 1 0 11868 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_129
timestamp 1667941163
transform 1 0 12972 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1667941163
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_148
timestamp 1667941163
transform 1 0 14720 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_161
timestamp 1667941163
transform 1 0 15916 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_169
timestamp 1667941163
transform 1 0 16652 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_175
timestamp 1667941163
transform 1 0 17204 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_181
timestamp 1667941163
transform 1 0 17756 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_193
timestamp 1667941163
transform 1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1667941163
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_221
timestamp 1667941163
transform 1 0 21436 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_227
timestamp 1667941163
transform 1 0 21988 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_230
timestamp 1667941163
transform 1 0 22264 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_242
timestamp 1667941163
transform 1 0 23368 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1667941163
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1667941163
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1667941163
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1667941163
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1667941163
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1667941163
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_321
timestamp 1667941163
transform 1 0 30636 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_328
timestamp 1667941163
transform 1 0 31280 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_340
timestamp 1667941163
transform 1 0 32384 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_352
timestamp 1667941163
transform 1 0 33488 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_377
timestamp 1667941163
transform 1 0 35788 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_385
timestamp 1667941163
transform 1 0 36524 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_9
timestamp 1667941163
transform 1 0 1932 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_16
timestamp 1667941163
transform 1 0 2576 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_28
timestamp 1667941163
transform 1 0 3680 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_40
timestamp 1667941163
transform 1 0 4784 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_52
timestamp 1667941163
transform 1 0 5888 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_62
timestamp 1667941163
transform 1 0 6808 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_68
timestamp 1667941163
transform 1 0 7360 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_80
timestamp 1667941163
transform 1 0 8464 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_92
timestamp 1667941163
transform 1 0 9568 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_96
timestamp 1667941163
transform 1 0 9936 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_103
timestamp 1667941163
transform 1 0 10580 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1667941163
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_132
timestamp 1667941163
transform 1 0 13248 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_145
timestamp 1667941163
transform 1 0 14444 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_39_162
timestamp 1667941163
transform 1 0 16008 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_174
timestamp 1667941163
transform 1 0 17112 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_180
timestamp 1667941163
transform 1 0 17664 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_192
timestamp 1667941163
transform 1 0 18768 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_204
timestamp 1667941163
transform 1 0 19872 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_216
timestamp 1667941163
transform 1 0 20976 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_229
timestamp 1667941163
transform 1 0 22172 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_234
timestamp 1667941163
transform 1 0 22632 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_246
timestamp 1667941163
transform 1 0 23736 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_258
timestamp 1667941163
transform 1 0 24840 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_270
timestamp 1667941163
transform 1 0 25944 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1667941163
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1667941163
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1667941163
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1667941163
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1667941163
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1667941163
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1667941163
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_373
timestamp 1667941163
transform 1 0 35420 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_377
timestamp 1667941163
transform 1 0 35788 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_381
timestamp 1667941163
transform 1 0 36156 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_385
timestamp 1667941163
transform 1 0 36524 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1667941163
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1667941163
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1667941163
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1667941163
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_65
timestamp 1667941163
transform 1 0 7084 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1667941163
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_98
timestamp 1667941163
transform 1 0 10120 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_106
timestamp 1667941163
transform 1 0 10856 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_116
timestamp 1667941163
transform 1 0 11776 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_128
timestamp 1667941163
transform 1 0 12880 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_134
timestamp 1667941163
transform 1 0 13432 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1667941163
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_152
timestamp 1667941163
transform 1 0 15088 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_165
timestamp 1667941163
transform 1 0 16284 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_172
timestamp 1667941163
transform 1 0 16928 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_179
timestamp 1667941163
transform 1 0 17572 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_185
timestamp 1667941163
transform 1 0 18124 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_191
timestamp 1667941163
transform 1 0 18676 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1667941163
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1667941163
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1667941163
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1667941163
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1667941163
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1667941163
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1667941163
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1667941163
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_289
timestamp 1667941163
transform 1 0 27692 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_297
timestamp 1667941163
transform 1 0 28428 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_303
timestamp 1667941163
transform 1 0 28980 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1667941163
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1667941163
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1667941163
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1667941163
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1667941163
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1667941163
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_377
timestamp 1667941163
transform 1 0 35788 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_385
timestamp 1667941163
transform 1 0 36524 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1667941163
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1667941163
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1667941163
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1667941163
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1667941163
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_69
timestamp 1667941163
transform 1 0 7452 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_77
timestamp 1667941163
transform 1 0 8188 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_81
timestamp 1667941163
transform 1 0 8556 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_88
timestamp 1667941163
transform 1 0 9200 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_97
timestamp 1667941163
transform 1 0 10028 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1667941163
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_117
timestamp 1667941163
transform 1 0 11868 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_134
timestamp 1667941163
transform 1 0 13432 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_142
timestamp 1667941163
transform 1 0 14168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_146
timestamp 1667941163
transform 1 0 14536 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_153
timestamp 1667941163
transform 1 0 15180 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1667941163
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_180
timestamp 1667941163
transform 1 0 17664 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_189
timestamp 1667941163
transform 1 0 18492 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_195
timestamp 1667941163
transform 1 0 19044 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_201
timestamp 1667941163
transform 1 0 19596 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_213
timestamp 1667941163
transform 1 0 20700 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_221
timestamp 1667941163
transform 1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1667941163
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1667941163
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_261
timestamp 1667941163
transform 1 0 25116 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_272
timestamp 1667941163
transform 1 0 26128 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1667941163
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1667941163
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1667941163
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1667941163
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1667941163
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1667941163
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_354
timestamp 1667941163
transform 1 0 33672 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_366
timestamp 1667941163
transform 1 0 34776 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_376
timestamp 1667941163
transform 1 0 35696 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_384
timestamp 1667941163
transform 1 0 36432 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_8
timestamp 1667941163
transform 1 0 1840 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_14
timestamp 1667941163
transform 1 0 2392 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_26
timestamp 1667941163
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1667941163
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1667941163
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1667941163
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1667941163
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_96
timestamp 1667941163
transform 1 0 9936 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_103
timestamp 1667941163
transform 1 0 10580 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_110
timestamp 1667941163
transform 1 0 11224 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_123
timestamp 1667941163
transform 1 0 12420 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_136
timestamp 1667941163
transform 1 0 13616 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_148
timestamp 1667941163
transform 1 0 14720 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_161
timestamp 1667941163
transform 1 0 15916 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_174
timestamp 1667941163
transform 1 0 17112 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_181
timestamp 1667941163
transform 1 0 17756 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_188
timestamp 1667941163
transform 1 0 18400 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1667941163
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_201
timestamp 1667941163
transform 1 0 19596 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_213
timestamp 1667941163
transform 1 0 20700 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_225
timestamp 1667941163
transform 1 0 21804 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_237
timestamp 1667941163
transform 1 0 22908 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_249
timestamp 1667941163
transform 1 0 24012 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1667941163
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1667941163
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1667941163
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1667941163
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1667941163
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1667941163
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1667941163
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1667941163
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1667941163
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1667941163
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_385
timestamp 1667941163
transform 1 0 36524 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1667941163
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1667941163
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1667941163
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1667941163
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1667941163
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1667941163
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_81
timestamp 1667941163
transform 1 0 8556 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_89
timestamp 1667941163
transform 1 0 9292 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_95
timestamp 1667941163
transform 1 0 9844 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_102
timestamp 1667941163
transform 1 0 10488 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1667941163
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_132
timestamp 1667941163
transform 1 0 13248 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_138
timestamp 1667941163
transform 1 0 13800 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_148
timestamp 1667941163
transform 1 0 14720 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1667941163
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1667941163
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_173
timestamp 1667941163
transform 1 0 17020 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_177
timestamp 1667941163
transform 1 0 17388 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_184
timestamp 1667941163
transform 1 0 18032 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_191
timestamp 1667941163
transform 1 0 18676 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_197
timestamp 1667941163
transform 1 0 19228 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_203
timestamp 1667941163
transform 1 0 19780 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_209
timestamp 1667941163
transform 1 0 20332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_221
timestamp 1667941163
transform 1 0 21436 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1667941163
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1667941163
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1667941163
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1667941163
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1667941163
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1667941163
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1667941163
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1667941163
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1667941163
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1667941163
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1667941163
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1667941163
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_385
timestamp 1667941163
transform 1 0 36524 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_7
timestamp 1667941163
transform 1 0 1748 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_13
timestamp 1667941163
transform 1 0 2300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_25
timestamp 1667941163
transform 1 0 3404 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_53
timestamp 1667941163
transform 1 0 5980 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_58
timestamp 1667941163
transform 1 0 6440 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_64
timestamp 1667941163
transform 1 0 6992 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_74
timestamp 1667941163
transform 1 0 7912 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_81
timestamp 1667941163
transform 1 0 8556 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_91
timestamp 1667941163
transform 1 0 9476 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_95
timestamp 1667941163
transform 1 0 9844 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_103
timestamp 1667941163
transform 1 0 10580 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_107
timestamp 1667941163
transform 1 0 10948 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_120
timestamp 1667941163
transform 1 0 12144 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_128
timestamp 1667941163
transform 1 0 12880 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1667941163
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_146
timestamp 1667941163
transform 1 0 14536 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_159
timestamp 1667941163
transform 1 0 15732 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_170
timestamp 1667941163
transform 1 0 16744 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_183
timestamp 1667941163
transform 1 0 17940 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_190
timestamp 1667941163
transform 1 0 18584 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_201
timestamp 1667941163
transform 1 0 19596 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_207
timestamp 1667941163
transform 1 0 20148 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_219
timestamp 1667941163
transform 1 0 21252 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_231
timestamp 1667941163
transform 1 0 22356 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_243
timestamp 1667941163
transform 1 0 23460 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1667941163
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1667941163
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1667941163
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1667941163
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1667941163
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1667941163
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1667941163
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1667941163
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1667941163
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1667941163
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1667941163
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_377
timestamp 1667941163
transform 1 0 35788 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_385
timestamp 1667941163
transform 1 0 36524 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_9
timestamp 1667941163
transform 1 0 1932 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_16
timestamp 1667941163
transform 1 0 2576 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_28
timestamp 1667941163
transform 1 0 3680 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_31
timestamp 1667941163
transform 1 0 3956 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_37
timestamp 1667941163
transform 1 0 4508 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_49
timestamp 1667941163
transform 1 0 5612 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1667941163
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_65
timestamp 1667941163
transform 1 0 7084 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_75
timestamp 1667941163
transform 1 0 8004 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_79
timestamp 1667941163
transform 1 0 8372 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_82
timestamp 1667941163
transform 1 0 8648 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_89
timestamp 1667941163
transform 1 0 9292 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_96
timestamp 1667941163
transform 1 0 9936 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_103
timestamp 1667941163
transform 1 0 10580 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_109
timestamp 1667941163
transform 1 0 11132 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_117
timestamp 1667941163
transform 1 0 11868 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_121
timestamp 1667941163
transform 1 0 12236 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_134
timestamp 1667941163
transform 1 0 13432 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_147
timestamp 1667941163
transform 1 0 14628 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_153
timestamp 1667941163
transform 1 0 15180 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1667941163
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_186
timestamp 1667941163
transform 1 0 18216 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_193
timestamp 1667941163
transform 1 0 18860 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_199
timestamp 1667941163
transform 1 0 19412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_211
timestamp 1667941163
transform 1 0 20516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1667941163
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1667941163
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1667941163
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1667941163
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1667941163
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1667941163
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1667941163
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1667941163
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1667941163
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1667941163
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1667941163
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1667941163
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1667941163
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_373
timestamp 1667941163
transform 1 0 35420 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_377
timestamp 1667941163
transform 1 0 35788 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_384
timestamp 1667941163
transform 1 0 36432 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_7
timestamp 1667941163
transform 1 0 1748 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_13
timestamp 1667941163
transform 1 0 2300 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_17
timestamp 1667941163
transform 1 0 2668 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_24
timestamp 1667941163
transform 1 0 3312 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_33
timestamp 1667941163
transform 1 0 4140 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_39
timestamp 1667941163
transform 1 0 4692 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_45
timestamp 1667941163
transform 1 0 5244 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_51
timestamp 1667941163
transform 1 0 5796 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_54
timestamp 1667941163
transform 1 0 6072 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_58
timestamp 1667941163
transform 1 0 6440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_62
timestamp 1667941163
transform 1 0 6808 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_69
timestamp 1667941163
transform 1 0 7452 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_82
timestamp 1667941163
transform 1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_91
timestamp 1667941163
transform 1 0 9476 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_101
timestamp 1667941163
transform 1 0 10396 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_110
timestamp 1667941163
transform 1 0 11224 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_117
timestamp 1667941163
transform 1 0 11868 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_124
timestamp 1667941163
transform 1 0 12512 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_137
timestamp 1667941163
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_145
timestamp 1667941163
transform 1 0 14444 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_152
timestamp 1667941163
transform 1 0 15088 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_165
timestamp 1667941163
transform 1 0 16284 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_178
timestamp 1667941163
transform 1 0 17480 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_185
timestamp 1667941163
transform 1 0 18124 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1667941163
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_201
timestamp 1667941163
transform 1 0 19596 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_213
timestamp 1667941163
transform 1 0 20700 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_225
timestamp 1667941163
transform 1 0 21804 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_237
timestamp 1667941163
transform 1 0 22908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_249
timestamp 1667941163
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1667941163
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_277
timestamp 1667941163
transform 1 0 26588 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_281
timestamp 1667941163
transform 1 0 26956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_285
timestamp 1667941163
transform 1 0 27324 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_297
timestamp 1667941163
transform 1 0 28428 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_305
timestamp 1667941163
transform 1 0 29164 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1667941163
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1667941163
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1667941163
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1667941163
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1667941163
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_381
timestamp 1667941163
transform 1 0 36156 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_384
timestamp 1667941163
transform 1 0 36432 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_8
timestamp 1667941163
transform 1 0 1840 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_15
timestamp 1667941163
transform 1 0 2484 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_22
timestamp 1667941163
transform 1 0 3128 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_28
timestamp 1667941163
transform 1 0 3680 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_34
timestamp 1667941163
transform 1 0 4232 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_42
timestamp 1667941163
transform 1 0 4968 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_48
timestamp 1667941163
transform 1 0 5520 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_54
timestamp 1667941163
transform 1 0 6072 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_62
timestamp 1667941163
transform 1 0 6808 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_69
timestamp 1667941163
transform 1 0 7452 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_76
timestamp 1667941163
transform 1 0 8096 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_85
timestamp 1667941163
transform 1 0 8924 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_98
timestamp 1667941163
transform 1 0 10120 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_106
timestamp 1667941163
transform 1 0 10856 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_110
timestamp 1667941163
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_117
timestamp 1667941163
transform 1 0 11868 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_124
timestamp 1667941163
transform 1 0 12512 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_137
timestamp 1667941163
transform 1 0 13708 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_143
timestamp 1667941163
transform 1 0 14260 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_153
timestamp 1667941163
transform 1 0 15180 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_166
timestamp 1667941163
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_178
timestamp 1667941163
transform 1 0 17480 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_185
timestamp 1667941163
transform 1 0 18124 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_192
timestamp 1667941163
transform 1 0 18768 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_198
timestamp 1667941163
transform 1 0 19320 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_204
timestamp 1667941163
transform 1 0 19872 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_216
timestamp 1667941163
transform 1 0 20976 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1667941163
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1667941163
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1667941163
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1667941163
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1667941163
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1667941163
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1667941163
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1667941163
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1667941163
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1667941163
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1667941163
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1667941163
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_373
timestamp 1667941163
transform 1 0 35420 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_384
timestamp 1667941163
transform 1 0 36432 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_8
timestamp 1667941163
transform 1 0 1840 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_15
timestamp 1667941163
transform 1 0 2484 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_22
timestamp 1667941163
transform 1 0 3128 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_34
timestamp 1667941163
transform 1 0 4232 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_38
timestamp 1667941163
transform 1 0 4600 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_41
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_47
timestamp 1667941163
transform 1 0 5428 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_53
timestamp 1667941163
transform 1 0 5980 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1667941163
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1667941163
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_92
timestamp 1667941163
transform 1 0 9568 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_99
timestamp 1667941163
transform 1 0 10212 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_112
timestamp 1667941163
transform 1 0 11408 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_125
timestamp 1667941163
transform 1 0 12604 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_138
timestamp 1667941163
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_146
timestamp 1667941163
transform 1 0 14536 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_159
timestamp 1667941163
transform 1 0 15732 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_163
timestamp 1667941163
transform 1 0 16100 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_173
timestamp 1667941163
transform 1 0 17020 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_180
timestamp 1667941163
transform 1 0 17664 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_187
timestamp 1667941163
transform 1 0 18308 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_48_193
timestamp 1667941163
transform 1 0 18860 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1667941163
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1667941163
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1667941163
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1667941163
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1667941163
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1667941163
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1667941163
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1667941163
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1667941163
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1667941163
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_320
timestamp 1667941163
transform 1 0 30544 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_332
timestamp 1667941163
transform 1 0 31648 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_344
timestamp 1667941163
transform 1 0 32752 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_356
timestamp 1667941163
transform 1 0 33856 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_377
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_385
timestamp 1667941163
transform 1 0 36524 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_15
timestamp 1667941163
transform 1 0 2484 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_19
timestamp 1667941163
transform 1 0 2852 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_40
timestamp 1667941163
transform 1 0 4784 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_48
timestamp 1667941163
transform 1 0 5520 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_54
timestamp 1667941163
transform 1 0 6072 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_79
timestamp 1667941163
transform 1 0 8372 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_86
timestamp 1667941163
transform 1 0 9016 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_93
timestamp 1667941163
transform 1 0 9660 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_106
timestamp 1667941163
transform 1 0 10856 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_130
timestamp 1667941163
transform 1 0 13064 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_147
timestamp 1667941163
transform 1 0 14628 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_164
timestamp 1667941163
transform 1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_180
timestamp 1667941163
transform 1 0 17664 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_187
timestamp 1667941163
transform 1 0 18308 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1667941163
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1667941163
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1667941163
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1667941163
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1667941163
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1667941163
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1667941163
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1667941163
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1667941163
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1667941163
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1667941163
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1667941163
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1667941163
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1667941163
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_385
timestamp 1667941163
transform 1 0 36524 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_8
timestamp 1667941163
transform 1 0 1840 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_15
timestamp 1667941163
transform 1 0 2484 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_22
timestamp 1667941163
transform 1 0 3128 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_34
timestamp 1667941163
transform 1 0 4232 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_41
timestamp 1667941163
transform 1 0 4876 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_47
timestamp 1667941163
transform 1 0 5428 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_54
timestamp 1667941163
transform 1 0 6072 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_82
timestamp 1667941163
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_107
timestamp 1667941163
transform 1 0 10948 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_124
timestamp 1667941163
transform 1 0 12512 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_50_137
timestamp 1667941163
transform 1 0 13708 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_152
timestamp 1667941163
transform 1 0 15088 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_169
timestamp 1667941163
transform 1 0 16652 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_176
timestamp 1667941163
transform 1 0 17296 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_188
timestamp 1667941163
transform 1 0 18400 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1667941163
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1667941163
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1667941163
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1667941163
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1667941163
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1667941163
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1667941163
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1667941163
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1667941163
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1667941163
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1667941163
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1667941163
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1667941163
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1667941163
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1667941163
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_377
timestamp 1667941163
transform 1 0 35788 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_381
timestamp 1667941163
transform 1 0 36156 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_384
timestamp 1667941163
transform 1 0 36432 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_26
timestamp 1667941163
transform 1 0 3496 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_54
timestamp 1667941163
transform 1 0 6072 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_62
timestamp 1667941163
transform 1 0 6808 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_70
timestamp 1667941163
transform 1 0 7544 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_92
timestamp 1667941163
transform 1 0 9568 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_103
timestamp 1667941163
transform 1 0 10580 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1667941163
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_117
timestamp 1667941163
transform 1 0 11868 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_121
timestamp 1667941163
transform 1 0 12236 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_128
timestamp 1667941163
transform 1 0 12880 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_132
timestamp 1667941163
transform 1 0 13248 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_136
timestamp 1667941163
transform 1 0 13616 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_143
timestamp 1667941163
transform 1 0 14260 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_150
timestamp 1667941163
transform 1 0 14904 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_163
timestamp 1667941163
transform 1 0 16100 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1667941163
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_173
timestamp 1667941163
transform 1 0 17020 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_185
timestamp 1667941163
transform 1 0 18124 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_197
timestamp 1667941163
transform 1 0 19228 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_209
timestamp 1667941163
transform 1 0 20332 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_221
timestamp 1667941163
transform 1 0 21436 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1667941163
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1667941163
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1667941163
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1667941163
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1667941163
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1667941163
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1667941163
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1667941163
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1667941163
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1667941163
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1667941163
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_373
timestamp 1667941163
transform 1 0 35420 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_384
timestamp 1667941163
transform 1 0 36432 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_9
timestamp 1667941163
transform 1 0 1932 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_16
timestamp 1667941163
transform 1 0 2576 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_23
timestamp 1667941163
transform 1 0 3220 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1667941163
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_52
timestamp 1667941163
transform 1 0 5888 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_60
timestamp 1667941163
transform 1 0 6624 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_82
timestamp 1667941163
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_107
timestamp 1667941163
transform 1 0 10948 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_128
timestamp 1667941163
transform 1 0 12880 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_135
timestamp 1667941163
transform 1 0 13524 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1667941163
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_152
timestamp 1667941163
transform 1 0 15088 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_159
timestamp 1667941163
transform 1 0 15732 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1667941163
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1667941163
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1667941163
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1667941163
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1667941163
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1667941163
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1667941163
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1667941163
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1667941163
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1667941163
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1667941163
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1667941163
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1667941163
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1667941163
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1667941163
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1667941163
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1667941163
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1667941163
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1667941163
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_377
timestamp 1667941163
transform 1 0 35788 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_385
timestamp 1667941163
transform 1 0 36524 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_29
timestamp 1667941163
transform 1 0 3772 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_54
timestamp 1667941163
transform 1 0 6072 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_62
timestamp 1667941163
transform 1 0 6808 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_69
timestamp 1667941163
transform 1 0 7452 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_76
timestamp 1667941163
transform 1 0 8096 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_101
timestamp 1667941163
transform 1 0 10396 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_108
timestamp 1667941163
transform 1 0 11040 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_128
timestamp 1667941163
transform 1 0 12880 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_145
timestamp 1667941163
transform 1 0 14444 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_158
timestamp 1667941163
transform 1 0 15640 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 1667941163
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1667941163
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1667941163
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1667941163
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1667941163
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1667941163
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1667941163
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1667941163
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1667941163
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1667941163
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1667941163
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1667941163
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1667941163
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1667941163
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1667941163
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1667941163
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1667941163
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1667941163
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_385
timestamp 1667941163
transform 1 0 36524 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_15
timestamp 1667941163
transform 1 0 2484 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_22
timestamp 1667941163
transform 1 0 3128 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_34
timestamp 1667941163
transform 1 0 4232 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_41
timestamp 1667941163
transform 1 0 4876 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_48
timestamp 1667941163
transform 1 0 5520 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_55
timestamp 1667941163
transform 1 0 6164 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_82
timestamp 1667941163
transform 1 0 8648 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_89
timestamp 1667941163
transform 1 0 9292 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_54_98
timestamp 1667941163
transform 1 0 10120 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_104
timestamp 1667941163
transform 1 0 10672 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_108
timestamp 1667941163
transform 1 0 11040 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_115
timestamp 1667941163
transform 1 0 11684 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_122
timestamp 1667941163
transform 1 0 12328 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_126
timestamp 1667941163
transform 1 0 12696 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_130
timestamp 1667941163
transform 1 0 13064 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_54_137
timestamp 1667941163
transform 1 0 13708 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_150
timestamp 1667941163
transform 1 0 14904 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_162
timestamp 1667941163
transform 1 0 16008 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_174
timestamp 1667941163
transform 1 0 17112 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_186
timestamp 1667941163
transform 1 0 18216 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_194
timestamp 1667941163
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1667941163
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1667941163
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_233
timestamp 1667941163
transform 1 0 22540 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_237
timestamp 1667941163
transform 1 0 22908 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_243
timestamp 1667941163
transform 1 0 23460 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1667941163
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1667941163
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1667941163
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1667941163
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1667941163
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1667941163
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1667941163
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1667941163
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1667941163
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1667941163
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_381
timestamp 1667941163
transform 1 0 36156 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_385
timestamp 1667941163
transform 1 0 36524 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_8
timestamp 1667941163
transform 1 0 1840 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_32
timestamp 1667941163
transform 1 0 4048 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_39
timestamp 1667941163
transform 1 0 4692 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_46
timestamp 1667941163
transform 1 0 5336 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_53
timestamp 1667941163
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_62
timestamp 1667941163
transform 1 0 6808 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_69
timestamp 1667941163
transform 1 0 7452 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_75
timestamp 1667941163
transform 1 0 8004 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_99
timestamp 1667941163
transform 1 0 10212 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1667941163
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1667941163
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_119
timestamp 1667941163
transform 1 0 12052 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_123
timestamp 1667941163
transform 1 0 12420 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_130
timestamp 1667941163
transform 1 0 13064 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_143
timestamp 1667941163
transform 1 0 14260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_155
timestamp 1667941163
transform 1 0 15364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1667941163
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1667941163
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1667941163
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1667941163
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1667941163
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1667941163
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1667941163
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1667941163
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1667941163
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1667941163
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1667941163
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1667941163
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1667941163
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1667941163
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1667941163
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1667941163
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1667941163
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_373
timestamp 1667941163
transform 1 0 35420 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_384
timestamp 1667941163
transform 1 0 36432 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_26
timestamp 1667941163
transform 1 0 3496 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_35
timestamp 1667941163
transform 1 0 4324 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_42
timestamp 1667941163
transform 1 0 4968 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_49
timestamp 1667941163
transform 1 0 5612 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_56
timestamp 1667941163
transform 1 0 6256 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_60
timestamp 1667941163
transform 1 0 6624 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_82
timestamp 1667941163
transform 1 0 8648 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_108
timestamp 1667941163
transform 1 0 11040 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_114
timestamp 1667941163
transform 1 0 11592 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_125
timestamp 1667941163
transform 1 0 12604 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_138
timestamp 1667941163
transform 1 0 13800 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_145
timestamp 1667941163
transform 1 0 14444 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_157
timestamp 1667941163
transform 1 0 15548 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_169
timestamp 1667941163
transform 1 0 16652 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_181
timestamp 1667941163
transform 1 0 17756 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_193
timestamp 1667941163
transform 1 0 18860 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1667941163
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1667941163
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1667941163
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1667941163
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1667941163
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1667941163
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1667941163
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1667941163
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1667941163
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1667941163
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1667941163
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1667941163
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1667941163
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_381
timestamp 1667941163
transform 1 0 36156 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_384
timestamp 1667941163
transform 1 0 36432 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_29
timestamp 1667941163
transform 1 0 3772 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_54
timestamp 1667941163
transform 1 0 6072 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_62
timestamp 1667941163
transform 1 0 6808 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_77
timestamp 1667941163
transform 1 0 8188 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_101
timestamp 1667941163
transform 1 0 10396 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_107
timestamp 1667941163
transform 1 0 10948 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1667941163
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_120
timestamp 1667941163
transform 1 0 12144 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_126
timestamp 1667941163
transform 1 0 12696 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_57_135
timestamp 1667941163
transform 1 0 13524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_144
timestamp 1667941163
transform 1 0 14352 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_150
timestamp 1667941163
transform 1 0 14904 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_156
timestamp 1667941163
transform 1 0 15456 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1667941163
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1667941163
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1667941163
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1667941163
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1667941163
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1667941163
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1667941163
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1667941163
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1667941163
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1667941163
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_317
timestamp 1667941163
transform 1 0 30268 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_325
timestamp 1667941163
transform 1 0 31004 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_331
timestamp 1667941163
transform 1 0 31556 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1667941163
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1667941163
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_379
timestamp 1667941163
transform 1 0 35972 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_384
timestamp 1667941163
transform 1 0 36432 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_26
timestamp 1667941163
transform 1 0 3496 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_33
timestamp 1667941163
transform 1 0 4140 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_60
timestamp 1667941163
transform 1 0 6624 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_67
timestamp 1667941163
transform 1 0 7268 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_74
timestamp 1667941163
transform 1 0 7912 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_58_81
timestamp 1667941163
transform 1 0 8556 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_89
timestamp 1667941163
transform 1 0 9292 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_95
timestamp 1667941163
transform 1 0 9844 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_101
timestamp 1667941163
transform 1 0 10396 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_107
timestamp 1667941163
transform 1 0 10948 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_124
timestamp 1667941163
transform 1 0 12512 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_131
timestamp 1667941163
transform 1 0 13156 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_138
timestamp 1667941163
transform 1 0 13800 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_145
timestamp 1667941163
transform 1 0 14444 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_151
timestamp 1667941163
transform 1 0 14996 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_157
timestamp 1667941163
transform 1 0 15548 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_163
timestamp 1667941163
transform 1 0 16100 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_175
timestamp 1667941163
transform 1 0 17204 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_187
timestamp 1667941163
transform 1 0 18308 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1667941163
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1667941163
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1667941163
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1667941163
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1667941163
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1667941163
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1667941163
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1667941163
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1667941163
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1667941163
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1667941163
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1667941163
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1667941163
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1667941163
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_370
timestamp 1667941163
transform 1 0 35144 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_376
timestamp 1667941163
transform 1 0 35696 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_384
timestamp 1667941163
transform 1 0 36432 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_8
timestamp 1667941163
transform 1 0 1840 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_32
timestamp 1667941163
transform 1 0 4048 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_42
timestamp 1667941163
transform 1 0 4968 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_50
timestamp 1667941163
transform 1 0 5704 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_62
timestamp 1667941163
transform 1 0 6808 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_69
timestamp 1667941163
transform 1 0 7452 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_59_98
timestamp 1667941163
transform 1 0 10120 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_106
timestamp 1667941163
transform 1 0 10856 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_110
timestamp 1667941163
transform 1 0 11224 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_129
timestamp 1667941163
transform 1 0 12972 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_136
timestamp 1667941163
transform 1 0 13616 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_142
timestamp 1667941163
transform 1 0 14168 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_148
timestamp 1667941163
transform 1 0 14720 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_154
timestamp 1667941163
transform 1 0 15272 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_166
timestamp 1667941163
transform 1 0 16376 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_180
timestamp 1667941163
transform 1 0 17664 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_192
timestamp 1667941163
transform 1 0 18768 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_204
timestamp 1667941163
transform 1 0 19872 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_216
timestamp 1667941163
transform 1 0 20976 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1667941163
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1667941163
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1667941163
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1667941163
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1667941163
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1667941163
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1667941163
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1667941163
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1667941163
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1667941163
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1667941163
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1667941163
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_385
timestamp 1667941163
transform 1 0 36524 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_25
timestamp 1667941163
transform 1 0 3404 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_37
timestamp 1667941163
transform 1 0 4508 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_47
timestamp 1667941163
transform 1 0 5428 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_76
timestamp 1667941163
transform 1 0 8096 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_82
timestamp 1667941163
transform 1 0 8648 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_108
timestamp 1667941163
transform 1 0 11040 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_125
timestamp 1667941163
transform 1 0 12604 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_131
timestamp 1667941163
transform 1 0 13156 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_137
timestamp 1667941163
transform 1 0 13708 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_145
timestamp 1667941163
transform 1 0 14444 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_151
timestamp 1667941163
transform 1 0 14996 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_160
timestamp 1667941163
transform 1 0 15824 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_167
timestamp 1667941163
transform 1 0 16468 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_179
timestamp 1667941163
transform 1 0 17572 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_191
timestamp 1667941163
transform 1 0 18676 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1667941163
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1667941163
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1667941163
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1667941163
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1667941163
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1667941163
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1667941163
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_289
timestamp 1667941163
transform 1 0 27692 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_294
timestamp 1667941163
transform 1 0 28152 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_300
timestamp 1667941163
transform 1 0 28704 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1667941163
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1667941163
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1667941163
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1667941163
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1667941163
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_377
timestamp 1667941163
transform 1 0 35788 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_385
timestamp 1667941163
transform 1 0 36524 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_25
timestamp 1667941163
transform 1 0 3404 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1667941163
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_61
timestamp 1667941163
transform 1 0 6716 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_88
timestamp 1667941163
transform 1 0 9200 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_97
timestamp 1667941163
transform 1 0 10028 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_104
timestamp 1667941163
transform 1 0 10672 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_110
timestamp 1667941163
transform 1 0 11224 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_125
timestamp 1667941163
transform 1 0 12604 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_131
timestamp 1667941163
transform 1 0 13156 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_137
timestamp 1667941163
transform 1 0 13708 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_143
timestamp 1667941163
transform 1 0 14260 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_149
timestamp 1667941163
transform 1 0 14812 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_155
timestamp 1667941163
transform 1 0 15364 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1667941163
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1667941163
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1667941163
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1667941163
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1667941163
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1667941163
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1667941163
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1667941163
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1667941163
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1667941163
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1667941163
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1667941163
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1667941163
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1667941163
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1667941163
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1667941163
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1667941163
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1667941163
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1667941163
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_373
timestamp 1667941163
transform 1 0 35420 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_376
timestamp 1667941163
transform 1 0 35696 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_384
timestamp 1667941163
transform 1 0 36432 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_26
timestamp 1667941163
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_41
timestamp 1667941163
transform 1 0 4876 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_48
timestamp 1667941163
transform 1 0 5520 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_75
timestamp 1667941163
transform 1 0 8004 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_82
timestamp 1667941163
transform 1 0 8648 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_108
timestamp 1667941163
transform 1 0 11040 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_114
timestamp 1667941163
transform 1 0 11592 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_120
timestamp 1667941163
transform 1 0 12144 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_131
timestamp 1667941163
transform 1 0 13156 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_137
timestamp 1667941163
transform 1 0 13708 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_145
timestamp 1667941163
transform 1 0 14444 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_151
timestamp 1667941163
transform 1 0 14996 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_157
timestamp 1667941163
transform 1 0 15548 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_163
timestamp 1667941163
transform 1 0 16100 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_169
timestamp 1667941163
transform 1 0 16652 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_181
timestamp 1667941163
transform 1 0 17756 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_193
timestamp 1667941163
transform 1 0 18860 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1667941163
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1667941163
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1667941163
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1667941163
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1667941163
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1667941163
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1667941163
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1667941163
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1667941163
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1667941163
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1667941163
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1667941163
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1667941163
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1667941163
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_373
timestamp 1667941163
transform 1 0 35420 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_376
timestamp 1667941163
transform 1 0 35696 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_384
timestamp 1667941163
transform 1 0 36432 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_13
timestamp 1667941163
transform 1 0 2300 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_40
timestamp 1667941163
transform 1 0 4784 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_48
timestamp 1667941163
transform 1 0 5520 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_54
timestamp 1667941163
transform 1 0 6072 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_63
timestamp 1667941163
transform 1 0 6900 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_75
timestamp 1667941163
transform 1 0 8004 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_102
timestamp 1667941163
transform 1 0 10488 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_63_109
timestamp 1667941163
transform 1 0 11132 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_118
timestamp 1667941163
transform 1 0 11960 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_124
timestamp 1667941163
transform 1 0 12512 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_131
timestamp 1667941163
transform 1 0 13156 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_137
timestamp 1667941163
transform 1 0 13708 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_144
timestamp 1667941163
transform 1 0 14352 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_150
timestamp 1667941163
transform 1 0 14904 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_156
timestamp 1667941163
transform 1 0 15456 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_162
timestamp 1667941163
transform 1 0 16008 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_174
timestamp 1667941163
transform 1 0 17112 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_186
timestamp 1667941163
transform 1 0 18216 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_198
timestamp 1667941163
transform 1 0 19320 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_210
timestamp 1667941163
transform 1 0 20424 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 1667941163
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1667941163
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1667941163
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1667941163
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1667941163
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1667941163
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1667941163
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1667941163
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1667941163
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1667941163
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1667941163
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1667941163
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_361
timestamp 1667941163
transform 1 0 34316 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_369
timestamp 1667941163
transform 1 0 35052 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_376
timestamp 1667941163
transform 1 0 35696 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_384
timestamp 1667941163
transform 1 0 36432 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_25
timestamp 1667941163
transform 1 0 3404 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_33
timestamp 1667941163
transform 1 0 4140 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_54
timestamp 1667941163
transform 1 0 6072 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_79
timestamp 1667941163
transform 1 0 8372 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1667941163
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_107
timestamp 1667941163
transform 1 0 10948 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_111
timestamp 1667941163
transform 1 0 11316 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_119
timestamp 1667941163
transform 1 0 12052 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_125
timestamp 1667941163
transform 1 0 12604 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1667941163
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1667941163
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_145
timestamp 1667941163
transform 1 0 14444 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_149
timestamp 1667941163
transform 1 0 14812 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_153
timestamp 1667941163
transform 1 0 15180 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_159
timestamp 1667941163
transform 1 0 15732 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_165
timestamp 1667941163
transform 1 0 16284 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_174
timestamp 1667941163
transform 1 0 17112 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_180
timestamp 1667941163
transform 1 0 17664 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_184
timestamp 1667941163
transform 1 0 18032 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1667941163
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1667941163
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_205
timestamp 1667941163
transform 1 0 19964 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_210
timestamp 1667941163
transform 1 0 20424 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_222
timestamp 1667941163
transform 1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_231
timestamp 1667941163
transform 1 0 22356 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_239
timestamp 1667941163
transform 1 0 23092 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_244
timestamp 1667941163
transform 1 0 23552 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_250
timestamp 1667941163
transform 1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_258
timestamp 1667941163
transform 1 0 24840 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_266
timestamp 1667941163
transform 1 0 25576 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_278
timestamp 1667941163
transform 1 0 26680 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_287
timestamp 1667941163
transform 1 0 27508 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_293
timestamp 1667941163
transform 1 0 28060 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1667941163
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1667941163
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_314
timestamp 1667941163
transform 1 0 29992 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_322
timestamp 1667941163
transform 1 0 30728 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_334
timestamp 1667941163
transform 1 0 31832 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_343
timestamp 1667941163
transform 1 0 32660 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_351
timestamp 1667941163
transform 1 0 33396 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1667941163
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1667941163
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_370
timestamp 1667941163
transform 1 0 35144 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_378
timestamp 1667941163
transform 1 0 35880 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 36892 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 36892 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 36892 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 36892 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 36892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 36892 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 36892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 36892 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 36892 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 36892 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 36892 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 36892 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 36892 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 36892 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 36892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 36892 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 36892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 36892 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 36892 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 36892 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 36892 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 36892 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 36892 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 36892 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 36892 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 36892 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 36892 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 36892 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 36892 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 36892 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 36892 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 36892 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 36892 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 36892 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 36892 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 36892 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 36892 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 36892 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 36892 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 36892 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 36892 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 36892 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 36892 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 36892 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 36892 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 36892 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 36892 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 36892 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 36892 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 36892 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 36892 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 36892 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 36892 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 36892 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 36892 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 36892 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 36892 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 36892 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 36892 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 36892 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 36892 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _134_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 12328 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _135_
timestamp 1667941163
transform 1 0 9660 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _136_
timestamp 1667941163
transform 1 0 13248 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _137_
timestamp 1667941163
transform -1 0 17756 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _138_
timestamp 1667941163
transform 1 0 15548 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _139_
timestamp 1667941163
transform 1 0 10764 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _140_
timestamp 1667941163
transform 1 0 9016 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _141_
timestamp 1667941163
transform 1 0 13248 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _142_
timestamp 1667941163
transform 1 0 14260 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _143_
timestamp 1667941163
transform 1 0 11408 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _144_
timestamp 1667941163
transform 1 0 14260 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _145_
timestamp 1667941163
transform -1 0 18676 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _146_
timestamp 1667941163
transform -1 0 12236 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _147_
timestamp 1667941163
transform -1 0 18584 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _148_
timestamp 1667941163
transform 1 0 17388 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _149_
timestamp 1667941163
transform 1 0 16468 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _150_
timestamp 1667941163
transform 1 0 13340 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _151_
timestamp 1667941163
transform 1 0 12144 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _152_
timestamp 1667941163
transform 1 0 14812 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _153_
timestamp 1667941163
transform -1 0 18032 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _154_
timestamp 1667941163
transform -1 0 12880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _155_
timestamp 1667941163
transform 1 0 8740 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _156_
timestamp 1667941163
transform 1 0 11408 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _157_
timestamp 1667941163
transform 1 0 10948 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _158_
timestamp 1667941163
transform 1 0 13340 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _159_
timestamp 1667941163
transform 1 0 8648 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _160_
timestamp 1667941163
transform 1 0 10304 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _161_
timestamp 1667941163
transform 1 0 12236 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _162_
timestamp 1667941163
transform -1 0 16100 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _163_
timestamp 1667941163
transform 1 0 10764 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _164_
timestamp 1667941163
transform 1 0 10672 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _165_
timestamp 1667941163
transform 1 0 10948 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _166_
timestamp 1667941163
transform -1 0 18400 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _167_
timestamp 1667941163
transform 1 0 11868 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _168_
timestamp 1667941163
transform -1 0 14260 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _169_
timestamp 1667941163
transform 1 0 10304 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _170_
timestamp 1667941163
transform 1 0 12236 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _171_
timestamp 1667941163
transform 1 0 10948 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _172_
timestamp 1667941163
transform 1 0 14628 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _173_
timestamp 1667941163
transform 1 0 10304 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _174_
timestamp 1667941163
transform 1 0 9844 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _175_
timestamp 1667941163
transform 1 0 13340 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _176_
timestamp 1667941163
transform 1 0 11592 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1667941163
transform -1 0 9200 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _178_
timestamp 1667941163
transform 1 0 12880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _179_
timestamp 1667941163
transform 1 0 7176 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp 1667941163
transform -1 0 15732 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _181_
timestamp 1667941163
transform -1 0 18768 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp 1667941163
transform -1 0 10580 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1667941163
transform 1 0 6532 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1667941163
transform 1 0 14260 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _185_
timestamp 1667941163
transform 1 0 14904 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _186_
timestamp 1667941163
transform -1 0 16928 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _187_
timestamp 1667941163
transform 1 0 6164 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp 1667941163
transform -1 0 17572 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _189_
timestamp 1667941163
transform 1 0 14444 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _190_
timestamp 1667941163
transform 1 0 17112 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _191_
timestamp 1667941163
transform 1 0 6532 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _192_
timestamp 1667941163
transform 1 0 9752 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _193_
timestamp 1667941163
transform -1 0 9384 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _194_
timestamp 1667941163
transform -1 0 11040 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _195_
timestamp 1667941163
transform 1 0 7176 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _196_
timestamp 1667941163
transform -1 0 7728 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _197_
timestamp 1667941163
transform 1 0 15548 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _198_
timestamp 1667941163
transform 1 0 14260 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _199_
timestamp 1667941163
transform 1 0 7820 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _200_
timestamp 1667941163
transform 1 0 12880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _201_
timestamp 1667941163
transform -1 0 16284 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _202_
timestamp 1667941163
transform 1 0 13800 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _203_
timestamp 1667941163
transform 1 0 9384 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _204_
timestamp 1667941163
transform 1 0 10948 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _205_
timestamp 1667941163
transform 1 0 12052 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _206_
timestamp 1667941163
transform 1 0 12236 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _207_
timestamp 1667941163
transform 1 0 12788 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _208_
timestamp 1667941163
transform 1 0 18032 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _209_
timestamp 1667941163
transform 1 0 12788 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _210_
timestamp 1667941163
transform -1 0 18308 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _211_
timestamp 1667941163
transform -1 0 11224 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _212_
timestamp 1667941163
transform -1 0 18124 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _213_
timestamp 1667941163
transform -1 0 9844 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _214_
timestamp 1667941163
transform 1 0 11960 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _215_
timestamp 1667941163
transform -1 0 18124 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _216_
timestamp 1667941163
transform -1 0 30544 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _217_
timestamp 1667941163
transform 1 0 19320 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _218_
timestamp 1667941163
transform 1 0 14076 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _219_
timestamp 1667941163
transform -1 0 13708 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 1667941163
transform 1 0 6900 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _221_
timestamp 1667941163
transform -1 0 13800 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1667941163
transform -1 0 18768 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _223_
timestamp 1667941163
transform 1 0 9292 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _224_
timestamp 1667941163
transform -1 0 2024 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _225_
timestamp 1667941163
transform 1 0 5244 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _226_
timestamp 1667941163
transform -1 0 15916 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _227_
timestamp 1667941163
transform -1 0 30728 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1667941163
transform -1 0 31280 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _229_
timestamp 1667941163
transform -1 0 11040 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _230_
timestamp 1667941163
transform -1 0 31464 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _231_
timestamp 1667941163
transform -1 0 6164 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _232_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14352 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _233_
timestamp 1667941163
transform -1 0 18492 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _234_
timestamp 1667941163
transform -1 0 27324 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1667941163
transform -1 0 24656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _236_
timestamp 1667941163
transform -1 0 14904 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _237_
timestamp 1667941163
transform 1 0 15088 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _238_
timestamp 1667941163
transform 1 0 34868 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 1667941163
transform -1 0 22908 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 1667941163
transform 1 0 6532 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _241_
timestamp 1667941163
transform -1 0 13156 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _242_
timestamp 1667941163
transform -1 0 13432 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1667941163
transform 1 0 9108 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _244_
timestamp 1667941163
transform 1 0 5796 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _245_
timestamp 1667941163
transform 1 0 35972 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _246_
timestamp 1667941163
transform 1 0 10212 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _247_
timestamp 1667941163
transform 1 0 9936 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1667941163
transform 1 0 13524 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 1667941163
transform -1 0 15180 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _250_
timestamp 1667941163
transform 1 0 23000 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1667941163
transform -1 0 13156 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1667941163
transform -1 0 28980 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1667941163
transform 1 0 8280 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1667941163
transform -1 0 13800 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1667941163
transform 1 0 12512 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _256_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 4508 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 1667941163
transform 1 0 2852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 1667941163
transform 1 0 2208 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1667941163
transform 1 0 2300 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp 1667941163
transform 1 0 5244 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _261_
timestamp 1667941163
transform -1 0 1840 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp 1667941163
transform 1 0 2392 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _263_
timestamp 1667941163
transform -1 0 4232 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1667941163
transform -1 0 4876 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1667941163
transform 1 0 6532 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 1667941163
transform 1 0 5980 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _267_
timestamp 1667941163
transform -1 0 2300 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _268_
timestamp 1667941163
transform 1 0 6532 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _269_
timestamp 1667941163
transform 1 0 4692 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1667941163
transform -1 0 4232 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1667941163
transform -1 0 1840 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _272_
timestamp 1667941163
transform -1 0 4876 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1667941163
transform 1 0 7820 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _274_
timestamp 1667941163
transform -1 0 7452 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _275_
timestamp 1667941163
transform -1 0 7452 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _276_
timestamp 1667941163
transform -1 0 7912 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _277_
timestamp 1667941163
transform -1 0 6808 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _278_
timestamp 1667941163
transform -1 0 5428 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _279_
timestamp 1667941163
transform 1 0 6532 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1667941163
transform 1 0 4416 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _281_
timestamp 1667941163
transform 1 0 2944 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _282_
timestamp 1667941163
transform 1 0 2208 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _283_
timestamp 1667941163
transform 1 0 2852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _284_
timestamp 1667941163
transform 1 0 2208 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _285_
timestamp 1667941163
transform 1 0 2852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _286_
timestamp 1667941163
transform 1 0 5060 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _287_
timestamp 1667941163
transform 1 0 5888 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _288_
timestamp 1667941163
transform -1 0 1840 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _289_
timestamp 1667941163
transform -1 0 4968 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _290_
timestamp 1667941163
transform 1 0 3036 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _291_
timestamp 1667941163
transform -1 0 1840 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _292_
timestamp 1667941163
transform 1 0 2852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _293_
timestamp 1667941163
transform 1 0 6532 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _294_
timestamp 1667941163
transform 1 0 5704 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1667941163
transform 1 0 7176 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1667941163
transform 1 0 8280 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1667941163
transform -1 0 7268 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1667941163
transform -1 0 7452 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1667941163
transform -1 0 5612 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _300_
timestamp 1667941163
transform 1 0 8372 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _301_
timestamp 1667941163
transform -1 0 5520 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _302_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 10948 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _303_
timestamp 1667941163
transform 1 0 4232 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _304_
timestamp 1667941163
transform -1 0 4784 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _305_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 10396 0 -1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _306_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 8464 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _307_
timestamp 1667941163
transform 1 0 4140 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _308_
timestamp 1667941163
transform -1 0 4048 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _309_
timestamp 1667941163
transform 1 0 1932 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _310_
timestamp 1667941163
transform -1 0 3496 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _311_
timestamp 1667941163
transform -1 0 8004 0 1 35904
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _312_
timestamp 1667941163
transform 1 0 7084 0 -1 35904
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _313_
timestamp 1667941163
transform -1 0 10212 0 -1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _314_
timestamp 1667941163
transform 1 0 1932 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _315_
timestamp 1667941163
transform -1 0 4048 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _316_
timestamp 1667941163
transform 1 0 1656 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _317_
timestamp 1667941163
transform -1 0 6624 0 1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _318_
timestamp 1667941163
transform 1 0 3956 0 -1 35904
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _319_
timestamp 1667941163
transform 1 0 2668 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _320_
timestamp 1667941163
transform 1 0 6532 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _321_
timestamp 1667941163
transform 1 0 4232 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _322_
timestamp 1667941163
transform -1 0 10948 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _323_
timestamp 1667941163
transform -1 0 10120 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _324_
timestamp 1667941163
transform 1 0 7636 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _325_
timestamp 1667941163
transform 1 0 1564 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _326_
timestamp 1667941163
transform -1 0 8188 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _327_
timestamp 1667941163
transform 1 0 6532 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _328_
timestamp 1667941163
transform -1 0 5888 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _329_
timestamp 1667941163
transform -1 0 8096 0 1 34816
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _330_
timestamp 1667941163
transform -1 0 10488 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _331_
timestamp 1667941163
transform 1 0 9108 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _332_
timestamp 1667941163
transform -1 0 8648 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _333_
timestamp 1667941163
transform -1 0 10948 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _334_
timestamp 1667941163
transform 1 0 6808 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _335_
timestamp 1667941163
transform -1 0 8648 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _336_
timestamp 1667941163
transform -1 0 11040 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _337_
timestamp 1667941163
transform 1 0 6716 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _338_
timestamp 1667941163
transform 1 0 1564 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _339_
timestamp 1667941163
transform 1 0 1564 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _340_
timestamp 1667941163
transform -1 0 3404 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _341_
timestamp 1667941163
transform -1 0 6072 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _342_
timestamp 1667941163
transform 1 0 9108 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _343_
timestamp 1667941163
transform 1 0 1564 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _351_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 14352 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _352_
timestamp 1667941163
transform 1 0 14904 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _353_
timestamp 1667941163
transform 1 0 2300 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _354_
timestamp 1667941163
transform 1 0 11684 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _355_
timestamp 1667941163
transform 1 0 31740 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _356_
timestamp 1667941163
transform -1 0 35696 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _357_
timestamp 1667941163
transform -1 0 18860 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _358_
timestamp 1667941163
transform -1 0 27416 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _359_
timestamp 1667941163
transform 1 0 1932 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _360_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 22264 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _361_
timestamp 1667941163
transform 1 0 2300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _362_
timestamp 1667941163
transform 1 0 15640 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _363_
timestamp 1667941163
transform -1 0 25116 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _364_
timestamp 1667941163
transform -1 0 2576 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _365_
timestamp 1667941163
transform -1 0 25668 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _366_
timestamp 1667941163
transform -1 0 33304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _367_
timestamp 1667941163
transform 1 0 2300 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _368_
timestamp 1667941163
transform -1 0 36156 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _369_
timestamp 1667941163
transform -1 0 5980 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _370_
timestamp 1667941163
transform 1 0 35880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _371_
timestamp 1667941163
transform 1 0 10856 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _372_
timestamp 1667941163
transform -1 0 28152 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _373_
timestamp 1667941163
transform 1 0 16284 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _374_
timestamp 1667941163
transform 1 0 1748 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _375_
timestamp 1667941163
transform -1 0 4232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _376_
timestamp 1667941163
transform 1 0 1564 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _377_
timestamp 1667941163
transform -1 0 33672 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _378_
timestamp 1667941163
transform -1 0 17112 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _379_
timestamp 1667941163
transform -1 0 31556 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _380_
timestamp 1667941163
transform 1 0 21160 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _381_
timestamp 1667941163
transform -1 0 36156 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _382_
timestamp 1667941163
transform 1 0 13616 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _383_
timestamp 1667941163
transform 1 0 13156 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _384_
timestamp 1667941163
transform -1 0 6624 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _385_
timestamp 1667941163
transform -1 0 26128 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _386_
timestamp 1667941163
transform 1 0 10856 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _387_
timestamp 1667941163
transform 1 0 14352 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _388_
timestamp 1667941163
transform 1 0 11684 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _389_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 13800 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _390_
timestamp 1667941163
transform 1 0 9292 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _391_
timestamp 1667941163
transform -1 0 16284 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _392_
timestamp 1667941163
transform 1 0 10580 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _393__87 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 17296 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _393_
timestamp 1667941163
transform -1 0 17664 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _394_
timestamp 1667941163
transform 1 0 14260 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _395_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 14444 0 -1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _396_
timestamp 1667941163
transform 1 0 11684 0 1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _397_
timestamp 1667941163
transform -1 0 13708 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _398_
timestamp 1667941163
transform -1 0 15732 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _399_
timestamp 1667941163
transform -1 0 16652 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _400_
timestamp 1667941163
transform 1 0 11316 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _401_
timestamp 1667941163
transform -1 0 8464 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _402__88
timestamp 1667941163
transform -1 0 14720 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _402_
timestamp 1667941163
transform 1 0 14628 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _403_
timestamp 1667941163
transform -1 0 17204 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _404_
timestamp 1667941163
transform -1 0 8188 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _405_
timestamp 1667941163
transform 1 0 10396 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _406_
timestamp 1667941163
transform 1 0 8832 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _407_
timestamp 1667941163
transform -1 0 15916 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _408_
timestamp 1667941163
transform -1 0 15640 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _409_
timestamp 1667941163
transform -1 0 8648 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _410_
timestamp 1667941163
transform 1 0 7360 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _411_
timestamp 1667941163
transform -1 0 15916 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _412_
timestamp 1667941163
transform -1 0 12420 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _413_
timestamp 1667941163
transform -1 0 8004 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _414_
timestamp 1667941163
transform -1 0 7912 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _415_
timestamp 1667941163
transform 1 0 15180 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _416__89
timestamp 1667941163
transform 1 0 16836 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _416_
timestamp 1667941163
transform -1 0 16284 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _417_
timestamp 1667941163
transform -1 0 17480 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _418_
timestamp 1667941163
transform -1 0 15916 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _419_
timestamp 1667941163
transform 1 0 9568 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _420_
timestamp 1667941163
transform -1 0 15180 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _421_
timestamp 1667941163
transform -1 0 8648 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _422_
timestamp 1667941163
transform 1 0 14628 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _423_
timestamp 1667941163
transform -1 0 17112 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _424_
timestamp 1667941163
transform 1 0 14260 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _425_
timestamp 1667941163
transform -1 0 12972 0 -1 34816
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _426_
timestamp 1667941163
transform 1 0 11316 0 1 33728
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _427_
timestamp 1667941163
transform 1 0 10028 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _428__90
timestamp 1667941163
transform -1 0 11224 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _428_
timestamp 1667941163
transform 1 0 12880 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _429_
timestamp 1667941163
transform -1 0 12604 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _430_
timestamp 1667941163
transform 1 0 9108 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _431_
timestamp 1667941163
transform -1 0 17664 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _432_
timestamp 1667941163
transform 1 0 10948 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _433_
timestamp 1667941163
transform 1 0 11408 0 1 34816
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _434_
timestamp 1667941163
transform -1 0 15640 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _435_
timestamp 1667941163
transform -1 0 13616 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _436_
timestamp 1667941163
transform -1 0 13800 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _437_
timestamp 1667941163
transform 1 0 12052 0 -1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _438_
timestamp 1667941163
transform 1 0 12052 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _439_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 14260 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _440_
timestamp 1667941163
transform 1 0 12236 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _440__91
timestamp 1667941163
transform -1 0 10672 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _441_
timestamp 1667941163
transform -1 0 15732 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _442_
timestamp 1667941163
transform 1 0 12604 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _443_
timestamp 1667941163
transform 1 0 13616 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _444_
timestamp 1667941163
transform -1 0 15088 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _445_
timestamp 1667941163
transform 1 0 12236 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _446_
timestamp 1667941163
transform 1 0 12144 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _447_
timestamp 1667941163
transform 1 0 11316 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _448_
timestamp 1667941163
transform 1 0 11040 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _449_
timestamp 1667941163
transform 1 0 14996 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _450_
timestamp 1667941163
transform -1 0 18216 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _451_
timestamp 1667941163
transform 1 0 15272 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _452__92
timestamp 1667941163
transform 1 0 17204 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _452_
timestamp 1667941163
transform 1 0 17112 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _453_
timestamp 1667941163
transform 1 0 12236 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _454_
timestamp 1667941163
transform -1 0 16376 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _455_
timestamp 1667941163
transform 1 0 11776 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _456_
timestamp 1667941163
transform 1 0 13892 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _457_
timestamp 1667941163
transform 1 0 13432 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _458_
timestamp 1667941163
transform -1 0 17020 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _459_
timestamp 1667941163
transform 1 0 15548 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _460_
timestamp 1667941163
transform 1 0 15088 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _461_
timestamp 1667941163
transform 1 0 12052 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _462_
timestamp 1667941163
transform 1 0 16836 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _462__93
timestamp 1667941163
transform -1 0 16468 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _463_
timestamp 1667941163
transform -1 0 14628 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _464_
timestamp 1667941163
transform 1 0 12880 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _465_
timestamp 1667941163
transform -1 0 16376 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _466_
timestamp 1667941163
transform -1 0 13800 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _467_
timestamp 1667941163
transform 1 0 13432 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _468_
timestamp 1667941163
transform 1 0 9292 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _469_
timestamp 1667941163
transform 1 0 10396 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 36432 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1667941163
transform 1 0 16836 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1667941163
transform -1 0 15180 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1667941163
transform -1 0 36432 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1667941163
transform -1 0 4876 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1667941163
transform -1 0 1840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1667941163
transform 1 0 10396 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1667941163
transform 1 0 13432 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1667941163
transform -1 0 36432 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1667941163
transform 1 0 1564 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1667941163
transform 1 0 36156 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1667941163
transform 1 0 9108 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1667941163
transform -1 0 35880 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1667941163
transform 1 0 1564 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1667941163
transform 1 0 1564 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1667941163
transform -1 0 25576 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1667941163
transform -1 0 34408 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1667941163
transform 1 0 35512 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1667941163
transform 1 0 23276 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1667941163
transform -1 0 36432 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1667941163
transform 1 0 1564 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1667941163
transform -1 0 3496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1667941163
transform 1 0 10396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1667941163
transform -1 0 32660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1667941163
transform 1 0 36156 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1667941163
transform 1 0 36156 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1667941163
transform 1 0 24564 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1667941163
transform -1 0 5704 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input29
timestamp 1667941163
transform -1 0 36432 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1667941163
transform -1 0 10028 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1667941163
transform -1 0 36432 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1667941163
transform -1 0 1840 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1667941163
transform 1 0 29716 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1667941163
transform 1 0 1564 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input35
timestamp 1667941163
transform -1 0 2484 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1667941163
transform 1 0 12972 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1667941163
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1667941163
transform -1 0 2576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1667941163
transform 1 0 21988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input40 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 30360 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1667941163
transform -1 0 1932 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1667941163
transform 1 0 36064 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1667941163
transform 1 0 36064 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1667941163
transform 1 0 27140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1667941163
transform 1 0 36064 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1667941163
transform 1 0 6532 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1667941163
transform -1 0 1932 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1667941163
transform 1 0 36064 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1667941163
transform 1 0 20056 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1667941163
transform 1 0 36064 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1667941163
transform -1 0 27508 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1667941163
transform -1 0 1932 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1667941163
transform -1 0 1932 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1667941163
transform -1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1667941163
transform 1 0 18124 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1667941163
transform 1 0 36064 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1667941163
transform -1 0 1932 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1667941163
transform 1 0 34776 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1667941163
transform 1 0 36064 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1667941163
transform 1 0 3956 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1667941163
transform 1 0 31004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1667941163
transform -1 0 15272 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1667941163
transform -1 0 1932 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1667941163
transform 1 0 36064 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1667941163
transform 1 0 11684 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1667941163
transform 1 0 21988 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1667941163
transform 1 0 33580 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1667941163
transform 1 0 1564 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1667941163
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1667941163
transform -1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1667941163
transform 1 0 36064 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1667941163
transform 1 0 28428 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1667941163
transform 1 0 16836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1667941163
transform -1 0 35696 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1667941163
transform 1 0 36064 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1667941163
transform -1 0 5520 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1667941163
transform 1 0 36064 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1667941163
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1667941163
transform -1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1667941163
transform -1 0 1932 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1667941163
transform 1 0 36064 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1667941163
transform -1 0 20424 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1667941163
transform 1 0 32292 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1667941163
transform -1 0 8004 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1667941163
transform 1 0 25852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1667941163
transform -1 0 1932 0 -1 13056
box -38 -48 406 592
<< labels >>
flabel metal3 s 200 19728 800 19848 0 FreeSans 480 0 0 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_
port 0 nsew signal tristate
flabel metal3 s 37200 33328 37800 33448 0 FreeSans 480 0 0 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_
port 1 nsew signal tristate
flabel metal3 s 37200 8168 37800 8288 0 FreeSans 480 0 0 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_
port 2 nsew signal tristate
flabel metal2 s 27066 200 27122 800 0 FreeSans 224 90 0 0 bottom_grid_top_width_0_height_0_subtile_0__pin_clk_0_
port 3 nsew signal tristate
flabel metal3 s 37200 31968 37800 32088 0 FreeSans 480 0 0 0 ccff_head
port 4 nsew signal input
flabel metal3 s 37200 24488 37800 24608 0 FreeSans 480 0 0 0 ccff_tail
port 5 nsew signal tristate
flabel metal2 s 16118 39200 16174 39800 0 FreeSans 224 90 0 0 chanx_left_in[0]
port 6 nsew signal input
flabel metal2 s 14830 39200 14886 39800 0 FreeSans 224 90 0 0 chanx_left_in[10]
port 7 nsew signal input
flabel metal3 s 37200 15648 37800 15768 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 8 nsew signal input
flabel metal2 s 662 39200 718 39800 0 FreeSans 224 90 0 0 chanx_left_in[12]
port 9 nsew signal input
flabel metal3 s 200 4768 800 4888 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 10 nsew signal input
flabel metal3 s 200 36048 800 36168 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 11 nsew signal input
flabel metal2 s 13542 200 13598 800 0 FreeSans 224 90 0 0 chanx_left_in[15]
port 12 nsew signal input
flabel metal3 s 37200 29928 37800 30048 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 13 nsew signal input
flabel metal3 s 200 28568 800 28688 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 14 nsew signal input
flabel metal3 s 37200 26528 37800 26648 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 15 nsew signal input
flabel metal2 s 8390 200 8446 800 0 FreeSans 224 90 0 0 chanx_left_in[1]
port 16 nsew signal input
flabel metal2 s 35438 39200 35494 39800 0 FreeSans 224 90 0 0 chanx_left_in[2]
port 17 nsew signal input
flabel metal3 s 200 30608 800 30728 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 18 nsew signal input
flabel metal3 s 200 14288 800 14408 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 19 nsew signal input
flabel metal2 s 25134 39200 25190 39800 0 FreeSans 224 90 0 0 chanx_left_in[5]
port 20 nsew signal input
flabel metal2 s 34150 200 34206 800 0 FreeSans 224 90 0 0 chanx_left_in[6]
port 21 nsew signal input
flabel metal2 s 35438 200 35494 800 0 FreeSans 224 90 0 0 chanx_left_in[7]
port 22 nsew signal input
flabel metal2 s 23202 39200 23258 39800 0 FreeSans 224 90 0 0 chanx_left_in[8]
port 23 nsew signal input
flabel metal3 s 37200 27888 37800 28008 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 24 nsew signal input
flabel metal2 s 5814 39200 5870 39800 0 FreeSans 224 90 0 0 chanx_left_out[0]
port 25 nsew signal tristate
flabel metal3 s 200 23128 800 23248 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 26 nsew signal tristate
flabel metal3 s 37200 17008 37800 17128 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 27 nsew signal tristate
flabel metal2 s 19982 39200 20038 39800 0 FreeSans 224 90 0 0 chanx_left_out[12]
port 28 nsew signal tristate
flabel metal3 s 37200 4768 37800 4888 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 29 nsew signal tristate
flabel metal2 s 26422 39200 26478 39800 0 FreeSans 224 90 0 0 chanx_left_out[14]
port 30 nsew signal tristate
flabel metal3 s 200 3408 800 3528 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 31 nsew signal tristate
flabel metal3 s 200 10208 800 10328 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 32 nsew signal tristate
flabel metal3 s 200 1368 800 1488 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 33 nsew signal tristate
flabel metal2 s 18050 39200 18106 39800 0 FreeSans 224 90 0 0 chanx_left_out[18]
port 34 nsew signal tristate
flabel metal3 s 37200 38768 37800 38888 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 35 nsew signal tristate
flabel metal3 s 200 21088 800 21208 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 36 nsew signal tristate
flabel metal3 s 37200 688 37800 808 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 37 nsew signal tristate
flabel metal3 s 37200 13608 37800 13728 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 38 nsew signal tristate
flabel metal3 s 200 39448 800 39568 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 39 nsew signal tristate
flabel metal2 s 30286 200 30342 800 0 FreeSans 224 90 0 0 chanx_left_out[6]
port 40 nsew signal tristate
flabel metal2 s 14830 200 14886 800 0 FreeSans 224 90 0 0 chanx_left_out[7]
port 41 nsew signal tristate
flabel metal3 s 200 6808 800 6928 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 42 nsew signal tristate
flabel metal3 s 37200 35368 37800 35488 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 43 nsew signal tristate
flabel metal3 s 200 8848 800 8968 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 44 nsew signal input
flabel metal2 s 3238 200 3294 800 0 FreeSans 224 90 0 0 chanx_right_in[10]
port 45 nsew signal input
flabel metal2 s 9678 200 9734 800 0 FreeSans 224 90 0 0 chanx_right_in[11]
port 46 nsew signal input
flabel metal2 s 32218 200 32274 800 0 FreeSans 224 90 0 0 chanx_right_in[12]
port 47 nsew signal input
flabel metal3 s 37200 11568 37800 11688 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 48 nsew signal input
flabel metal3 s 37200 6128 37800 6248 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 49 nsew signal input
flabel metal2 s 23846 200 23902 800 0 FreeSans 224 90 0 0 chanx_right_in[15]
port 50 nsew signal input
flabel metal3 s 200 37408 800 37528 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 51 nsew signal input
flabel metal2 s 37370 200 37426 800 0 FreeSans 224 90 0 0 chanx_right_in[17]
port 52 nsew signal input
flabel metal2 s 9678 39200 9734 39800 0 FreeSans 224 90 0 0 chanx_right_in[18]
port 53 nsew signal input
flabel metal3 s 37200 10208 37800 10328 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 54 nsew signal input
flabel metal3 s 200 25168 800 25288 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 55 nsew signal input
flabel metal2 s 28998 200 29054 800 0 FreeSans 224 90 0 0 chanx_right_in[3]
port 56 nsew signal input
flabel metal3 s 200 17688 800 17808 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 57 nsew signal input
flabel metal3 s 200 31968 800 32088 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 58 nsew signal input
flabel metal2 s 12898 39200 12954 39800 0 FreeSans 224 90 0 0 chanx_right_in[6]
port 59 nsew signal input
flabel metal2 s 18694 200 18750 800 0 FreeSans 224 90 0 0 chanx_right_in[7]
port 60 nsew signal input
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 chanx_right_in[8]
port 61 nsew signal input
flabel metal2 s 21914 200 21970 800 0 FreeSans 224 90 0 0 chanx_right_in[9]
port 62 nsew signal input
flabel metal2 s 10966 39200 11022 39800 0 FreeSans 224 90 0 0 chanx_right_out[0]
port 63 nsew signal tristate
flabel metal2 s 21270 39200 21326 39800 0 FreeSans 224 90 0 0 chanx_right_out[10]
port 64 nsew signal tristate
flabel metal2 s 33506 39200 33562 39800 0 FreeSans 224 90 0 0 chanx_right_out[11]
port 65 nsew signal tristate
flabel metal3 s 200 26528 800 26648 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 66 nsew signal tristate
flabel metal2 s 4526 200 4582 800 0 FreeSans 224 90 0 0 chanx_right_out[13]
port 67 nsew signal tristate
flabel metal2 s 1306 200 1362 800 0 FreeSans 224 90 0 0 chanx_right_out[14]
port 68 nsew signal tristate
flabel metal2 s 36726 39200 36782 39800 0 FreeSans 224 90 0 0 chanx_right_out[15]
port 69 nsew signal tristate
flabel metal2 s 28354 39200 28410 39800 0 FreeSans 224 90 0 0 chanx_right_out[16]
port 70 nsew signal tristate
flabel metal2 s 16762 200 16818 800 0 FreeSans 224 90 0 0 chanx_right_out[17]
port 71 nsew signal tristate
flabel metal3 s 37200 37408 37800 37528 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 72 nsew signal tristate
flabel metal3 s 37200 2728 37800 2848 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 73 nsew signal tristate
flabel metal2 s 4526 39200 4582 39800 0 FreeSans 224 90 0 0 chanx_right_out[2]
port 74 nsew signal tristate
flabel metal3 s 37200 21088 37800 21208 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 75 nsew signal tristate
flabel metal2 s 6458 200 6514 800 0 FreeSans 224 90 0 0 chanx_right_out[4]
port 76 nsew signal tristate
flabel metal2 s 11610 200 11666 800 0 FreeSans 224 90 0 0 chanx_right_out[5]
port 77 nsew signal tristate
flabel metal3 s 200 15648 800 15768 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 78 nsew signal tristate
flabel metal3 s 37200 22448 37800 22568 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 79 nsew signal tristate
flabel metal2 s 19982 200 20038 800 0 FreeSans 224 90 0 0 chanx_right_out[8]
port 80 nsew signal tristate
flabel metal2 s 31574 39200 31630 39800 0 FreeSans 224 90 0 0 chanx_right_out[9]
port 81 nsew signal tristate
flabel metal2 s 30286 39200 30342 39800 0 FreeSans 224 90 0 0 pReset
port 82 nsew signal input
flabel metal2 s 2594 39200 2650 39800 0 FreeSans 224 90 0 0 prog_clk
port 83 nsew signal input
flabel metal2 s 7746 39200 7802 39800 0 FreeSans 224 90 0 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_
port 84 nsew signal tristate
flabel metal2 s 25134 200 25190 800 0 FreeSans 224 90 0 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_
port 85 nsew signal tristate
flabel metal3 s 200 12248 800 12368 0 FreeSans 480 0 0 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_
port 86 nsew signal tristate
flabel metal3 s 200 34008 800 34128 0 FreeSans 480 0 0 0 vccd1
port 87 nsew signal bidirectional
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 87 nsew signal bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 87 nsew signal bidirectional
flabel metal3 s 37200 19048 37800 19168 0 FreeSans 480 0 0 0 vssd1
port 88 nsew signal bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 88 nsew signal bidirectional
rlabel metal1 18998 37536 18998 37536 0 vccd1
rlabel metal1 18998 36992 18998 36992 0 vssd1
rlabel metal1 4554 29546 4554 29546 0 _000_
rlabel metal2 5566 29138 5566 29138 0 _001_
rlabel metal2 3082 29886 3082 29886 0 _002_
rlabel metal1 6900 31994 6900 31994 0 _003_
rlabel metal2 9246 31433 9246 31433 0 _004_
rlabel metal1 4186 27472 4186 27472 0 _005_
rlabel metal1 3680 31994 3680 31994 0 _006_
rlabel metal1 4186 29750 4186 29750 0 _007_
rlabel metal1 2744 33898 2744 33898 0 _008_
rlabel metal1 6210 33082 6210 33082 0 _009_
rlabel metal1 6900 33626 6900 33626 0 _010_
rlabel metal1 5152 32878 5152 32878 0 _011_
rlabel metal1 4048 29818 4048 29818 0 _012_
rlabel metal1 1702 32436 1702 32436 0 _013_
rlabel metal1 4692 31994 4692 31994 0 _014_
rlabel metal1 6033 33898 6033 33898 0 _015_
rlabel metal1 7176 32538 7176 32538 0 _016_
rlabel metal1 7084 34714 7084 34714 0 _017_
rlabel metal1 7820 34170 7820 34170 0 _018_
rlabel metal1 6210 34714 6210 34714 0 _019_
rlabel metal1 9009 37162 9009 37162 0 _020_
rlabel metal1 6532 32198 6532 32198 0 _021_
rlabel metal1 8365 30294 8365 30294 0 _022_
rlabel metal2 2346 30056 2346 30056 0 _023_
rlabel metal1 4823 28458 4823 28458 0 _024_
rlabel metal1 5934 28696 5934 28696 0 _025_
rlabel metal1 3910 31926 3910 31926 0 _026_
rlabel metal1 5290 32266 5290 32266 0 _027_
rlabel metal1 6256 31926 6256 31926 0 _028_
rlabel metal2 9890 35394 9890 35394 0 _029_
rlabel metal1 5198 27574 5198 27574 0 _030_
rlabel metal2 1702 28254 1702 28254 0 _031_
rlabel metal1 3128 28186 3128 28186 0 _032_
rlabel metal2 6670 32674 6670 32674 0 _033_
rlabel metal1 6716 32334 6716 32334 0 _034_
rlabel metal2 7314 31586 7314 31586 0 _035_
rlabel metal1 7590 34034 7590 34034 0 _036_
rlabel metal1 6486 34170 6486 34170 0 _037_
rlabel metal1 2698 34986 2698 34986 0 _038_
rlabel metal2 5474 33320 5474 33320 0 _039_
rlabel metal1 9108 36006 9108 36006 0 _040_
rlabel metal1 4239 36074 4239 36074 0 _041_
rlabel metal1 2346 28050 2346 28050 0 _042_
rlabel metal1 4738 32912 4738 32912 0 _043_
rlabel metal2 2898 28730 2898 28730 0 _044_
rlabel metal1 1794 28492 1794 28492 0 _045_
rlabel metal2 13570 26520 13570 26520 0 _046_
rlabel metal2 9522 25194 9522 25194 0 _047_
rlabel metal2 16054 27608 16054 27608 0 _048_
rlabel metal2 11086 28322 11086 28322 0 _049_
rlabel metal2 18170 29002 18170 29002 0 _050_
rlabel metal1 14490 30600 14490 30600 0 _051_
rlabel metal1 13570 32198 13570 32198 0 _052_
rlabel metal2 11914 31144 11914 31144 0 _053_
rlabel metal2 12466 27846 12466 27846 0 _054_
rlabel metal2 15502 28322 15502 28322 0 _055_
rlabel metal1 17296 29070 17296 29070 0 _056_
rlabel metal1 10534 29274 10534 29274 0 _057_
rlabel metal2 8234 25262 8234 25262 0 _058_
rlabel metal1 14628 20570 14628 20570 0 _059_
rlabel metal2 16974 19482 16974 19482 0 _060_
rlabel metal1 7636 21590 7636 21590 0 _061_
rlabel metal1 10764 22202 10764 22202 0 _062_
rlabel metal1 9154 22202 9154 22202 0 _063_
rlabel metal1 14812 21590 14812 21590 0 _064_
rlabel metal1 15410 21896 15410 21896 0 _065_
rlabel metal1 8418 24072 8418 24072 0 _066_
rlabel metal2 7590 19176 7590 19176 0 _067_
rlabel metal1 14352 22746 14352 22746 0 _068_
rlabel metal1 11040 24582 11040 24582 0 _069_
rlabel metal2 6302 26792 6302 26792 0 _070_
rlabel metal2 7682 26826 7682 26826 0 _071_
rlabel metal2 15410 23902 15410 23902 0 _072_
rlabel metal2 16054 24344 16054 24344 0 _073_
rlabel metal2 17250 26690 17250 26690 0 _074_
rlabel metal1 15686 25160 15686 25160 0 _075_
rlabel metal1 10120 27098 10120 27098 0 _076_
rlabel metal1 15272 28118 15272 28118 0 _077_
rlabel metal1 8418 27336 8418 27336 0 _078_
rlabel metal2 14858 23630 14858 23630 0 _079_
rlabel metal1 17158 24378 17158 24378 0 _080_
rlabel metal1 14490 29512 14490 29512 0 _081_
rlabel metal1 13110 34646 13110 34646 0 _082_
rlabel metal2 11546 34136 11546 34136 0 _083_
rlabel metal1 10120 29206 10120 29206 0 _084_
rlabel metal2 13202 29818 13202 29818 0 _085_
rlabel metal2 13018 34986 13018 34986 0 _086_
rlabel metal1 9200 24922 9200 24922 0 _087_
rlabel metal1 12558 27574 12558 27574 0 _088_
rlabel metal1 11224 24106 11224 24106 0 _089_
rlabel metal1 11822 33626 11822 33626 0 _090_
rlabel metal1 15088 31790 15088 31790 0 _091_
rlabel metal2 12650 26282 12650 26282 0 _092_
rlabel metal1 13846 28390 13846 28390 0 _093_
rlabel metal1 12282 25976 12282 25976 0 _094_
rlabel metal2 12282 25806 12282 25806 0 _095_
rlabel metal1 14306 22610 14306 22610 0 _096_
rlabel metal2 12374 22916 12374 22916 0 _097_
rlabel metal2 18262 25976 18262 25976 0 _098_
rlabel metal2 13110 26248 13110 26248 0 _099_
rlabel metal1 13662 23290 13662 23290 0 _100_
rlabel metal1 13754 24072 13754 24072 0 _101_
rlabel metal1 11730 24820 11730 24820 0 _102_
rlabel metal1 11178 23766 11178 23766 0 _103_
rlabel metal1 11546 26248 11546 26248 0 _104_
rlabel metal2 11546 22610 11546 22610 0 _105_
rlabel metal1 14628 29206 14628 29206 0 _106_
rlabel metal2 18446 26656 18446 26656 0 _107_
rlabel metal1 14490 30294 14490 30294 0 _108_
rlabel metal1 17204 26282 17204 26282 0 _109_
rlabel metal2 12466 29614 12466 29614 0 _110_
rlabel metal2 17894 26418 17894 26418 0 _111_
rlabel metal2 12006 29240 12006 29240 0 _112_
rlabel metal1 14122 25976 14122 25976 0 _113_
rlabel metal1 13202 29206 13202 29206 0 _114_
rlabel metal1 16790 28424 16790 28424 0 _115_
rlabel metal1 15364 27574 15364 27574 0 _116_
rlabel metal2 15318 26180 15318 26180 0 _117_
rlabel metal1 11132 31790 11132 31790 0 _118_
rlabel metal2 15686 34782 15686 34782 0 _119_
rlabel metal2 14398 27710 14398 27710 0 _120_
rlabel metal2 13110 28968 13110 28968 0 _121_
rlabel metal1 16376 24854 16376 24854 0 _122_
rlabel metal2 13570 33048 13570 33048 0 _123_
rlabel metal1 13064 32470 13064 32470 0 _124_
rlabel metal1 9338 27098 9338 27098 0 _125_
rlabel metal2 10626 25806 10626 25806 0 _126_
rlabel metal3 1188 19788 1188 19788 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_
rlabel via2 36294 33371 36294 33371 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_
rlabel metal2 36294 8279 36294 8279 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_
rlabel metal2 27094 1520 27094 1520 0 bottom_grid_top_width_0_height_0_subtile_0__pin_clk_0_
rlabel metal2 36386 32181 36386 32181 0 ccff_head
rlabel via2 36294 24565 36294 24565 0 ccff_tail
rlabel metal1 16836 37230 16836 37230 0 chanx_left_in[0]
rlabel metal1 14904 37230 14904 37230 0 chanx_left_in[10]
rlabel via2 36386 15691 36386 15691 0 chanx_left_in[11]
rlabel metal2 690 38430 690 38430 0 chanx_left_in[12]
rlabel metal2 1610 5015 1610 5015 0 chanx_left_in[13]
rlabel metal1 10534 35666 10534 35666 0 chanx_left_in[14]
rlabel metal2 13570 1554 13570 1554 0 chanx_left_in[15]
rlabel metal2 36386 29903 36386 29903 0 chanx_left_in[16]
rlabel metal2 1610 28849 1610 28849 0 chanx_left_in[17]
rlabel metal2 36386 26775 36386 26775 0 chanx_left_in[18]
rlabel metal1 8464 2278 8464 2278 0 chanx_left_in[1]
rlabel metal1 35282 37434 35282 37434 0 chanx_left_in[2]
rlabel metal1 1610 30634 1610 30634 0 chanx_left_in[3]
rlabel via2 1702 14331 1702 14331 0 chanx_left_in[4]
rlabel metal1 24978 37434 24978 37434 0 chanx_left_in[5]
rlabel metal1 34224 2346 34224 2346 0 chanx_left_in[6]
rlabel metal1 34592 2414 34592 2414 0 chanx_left_in[7]
rlabel metal2 23506 38233 23506 38233 0 chanx_left_in[8]
rlabel via2 36386 27965 36386 27965 0 chanx_left_in[9]
rlabel metal1 6302 36890 6302 36890 0 chanx_left_out[0]
rlabel metal3 1188 23188 1188 23188 0 chanx_left_out[10]
rlabel via2 36294 17051 36294 17051 0 chanx_left_out[11]
rlabel metal1 20148 37094 20148 37094 0 chanx_left_out[12]
rlabel metal2 36294 4913 36294 4913 0 chanx_left_out[13]
rlabel metal1 26864 37094 26864 37094 0 chanx_left_out[14]
rlabel metal3 1188 3468 1188 3468 0 chanx_left_out[15]
rlabel metal3 1188 10268 1188 10268 0 chanx_left_out[16]
rlabel metal3 1188 1428 1188 1428 0 chanx_left_out[17]
rlabel metal1 18216 37094 18216 37094 0 chanx_left_out[18]
rlabel metal2 35834 37859 35834 37859 0 chanx_left_out[1]
rlabel metal3 1188 21148 1188 21148 0 chanx_left_out[2]
rlabel metal2 36570 1785 36570 1785 0 chanx_left_out[3]
rlabel via2 36294 13685 36294 13685 0 chanx_left_out[4]
rlabel metal1 4370 32742 4370 32742 0 chanx_left_out[5]
rlabel metal2 30314 1520 30314 1520 0 chanx_left_out[6]
rlabel metal2 14858 1520 14858 1520 0 chanx_left_out[7]
rlabel metal3 1188 6868 1188 6868 0 chanx_left_out[8]
rlabel via2 36294 35445 36294 35445 0 chanx_left_out[9]
rlabel via2 1610 8925 1610 8925 0 chanx_right_in[0]
rlabel metal1 3312 2346 3312 2346 0 chanx_right_in[10]
rlabel metal1 10120 2346 10120 2346 0 chanx_right_in[11]
rlabel metal1 32384 2346 32384 2346 0 chanx_right_in[12]
rlabel metal2 36386 11679 36386 11679 0 chanx_right_in[13]
rlabel metal2 36386 6239 36386 6239 0 chanx_right_in[14]
rlabel metal1 23920 2278 23920 2278 0 chanx_right_in[15]
rlabel metal2 9982 34663 9982 34663 0 chanx_right_in[16]
rlabel metal1 36892 2958 36892 2958 0 chanx_right_in[17]
rlabel metal2 9798 36159 9798 36159 0 chanx_right_in[18]
rlabel via2 36386 10251 36386 10251 0 chanx_right_in[1]
rlabel via2 1610 25245 1610 25245 0 chanx_right_in[2]
rlabel metal1 29072 2278 29072 2278 0 chanx_right_in[3]
rlabel via2 1610 17765 1610 17765 0 chanx_right_in[4]
rlabel metal3 1464 32028 1464 32028 0 chanx_right_in[5]
rlabel metal1 13018 37230 13018 37230 0 chanx_right_in[6]
rlabel metal1 18768 2278 18768 2278 0 chanx_right_in[7]
rlabel metal2 2346 1870 2346 1870 0 chanx_right_in[8]
rlabel metal2 21942 1554 21942 1554 0 chanx_right_in[9]
rlabel metal1 11500 37094 11500 37094 0 chanx_right_out[0]
rlabel metal1 21758 37094 21758 37094 0 chanx_right_out[10]
rlabel metal1 33672 37094 33672 37094 0 chanx_right_out[11]
rlabel metal3 1234 26588 1234 26588 0 chanx_right_out[12]
rlabel metal2 4554 1520 4554 1520 0 chanx_right_out[13]
rlabel metal2 1334 1520 1334 1520 0 chanx_right_out[14]
rlabel metal1 36524 36346 36524 36346 0 chanx_right_out[15]
rlabel metal1 28520 37094 28520 37094 0 chanx_right_out[16]
rlabel metal2 16790 1520 16790 1520 0 chanx_right_out[17]
rlabel metal1 35558 36890 35558 36890 0 chanx_right_out[18]
rlabel metal2 36294 3077 36294 3077 0 chanx_right_out[1]
rlabel metal1 4968 36890 4968 36890 0 chanx_right_out[2]
rlabel metal2 36294 21233 36294 21233 0 chanx_right_out[3]
rlabel metal2 6486 1520 6486 1520 0 chanx_right_out[4]
rlabel metal2 11638 1520 11638 1520 0 chanx_right_out[5]
rlabel metal3 1188 15708 1188 15708 0 chanx_right_out[6]
rlabel via2 36294 22491 36294 22491 0 chanx_right_out[7]
rlabel metal2 20010 1520 20010 1520 0 chanx_right_out[8]
rlabel metal1 32154 37094 32154 37094 0 chanx_right_out[9]
rlabel metal1 8694 31246 8694 31246 0 mem_bottom_ipin_0.DFFR_0_.Q
rlabel metal1 12834 31858 12834 31858 0 mem_bottom_ipin_0.DFFR_1_.Q
rlabel metal2 18078 27812 18078 27812 0 mem_bottom_ipin_0.DFFR_2_.Q
rlabel metal1 5244 30158 5244 30158 0 mem_bottom_ipin_0.DFFR_3_.Q
rlabel metal2 8050 30226 8050 30226 0 mem_bottom_ipin_0.DFFR_4_.Q
rlabel metal1 12834 32368 12834 32368 0 mem_bottom_ipin_0.DFFR_5_.Q
rlabel metal1 8326 20026 8326 20026 0 mem_bottom_ipin_1.DFFR_0_.Q
rlabel metal1 16238 22032 16238 22032 0 mem_bottom_ipin_1.DFFR_1_.Q
rlabel metal2 13846 21675 13846 21675 0 mem_bottom_ipin_1.DFFR_2_.Q
rlabel via1 2254 33626 2254 33626 0 mem_bottom_ipin_1.DFFR_3_.Q
rlabel metal1 4830 33422 4830 33422 0 mem_bottom_ipin_1.DFFR_4_.Q
rlabel metal1 2346 34714 2346 34714 0 mem_bottom_ipin_1.DFFR_5_.Q
rlabel metal1 8970 34986 8970 34986 0 mem_bottom_ipin_2.DFFR_0_.Q
rlabel metal1 10856 34918 10856 34918 0 mem_bottom_ipin_2.DFFR_1_.Q
rlabel metal2 13294 33660 13294 33660 0 mem_bottom_ipin_2.DFFR_2_.Q
rlabel metal1 12374 32980 12374 32980 0 mem_bottom_ipin_2.DFFR_3_.Q
rlabel metal1 1886 35768 1886 35768 0 mem_bottom_ipin_2.DFFR_4_.Q
rlabel metal2 15594 35326 15594 35326 0 mem_bottom_ipin_2.DFFR_5_.Q
rlabel metal1 13386 35666 13386 35666 0 mem_top_ipin_0.DFFR_0_.Q
rlabel metal1 17158 25772 17158 25772 0 mem_top_ipin_0.DFFR_1_.Q
rlabel metal1 13524 33082 13524 33082 0 mem_top_ipin_0.DFFR_2_.Q
rlabel metal1 5796 27506 5796 27506 0 mem_top_ipin_0.DFFR_3_.Q
rlabel metal1 2438 31246 2438 31246 0 mem_top_ipin_0.DFFR_4_.Q
rlabel metal2 3726 29240 3726 29240 0 mem_top_ipin_0.DFFR_5_.Q
rlabel metal1 14398 31790 14398 31790 0 mem_top_ipin_1.DFFR_0_.Q
rlabel metal1 12926 34000 12926 34000 0 mem_top_ipin_1.DFFR_1_.Q
rlabel metal1 8878 34510 8878 34510 0 mem_top_ipin_1.DFFR_2_.Q
rlabel metal1 9246 37298 9246 37298 0 mem_top_ipin_1.DFFR_3_.Q
rlabel metal1 6762 37162 6762 37162 0 mem_top_ipin_1.DFFR_4_.Q
rlabel metal1 10212 36210 10212 36210 0 mem_top_ipin_1.DFFR_5_.Q
rlabel metal1 10902 22066 10902 22066 0 mem_top_ipin_2.DFFR_0_.Q
rlabel metal2 12742 24650 12742 24650 0 mem_top_ipin_2.DFFR_1_.Q
rlabel metal1 12236 21114 12236 21114 0 mem_top_ipin_2.DFFR_2_.Q
rlabel metal1 6670 29206 6670 29206 0 mem_top_ipin_2.DFFR_3_.Q
rlabel metal1 8740 29002 8740 29002 0 mem_top_ipin_2.DFFR_4_.Q
rlabel metal1 7176 28390 7176 28390 0 mem_top_ipin_2.DFFR_5_.Q
rlabel metal1 14536 32810 14536 32810 0 mem_top_ipin_3.DFFR_0_.Q
rlabel metal1 8602 32810 8602 32810 0 mem_top_ipin_3.DFFR_1_.Q
rlabel viali 16514 26355 16514 26355 0 mem_top_ipin_3.DFFR_2_.Q
rlabel metal1 11040 31858 11040 31858 0 mem_top_ipin_3.DFFR_3_.Q
rlabel metal1 11500 32402 11500 32402 0 mem_top_ipin_3.DFFR_4_.Q
rlabel metal2 13478 26095 13478 26095 0 mux_bottom_ipin_0.INVTX1_0_.out
rlabel metal1 8004 22066 8004 22066 0 mux_bottom_ipin_0.INVTX1_1_.out
rlabel metal1 13846 22066 13846 22066 0 mux_bottom_ipin_0.INVTX1_2_.out
rlabel metal1 15686 27948 15686 27948 0 mux_bottom_ipin_0.INVTX1_3_.out
rlabel metal1 10764 28594 10764 28594 0 mux_bottom_ipin_0.INVTX1_4_.out
rlabel metal1 17066 27506 17066 27506 0 mux_bottom_ipin_0.INVTX1_5_.out
rlabel metal1 16698 29546 16698 29546 0 mux_bottom_ipin_0.INVTX1_6_.out
rlabel metal1 14306 33286 14306 33286 0 mux_bottom_ipin_0.INVTX1_7_.out
rlabel metal2 13018 25296 13018 25296 0 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 11592 30634 11592 30634 0 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 16238 29444 16238 29444 0 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 19688 3026 19688 3026 0 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 10534 23630 10534 23630 0 mux_bottom_ipin_1.INVTX1_2_.out
rlabel metal1 16146 23018 16146 23018 0 mux_bottom_ipin_1.INVTX1_3_.out
rlabel metal2 30590 21522 30590 21522 0 mux_bottom_ipin_1.INVTX1_4_.out
rlabel metal2 15778 14756 15778 14756 0 mux_bottom_ipin_1.INVTX1_5_.out
rlabel metal1 6394 9622 6394 9622 0 mux_bottom_ipin_1.INVTX1_6_.out
rlabel metal1 17388 18666 17388 18666 0 mux_bottom_ipin_1.INVTX1_7_.out
rlabel metal1 11408 22678 11408 22678 0 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 15042 22134 15042 22134 0 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 15916 20842 15916 20842 0 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 7360 21454 7360 21454 0 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 13662 33320 13662 33320 0 mux_bottom_ipin_2.INVTX1_2_.out
rlabel metal1 9522 27370 9522 27370 0 mux_bottom_ipin_2.INVTX1_3_.out
rlabel metal2 26174 25704 26174 25704 0 mux_bottom_ipin_2.INVTX1_4_.out
rlabel metal1 12696 22066 12696 22066 0 mux_bottom_ipin_2.INVTX1_5_.out
rlabel metal1 13662 32334 13662 32334 0 mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 12650 29614 12650 29614 0 mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 16790 34476 16790 34476 0 mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 14904 30022 14904 30022 0 mux_top_ipin_0.INVTX1_2_.out
rlabel metal2 24518 16592 24518 16592 0 mux_top_ipin_0.INVTX1_3_.out
rlabel metal1 24633 27370 24633 27370 0 mux_top_ipin_0.INVTX1_4_.out
rlabel metal1 18124 24786 18124 24786 0 mux_top_ipin_0.INVTX1_5_.out
rlabel metal2 14766 22814 14766 22814 0 mux_top_ipin_0.INVTX1_6_.out
rlabel metal1 15318 8602 15318 8602 0 mux_top_ipin_0.INVTX1_7_.out
rlabel metal1 14352 27982 14352 27982 0 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 15226 26112 15226 26112 0 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 9430 26418 9430 26418 0 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 6624 26282 6624 26282 0 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 10212 20026 10212 20026 0 mux_top_ipin_1.INVTX1_2_.out
rlabel metal1 13524 21658 13524 21658 0 mux_top_ipin_1.INVTX1_3_.out
rlabel metal1 12742 36006 12742 36006 0 mux_top_ipin_1.INVTX1_4_.out
rlabel metal1 7314 23834 7314 23834 0 mux_top_ipin_1.INVTX1_5_.out
rlabel metal1 21114 31790 21114 31790 0 mux_top_ipin_1.INVTX1_6_.out
rlabel metal1 9338 29070 9338 29070 0 mux_top_ipin_1.INVTX1_7_.out
rlabel metal2 15778 24514 15778 24514 0 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 12006 35054 12006 35054 0 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 13156 29682 13156 29682 0 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 16560 34408 16560 34408 0 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 14950 25024 14950 25024 0 mux_top_ipin_2.INVTX1_2_.out
rlabel metal1 11914 28424 11914 28424 0 mux_top_ipin_2.INVTX1_3_.out
rlabel metal1 12144 24242 12144 24242 0 mux_top_ipin_2.INVTX1_6_.out
rlabel metal1 14628 22474 14628 22474 0 mux_top_ipin_2.INVTX1_7_.out
rlabel metal1 14030 23596 14030 23596 0 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 13294 26656 13294 26656 0 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 13248 22950 13248 22950 0 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 35949 9554 35949 9554 0 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 15042 25738 15042 25738 0 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 15134 29036 15134 29036 0 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 16146 28594 16146 28594 0 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 23046 3060 23046 3060 0 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 36110 31892 36110 31892 0 net1
rlabel metal1 1886 29206 1886 29206 0 net10
rlabel metal2 36018 30158 36018 30158 0 net11
rlabel metal2 14490 2992 14490 2992 0 net12
rlabel metal2 35558 36890 35558 36890 0 net13
rlabel metal2 25898 27404 25898 27404 0 net14
rlabel metal2 6394 6833 6394 6833 0 net15
rlabel metal2 25346 30668 25346 30668 0 net16
rlabel metal1 14214 21862 14214 21862 0 net17
rlabel metal1 35788 2482 35788 2482 0 net18
rlabel metal1 21620 19822 21620 19822 0 net19
rlabel metal1 14306 36822 14306 36822 0 net2
rlabel metal1 36294 28050 36294 28050 0 net20
rlabel metal1 4094 9010 4094 9010 0 net21
rlabel metal1 2438 22610 2438 22610 0 net22
rlabel metal1 11362 2550 11362 2550 0 net23
rlabel metal2 32430 14484 32430 14484 0 net24
rlabel metal2 36202 10030 36202 10030 0 net25
rlabel metal1 36064 6426 36064 6426 0 net26
rlabel metal1 13800 3162 13800 3162 0 net27
rlabel metal1 2645 19822 2645 19822 0 net28
rlabel metal1 15364 6290 15364 6290 0 net29
rlabel metal2 15134 36618 15134 36618 0 net3
rlabel metal1 14076 36754 14076 36754 0 net30
rlabel metal2 35926 23392 35926 23392 0 net31
rlabel metal1 2162 25126 2162 25126 0 net32
rlabel metal1 31556 3026 31556 3026 0 net33
rlabel metal1 25760 16082 25760 16082 0 net34
rlabel metal1 2254 26962 2254 26962 0 net35
rlabel metal1 25208 14382 25208 14382 0 net36
rlabel metal2 15870 5440 15870 5440 0 net37
rlabel metal2 2530 3060 2530 3060 0 net38
rlabel metal1 22310 23698 22310 23698 0 net39
rlabel metal2 36110 24191 36110 24191 0 net4
rlabel metal1 13754 36346 13754 36346 0 net40
rlabel metal1 1886 19788 1886 19788 0 net41
rlabel metal2 35006 33660 35006 33660 0 net42
rlabel metal2 36110 8908 36110 8908 0 net43
rlabel metal2 24702 2652 24702 2652 0 net44
rlabel metal1 35834 24786 35834 24786 0 net45
rlabel metal2 5934 21913 5934 21913 0 net46
rlabel metal1 1932 22746 1932 22746 0 net47
rlabel metal1 35995 17170 35995 17170 0 net48
rlabel metal1 19458 37230 19458 37230 0 net49
rlabel metal1 1794 27982 1794 27982 0 net5
rlabel metal2 36110 6766 36110 6766 0 net50
rlabel metal1 29946 37162 29946 37162 0 net51
rlabel metal1 1886 3468 1886 3468 0 net52
rlabel metal1 2162 19686 2162 19686 0 net53
rlabel metal1 1886 2992 1886 2992 0 net54
rlabel metal2 18170 37060 18170 37060 0 net55
rlabel metal1 36156 23834 36156 23834 0 net56
rlabel metal1 2116 21522 2116 21522 0 net57
rlabel metal1 34040 3026 34040 3026 0 net58
rlabel metal2 25622 15776 25622 15776 0 net59
rlabel metal1 2898 4998 2898 4998 0 net6
rlabel metal1 3680 32878 3680 32878 0 net60
rlabel metal2 25070 8432 25070 8432 0 net61
rlabel metal1 15456 2822 15456 2822 0 net62
rlabel metal1 2116 3706 2116 3706 0 net63
rlabel metal1 28980 23494 28980 23494 0 net64
rlabel metal2 11730 37060 11730 37060 0 net65
rlabel metal1 19550 36550 19550 36550 0 net66
rlabel metal2 33626 30940 33626 30940 0 net67
rlabel metal2 1610 27404 1610 27404 0 net68
rlabel metal2 4646 2618 4646 2618 0 net69
rlabel via2 2530 18819 2530 18819 0 net7
rlabel metal1 1840 2414 1840 2414 0 net70
rlabel metal1 22218 22984 22218 22984 0 net71
rlabel metal1 28290 35258 28290 35258 0 net72
rlabel metal1 15732 2550 15732 2550 0 net73
rlabel metal2 35650 34374 35650 34374 0 net74
rlabel metal1 35995 3502 35995 3502 0 net75
rlabel metal1 5934 36754 5934 36754 0 net76
rlabel metal2 36018 23052 36018 23052 0 net77
rlabel metal2 6578 4522 6578 4522 0 net78
rlabel metal1 13156 14042 13156 14042 0 net79
rlabel metal1 13984 2550 13984 2550 0 net8
rlabel metal1 2323 16082 2323 16082 0 net80
rlabel metal2 36110 21862 36110 21862 0 net81
rlabel metal1 21022 19686 21022 19686 0 net82
rlabel metal1 31924 37230 31924 37230 0 net83
rlabel metal1 13018 36584 13018 36584 0 net84
rlabel metal1 25898 2482 25898 2482 0 net85
rlabel metal2 1886 12988 1886 12988 0 net86
rlabel metal2 17526 29342 17526 29342 0 net87
rlabel metal2 14766 21216 14766 21216 0 net88
rlabel metal1 16514 23834 16514 23834 0 net89
rlabel metal1 23138 31790 23138 31790 0 net9
rlabel metal2 13018 29852 13018 29852 0 net90
rlabel metal1 11454 23154 11454 23154 0 net91
rlabel metal1 17296 26418 17296 26418 0 net92
rlabel metal2 16974 34714 16974 34714 0 net93
rlabel metal1 30406 37264 30406 37264 0 pReset
rlabel metal1 1610 30260 1610 30260 0 prog_clk
rlabel metal2 7774 38056 7774 38056 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_
rlabel metal2 25162 1520 25162 1520 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_
rlabel metal3 1188 12308 1188 12308 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_
<< properties >>
string FIXED_BBOX 0 0 38000 40000
<< end >>
