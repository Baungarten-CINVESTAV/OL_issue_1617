// This is the unpowered netlist.
module cbx_1__4_ (bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_,
    bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_,
    bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_,
    bottom_grid_top_width_0_height_0_subtile_0__pin_clk_0_,
    ccff_head,
    ccff_tail,
    pReset,
    prog_clk,
    top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_,
    top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_,
    top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_,
    top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_,
    top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_,
    top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_,
    top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_,
    top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_,
    vccd1,
    vssd1,
    chanx_left_in,
    chanx_left_out,
    chanx_right_in,
    chanx_right_out);
 output bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
 output bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
 output bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
 output bottom_grid_top_width_0_height_0_subtile_0__pin_clk_0_;
 input ccff_head;
 output ccff_tail;
 input pReset;
 input prog_clk;
 output top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
 output top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
 output top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
 output top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
 output top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
 output top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
 output top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
 output top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
 inout vccd1;
 inout vssd1;
 input [0:18] chanx_left_in;
 output [0:18] chanx_left_out;
 input [0:18] chanx_right_in;
 output [0:18] chanx_right_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire clknet_0_prog_clk;
 wire \mem_bottom_ipin_0.DFFR_0_.Q ;
 wire \mem_bottom_ipin_0.DFFR_1_.Q ;
 wire \mem_bottom_ipin_0.DFFR_2_.Q ;
 wire \mem_bottom_ipin_0.DFFR_3_.Q ;
 wire \mem_bottom_ipin_0.DFFR_4_.Q ;
 wire \mem_bottom_ipin_0.DFFR_5_.Q ;
 wire \mem_bottom_ipin_1.DFFR_0_.Q ;
 wire \mem_bottom_ipin_1.DFFR_1_.Q ;
 wire \mem_bottom_ipin_1.DFFR_2_.Q ;
 wire \mem_bottom_ipin_1.DFFR_3_.Q ;
 wire \mem_bottom_ipin_1.DFFR_4_.Q ;
 wire \mem_bottom_ipin_1.DFFR_5_.Q ;
 wire \mem_bottom_ipin_2.DFFR_0_.Q ;
 wire \mem_bottom_ipin_2.DFFR_1_.Q ;
 wire \mem_bottom_ipin_2.DFFR_2_.Q ;
 wire \mem_bottom_ipin_2.DFFR_3_.Q ;
 wire \mem_bottom_ipin_2.DFFR_4_.Q ;
 wire \mem_bottom_ipin_2.DFFR_5_.Q ;
 wire \mem_bottom_ipin_3.DFFR_0_.Q ;
 wire \mem_bottom_ipin_3.DFFR_1_.Q ;
 wire \mem_bottom_ipin_3.DFFR_2_.Q ;
 wire \mem_bottom_ipin_3.DFFR_3_.Q ;
 wire \mem_bottom_ipin_3.DFFR_4_.Q ;
 wire \mem_bottom_ipin_3.DFFR_5_.Q ;
 wire \mem_bottom_ipin_4.DFFR_0_.Q ;
 wire \mem_bottom_ipin_4.DFFR_1_.Q ;
 wire \mem_bottom_ipin_4.DFFR_2_.Q ;
 wire \mem_bottom_ipin_4.DFFR_3_.Q ;
 wire \mem_bottom_ipin_4.DFFR_4_.Q ;
 wire \mem_bottom_ipin_4.DFFR_5_.Q ;
 wire \mem_bottom_ipin_5.DFFR_0_.Q ;
 wire \mem_bottom_ipin_5.DFFR_1_.Q ;
 wire \mem_bottom_ipin_5.DFFR_2_.Q ;
 wire \mem_bottom_ipin_5.DFFR_3_.Q ;
 wire \mem_bottom_ipin_5.DFFR_4_.Q ;
 wire \mem_bottom_ipin_5.DFFR_5_.Q ;
 wire \mem_bottom_ipin_6.DFFR_0_.Q ;
 wire \mem_bottom_ipin_6.DFFR_1_.Q ;
 wire \mem_bottom_ipin_6.DFFR_2_.Q ;
 wire \mem_bottom_ipin_6.DFFR_3_.Q ;
 wire \mem_bottom_ipin_6.DFFR_4_.Q ;
 wire \mem_bottom_ipin_6.DFFR_5_.Q ;
 wire \mem_bottom_ipin_7.DFFR_0_.Q ;
 wire \mem_bottom_ipin_7.DFFR_1_.Q ;
 wire \mem_bottom_ipin_7.DFFR_2_.Q ;
 wire \mem_bottom_ipin_7.DFFR_3_.Q ;
 wire \mem_bottom_ipin_7.DFFR_4_.Q ;
 wire \mem_bottom_ipin_7.DFFR_5_.Q ;
 wire \mem_top_ipin_0.DFFR_0_.Q ;
 wire \mem_top_ipin_0.DFFR_1_.Q ;
 wire \mem_top_ipin_0.DFFR_2_.Q ;
 wire \mem_top_ipin_0.DFFR_3_.Q ;
 wire \mem_top_ipin_0.DFFR_4_.Q ;
 wire \mem_top_ipin_0.DFFR_5_.Q ;
 wire \mem_top_ipin_1.DFFR_0_.Q ;
 wire \mem_top_ipin_1.DFFR_1_.Q ;
 wire \mem_top_ipin_1.DFFR_2_.Q ;
 wire \mem_top_ipin_1.DFFR_3_.Q ;
 wire \mem_top_ipin_1.DFFR_4_.Q ;
 wire \mem_top_ipin_1.DFFR_5_.Q ;
 wire \mem_top_ipin_2.DFFR_0_.Q ;
 wire \mem_top_ipin_2.DFFR_1_.Q ;
 wire \mem_top_ipin_2.DFFR_2_.Q ;
 wire \mem_top_ipin_2.DFFR_3_.Q ;
 wire \mem_top_ipin_2.DFFR_4_.Q ;
 wire \mem_top_ipin_2.DFFR_5_.Q ;
 wire \mem_top_ipin_3.DFFR_0_.Q ;
 wire \mem_top_ipin_3.DFFR_1_.Q ;
 wire \mem_top_ipin_3.DFFR_2_.Q ;
 wire \mem_top_ipin_3.DFFR_3_.Q ;
 wire \mem_top_ipin_3.DFFR_4_.Q ;
 wire \mux_bottom_ipin_0.INVTX1_0_.out ;
 wire \mux_bottom_ipin_0.INVTX1_1_.out ;
 wire \mux_bottom_ipin_0.INVTX1_2_.out ;
 wire \mux_bottom_ipin_0.INVTX1_3_.out ;
 wire \mux_bottom_ipin_0.INVTX1_4_.out ;
 wire \mux_bottom_ipin_0.INVTX1_5_.out ;
 wire \mux_bottom_ipin_0.INVTX1_6_.out ;
 wire \mux_bottom_ipin_0.INVTX1_7_.out ;
 wire \mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_bottom_ipin_1.INVTX1_2_.out ;
 wire \mux_bottom_ipin_1.INVTX1_3_.out ;
 wire \mux_bottom_ipin_1.INVTX1_4_.out ;
 wire \mux_bottom_ipin_1.INVTX1_5_.out ;
 wire \mux_bottom_ipin_1.INVTX1_6_.out ;
 wire \mux_bottom_ipin_1.INVTX1_7_.out ;
 wire \mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_bottom_ipin_2.INVTX1_2_.out ;
 wire \mux_bottom_ipin_2.INVTX1_3_.out ;
 wire \mux_bottom_ipin_2.INVTX1_4_.out ;
 wire \mux_bottom_ipin_2.INVTX1_5_.out ;
 wire \mux_bottom_ipin_2.INVTX1_6_.out ;
 wire \mux_bottom_ipin_2.INVTX1_7_.out ;
 wire \mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_bottom_ipin_3.INVTX1_2_.out ;
 wire \mux_bottom_ipin_3.INVTX1_3_.out ;
 wire \mux_bottom_ipin_3.INVTX1_4_.out ;
 wire \mux_bottom_ipin_3.INVTX1_5_.out ;
 wire \mux_bottom_ipin_3.INVTX1_6_.out ;
 wire \mux_bottom_ipin_3.INVTX1_7_.out ;
 wire \mux_bottom_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_bottom_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_bottom_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_bottom_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_bottom_ipin_4.INVTX1_2_.out ;
 wire \mux_bottom_ipin_4.INVTX1_3_.out ;
 wire \mux_bottom_ipin_4.INVTX1_4_.out ;
 wire \mux_bottom_ipin_4.INVTX1_5_.out ;
 wire \mux_bottom_ipin_4.INVTX1_6_.out ;
 wire \mux_bottom_ipin_4.INVTX1_7_.out ;
 wire \mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_bottom_ipin_5.INVTX1_2_.out ;
 wire \mux_bottom_ipin_5.INVTX1_3_.out ;
 wire \mux_bottom_ipin_5.INVTX1_4_.out ;
 wire \mux_bottom_ipin_5.INVTX1_5_.out ;
 wire \mux_bottom_ipin_5.INVTX1_6_.out ;
 wire \mux_bottom_ipin_5.INVTX1_7_.out ;
 wire \mux_bottom_ipin_5.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_bottom_ipin_5.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_bottom_ipin_5.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_bottom_ipin_5.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_bottom_ipin_6.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_bottom_ipin_6.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_bottom_ipin_6.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_bottom_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_bottom_ipin_7.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_bottom_ipin_7.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_bottom_ipin_7.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_bottom_ipin_7.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire clknet_3_0__leaf_prog_clk;
 wire clknet_3_1__leaf_prog_clk;
 wire clknet_3_2__leaf_prog_clk;
 wire clknet_3_3__leaf_prog_clk;
 wire clknet_3_4__leaf_prog_clk;
 wire clknet_3_5__leaf_prog_clk;
 wire clknet_3_6__leaf_prog_clk;
 wire clknet_3_7__leaf_prog_clk;

 sky130_fd_sc_hd__inv_2 _236_ (.A(_077_),
    .Y(_049_));
 sky130_fd_sc_hd__buf_4 _237_ (.A(_072_),
    .X(_078_));
 sky130_fd_sc_hd__inv_2 _238_ (.A(_078_),
    .Y(_050_));
 sky130_fd_sc_hd__inv_2 _239_ (.A(_078_),
    .Y(_051_));
 sky130_fd_sc_hd__inv_2 _240_ (.A(_078_),
    .Y(_052_));
 sky130_fd_sc_hd__inv_2 _241_ (.A(_078_),
    .Y(_053_));
 sky130_fd_sc_hd__inv_2 _242_ (.A(_078_),
    .Y(_054_));
 sky130_fd_sc_hd__inv_2 _243_ (.A(_078_),
    .Y(_055_));
 sky130_fd_sc_hd__inv_2 _244_ (.A(_078_),
    .Y(_056_));
 sky130_fd_sc_hd__inv_2 _245_ (.A(_078_),
    .Y(_057_));
 sky130_fd_sc_hd__inv_2 _246_ (.A(_078_),
    .Y(_058_));
 sky130_fd_sc_hd__inv_2 _247_ (.A(_078_),
    .Y(_059_));
 sky130_fd_sc_hd__buf_4 _248_ (.A(_072_),
    .X(_079_));
 sky130_fd_sc_hd__inv_2 _249_ (.A(_079_),
    .Y(_060_));
 sky130_fd_sc_hd__inv_2 _250_ (.A(_079_),
    .Y(_061_));
 sky130_fd_sc_hd__inv_2 _251_ (.A(_079_),
    .Y(_062_));
 sky130_fd_sc_hd__inv_2 _252_ (.A(_079_),
    .Y(_063_));
 sky130_fd_sc_hd__inv_2 _253_ (.A(_079_),
    .Y(_064_));
 sky130_fd_sc_hd__inv_2 _254_ (.A(_079_),
    .Y(_065_));
 sky130_fd_sc_hd__inv_2 _255_ (.A(_079_),
    .Y(_066_));
 sky130_fd_sc_hd__inv_2 _256_ (.A(_079_),
    .Y(_067_));
 sky130_fd_sc_hd__inv_2 _257_ (.A(_079_),
    .Y(_068_));
 sky130_fd_sc_hd__inv_2 _258_ (.A(_079_),
    .Y(_069_));
 sky130_fd_sc_hd__inv_2 _259_ (.A(_072_),
    .Y(_070_));
 sky130_fd_sc_hd__inv_2 _260_ (.A(_072_),
    .Y(_071_));
 sky130_fd_sc_hd__inv_2 _261_ (.A(\mem_top_ipin_3.DFFR_3_.Q ),
    .Y(_220_));
 sky130_fd_sc_hd__inv_2 _262_ (.A(\mem_top_ipin_3.DFFR_0_.Q ),
    .Y(_223_));
 sky130_fd_sc_hd__inv_2 _263_ (.A(\mem_top_ipin_3.DFFR_2_.Q ),
    .Y(_219_));
 sky130_fd_sc_hd__inv_2 _264_ (.A(\mem_top_ipin_3.DFFR_1_.Q ),
    .Y(_218_));
 sky130_fd_sc_hd__inv_2 _265_ (.A(net45),
    .Y(_213_));
 sky130_fd_sc_hd__inv_2 _266_ (.A(\mem_top_ipin_3.DFFR_0_.Q ),
    .Y(_221_));
 sky130_fd_sc_hd__inv_2 _267_ (.A(\mem_top_ipin_3.DFFR_2_.Q ),
    .Y(_215_));
 sky130_fd_sc_hd__inv_2 _268_ (.A(\mem_top_ipin_3.DFFR_1_.Q ),
    .Y(_214_));
 sky130_fd_sc_hd__inv_2 _269_ (.A(\mem_top_ipin_3.DFFR_4_.Q ),
    .Y(_212_));
 sky130_fd_sc_hd__inv_2 _270_ (.A(\mem_top_ipin_3.DFFR_0_.Q ),
    .Y(_222_));
 sky130_fd_sc_hd__inv_2 _271_ (.A(\mem_top_ipin_3.DFFR_2_.Q ),
    .Y(_217_));
 sky130_fd_sc_hd__inv_2 _272_ (.A(\mem_top_ipin_3.DFFR_1_.Q ),
    .Y(_216_));
 sky130_fd_sc_hd__inv_2 _273_ (.A(\mem_top_ipin_2.DFFR_3_.Q ),
    .Y(_208_));
 sky130_fd_sc_hd__inv_2 _274_ (.A(\mem_top_ipin_2.DFFR_0_.Q ),
    .Y(_211_));
 sky130_fd_sc_hd__inv_2 _275_ (.A(\mem_top_ipin_2.DFFR_2_.Q ),
    .Y(_207_));
 sky130_fd_sc_hd__inv_2 _276_ (.A(\mem_top_ipin_2.DFFR_1_.Q ),
    .Y(_206_));
 sky130_fd_sc_hd__inv_2 _277_ (.A(\mem_top_ipin_2.DFFR_5_.Q ),
    .Y(_201_));
 sky130_fd_sc_hd__inv_2 _278_ (.A(\mem_top_ipin_2.DFFR_0_.Q ),
    .Y(_209_));
 sky130_fd_sc_hd__inv_2 _279_ (.A(\mem_top_ipin_2.DFFR_2_.Q ),
    .Y(_203_));
 sky130_fd_sc_hd__inv_2 _280_ (.A(\mem_top_ipin_2.DFFR_1_.Q ),
    .Y(_202_));
 sky130_fd_sc_hd__inv_2 _281_ (.A(\mem_top_ipin_2.DFFR_4_.Q ),
    .Y(_200_));
 sky130_fd_sc_hd__inv_2 _282_ (.A(\mem_top_ipin_2.DFFR_0_.Q ),
    .Y(_210_));
 sky130_fd_sc_hd__inv_2 _283_ (.A(\mem_top_ipin_2.DFFR_2_.Q ),
    .Y(_205_));
 sky130_fd_sc_hd__inv_2 _284_ (.A(\mem_top_ipin_2.DFFR_1_.Q ),
    .Y(_204_));
 sky130_fd_sc_hd__inv_2 _285_ (.A(\mem_top_ipin_1.DFFR_3_.Q ),
    .Y(_196_));
 sky130_fd_sc_hd__inv_2 _286_ (.A(\mem_top_ipin_1.DFFR_0_.Q ),
    .Y(_199_));
 sky130_fd_sc_hd__inv_2 _287_ (.A(\mem_top_ipin_1.DFFR_2_.Q ),
    .Y(_195_));
 sky130_fd_sc_hd__inv_2 _288_ (.A(\mem_top_ipin_1.DFFR_1_.Q ),
    .Y(_194_));
 sky130_fd_sc_hd__inv_2 _289_ (.A(\mem_top_ipin_1.DFFR_5_.Q ),
    .Y(_189_));
 sky130_fd_sc_hd__inv_2 _290_ (.A(\mem_top_ipin_1.DFFR_0_.Q ),
    .Y(_197_));
 sky130_fd_sc_hd__inv_2 _291_ (.A(\mem_top_ipin_1.DFFR_2_.Q ),
    .Y(_191_));
 sky130_fd_sc_hd__inv_2 _292_ (.A(\mem_top_ipin_1.DFFR_1_.Q ),
    .Y(_190_));
 sky130_fd_sc_hd__inv_2 _293_ (.A(\mem_top_ipin_1.DFFR_4_.Q ),
    .Y(_188_));
 sky130_fd_sc_hd__inv_2 _294_ (.A(\mem_top_ipin_1.DFFR_0_.Q ),
    .Y(_198_));
 sky130_fd_sc_hd__inv_2 _295_ (.A(\mem_top_ipin_1.DFFR_2_.Q ),
    .Y(_193_));
 sky130_fd_sc_hd__inv_2 _296_ (.A(\mem_top_ipin_1.DFFR_1_.Q ),
    .Y(_192_));
 sky130_fd_sc_hd__inv_2 _297_ (.A(\mem_top_ipin_0.DFFR_3_.Q ),
    .Y(_184_));
 sky130_fd_sc_hd__inv_2 _298_ (.A(\mem_top_ipin_0.DFFR_0_.Q ),
    .Y(_187_));
 sky130_fd_sc_hd__inv_2 _299_ (.A(\mem_top_ipin_0.DFFR_2_.Q ),
    .Y(_183_));
 sky130_fd_sc_hd__inv_2 _300_ (.A(\mem_top_ipin_0.DFFR_1_.Q ),
    .Y(_182_));
 sky130_fd_sc_hd__inv_2 _301_ (.A(\mem_top_ipin_0.DFFR_5_.Q ),
    .Y(_177_));
 sky130_fd_sc_hd__inv_2 _302_ (.A(\mem_top_ipin_0.DFFR_0_.Q ),
    .Y(_185_));
 sky130_fd_sc_hd__inv_2 _303_ (.A(\mem_top_ipin_0.DFFR_2_.Q ),
    .Y(_179_));
 sky130_fd_sc_hd__inv_2 _304_ (.A(\mem_top_ipin_0.DFFR_1_.Q ),
    .Y(_178_));
 sky130_fd_sc_hd__inv_2 _305_ (.A(\mem_top_ipin_0.DFFR_4_.Q ),
    .Y(_176_));
 sky130_fd_sc_hd__inv_2 _306_ (.A(\mem_top_ipin_0.DFFR_0_.Q ),
    .Y(_186_));
 sky130_fd_sc_hd__inv_2 _307_ (.A(\mem_top_ipin_0.DFFR_2_.Q ),
    .Y(_181_));
 sky130_fd_sc_hd__inv_2 _308_ (.A(\mem_top_ipin_0.DFFR_1_.Q ),
    .Y(_180_));
 sky130_fd_sc_hd__inv_2 _309_ (.A(\mem_bottom_ipin_7.DFFR_3_.Q ),
    .Y(_172_));
 sky130_fd_sc_hd__inv_2 _310_ (.A(\mem_bottom_ipin_7.DFFR_0_.Q ),
    .Y(_175_));
 sky130_fd_sc_hd__inv_2 _311_ (.A(\mem_bottom_ipin_7.DFFR_2_.Q ),
    .Y(_171_));
 sky130_fd_sc_hd__inv_2 _312_ (.A(\mem_bottom_ipin_7.DFFR_1_.Q ),
    .Y(_170_));
 sky130_fd_sc_hd__inv_2 _313_ (.A(\mem_bottom_ipin_7.DFFR_5_.Q ),
    .Y(_165_));
 sky130_fd_sc_hd__inv_2 _314_ (.A(\mem_bottom_ipin_7.DFFR_0_.Q ),
    .Y(_173_));
 sky130_fd_sc_hd__inv_2 _315_ (.A(\mem_bottom_ipin_7.DFFR_2_.Q ),
    .Y(_167_));
 sky130_fd_sc_hd__inv_2 _316_ (.A(\mem_bottom_ipin_7.DFFR_1_.Q ),
    .Y(_166_));
 sky130_fd_sc_hd__inv_2 _317_ (.A(\mem_bottom_ipin_7.DFFR_4_.Q ),
    .Y(_164_));
 sky130_fd_sc_hd__inv_2 _318_ (.A(\mem_bottom_ipin_7.DFFR_0_.Q ),
    .Y(_174_));
 sky130_fd_sc_hd__inv_2 _319_ (.A(\mem_bottom_ipin_7.DFFR_2_.Q ),
    .Y(_169_));
 sky130_fd_sc_hd__inv_2 _320_ (.A(\mem_bottom_ipin_7.DFFR_1_.Q ),
    .Y(_168_));
 sky130_fd_sc_hd__inv_2 _321_ (.A(\mem_bottom_ipin_6.DFFR_3_.Q ),
    .Y(_160_));
 sky130_fd_sc_hd__inv_2 _322_ (.A(\mem_bottom_ipin_6.DFFR_0_.Q ),
    .Y(_163_));
 sky130_fd_sc_hd__inv_2 _323_ (.A(\mem_bottom_ipin_6.DFFR_2_.Q ),
    .Y(_159_));
 sky130_fd_sc_hd__inv_2 _324_ (.A(\mem_bottom_ipin_6.DFFR_1_.Q ),
    .Y(_158_));
 sky130_fd_sc_hd__inv_2 _325_ (.A(\mem_bottom_ipin_6.DFFR_5_.Q ),
    .Y(_153_));
 sky130_fd_sc_hd__inv_2 _326_ (.A(\mem_bottom_ipin_6.DFFR_0_.Q ),
    .Y(_161_));
 sky130_fd_sc_hd__inv_2 _327_ (.A(\mem_bottom_ipin_6.DFFR_2_.Q ),
    .Y(_155_));
 sky130_fd_sc_hd__inv_2 _328_ (.A(\mem_bottom_ipin_6.DFFR_1_.Q ),
    .Y(_154_));
 sky130_fd_sc_hd__inv_2 _329_ (.A(\mem_bottom_ipin_6.DFFR_4_.Q ),
    .Y(_152_));
 sky130_fd_sc_hd__inv_2 _330_ (.A(\mem_bottom_ipin_6.DFFR_0_.Q ),
    .Y(_162_));
 sky130_fd_sc_hd__inv_2 _331_ (.A(\mem_bottom_ipin_6.DFFR_2_.Q ),
    .Y(_157_));
 sky130_fd_sc_hd__inv_2 _332_ (.A(\mem_bottom_ipin_6.DFFR_1_.Q ),
    .Y(_156_));
 sky130_fd_sc_hd__inv_2 _333_ (.A(\mem_bottom_ipin_5.DFFR_3_.Q ),
    .Y(_148_));
 sky130_fd_sc_hd__inv_2 _334_ (.A(\mem_bottom_ipin_5.DFFR_0_.Q ),
    .Y(_151_));
 sky130_fd_sc_hd__inv_2 _335_ (.A(\mem_bottom_ipin_5.DFFR_2_.Q ),
    .Y(_147_));
 sky130_fd_sc_hd__inv_2 _336_ (.A(\mem_bottom_ipin_5.DFFR_1_.Q ),
    .Y(_146_));
 sky130_fd_sc_hd__inv_2 _337_ (.A(\mem_bottom_ipin_5.DFFR_5_.Q ),
    .Y(_141_));
 sky130_fd_sc_hd__inv_2 _338_ (.A(\mem_bottom_ipin_5.DFFR_0_.Q ),
    .Y(_149_));
 sky130_fd_sc_hd__inv_2 _339_ (.A(\mem_bottom_ipin_5.DFFR_2_.Q ),
    .Y(_143_));
 sky130_fd_sc_hd__inv_2 _340_ (.A(\mem_bottom_ipin_5.DFFR_1_.Q ),
    .Y(_142_));
 sky130_fd_sc_hd__inv_2 _341_ (.A(\mem_bottom_ipin_5.DFFR_4_.Q ),
    .Y(_140_));
 sky130_fd_sc_hd__inv_2 _342_ (.A(\mem_bottom_ipin_5.DFFR_0_.Q ),
    .Y(_150_));
 sky130_fd_sc_hd__inv_2 _343_ (.A(\mem_bottom_ipin_5.DFFR_2_.Q ),
    .Y(_145_));
 sky130_fd_sc_hd__inv_2 _344_ (.A(\mem_bottom_ipin_5.DFFR_1_.Q ),
    .Y(_144_));
 sky130_fd_sc_hd__inv_2 _345_ (.A(\mem_bottom_ipin_4.DFFR_3_.Q ),
    .Y(_136_));
 sky130_fd_sc_hd__inv_2 _346_ (.A(\mem_bottom_ipin_4.DFFR_0_.Q ),
    .Y(_139_));
 sky130_fd_sc_hd__inv_2 _347_ (.A(\mem_bottom_ipin_4.DFFR_2_.Q ),
    .Y(_135_));
 sky130_fd_sc_hd__inv_2 _348_ (.A(\mem_bottom_ipin_4.DFFR_1_.Q ),
    .Y(_134_));
 sky130_fd_sc_hd__inv_2 _349_ (.A(\mem_bottom_ipin_4.DFFR_5_.Q ),
    .Y(_129_));
 sky130_fd_sc_hd__inv_2 _350_ (.A(\mem_bottom_ipin_4.DFFR_0_.Q ),
    .Y(_137_));
 sky130_fd_sc_hd__inv_2 _351_ (.A(\mem_bottom_ipin_4.DFFR_2_.Q ),
    .Y(_131_));
 sky130_fd_sc_hd__inv_2 _352_ (.A(\mem_bottom_ipin_4.DFFR_1_.Q ),
    .Y(_130_));
 sky130_fd_sc_hd__inv_2 _353_ (.A(\mem_bottom_ipin_4.DFFR_4_.Q ),
    .Y(_128_));
 sky130_fd_sc_hd__inv_2 _354_ (.A(\mem_bottom_ipin_4.DFFR_0_.Q ),
    .Y(_138_));
 sky130_fd_sc_hd__inv_2 _355_ (.A(\mem_bottom_ipin_4.DFFR_2_.Q ),
    .Y(_133_));
 sky130_fd_sc_hd__inv_2 _356_ (.A(\mem_bottom_ipin_4.DFFR_1_.Q ),
    .Y(_132_));
 sky130_fd_sc_hd__inv_2 _357_ (.A(\mem_bottom_ipin_3.DFFR_3_.Q ),
    .Y(_124_));
 sky130_fd_sc_hd__inv_2 _358_ (.A(\mem_bottom_ipin_3.DFFR_0_.Q ),
    .Y(_127_));
 sky130_fd_sc_hd__inv_2 _359_ (.A(\mem_bottom_ipin_3.DFFR_2_.Q ),
    .Y(_123_));
 sky130_fd_sc_hd__inv_2 _360_ (.A(\mem_bottom_ipin_3.DFFR_1_.Q ),
    .Y(_122_));
 sky130_fd_sc_hd__inv_2 _361_ (.A(\mem_bottom_ipin_3.DFFR_5_.Q ),
    .Y(_117_));
 sky130_fd_sc_hd__inv_2 _362_ (.A(\mem_bottom_ipin_3.DFFR_0_.Q ),
    .Y(_125_));
 sky130_fd_sc_hd__inv_2 _363_ (.A(\mem_bottom_ipin_3.DFFR_2_.Q ),
    .Y(_119_));
 sky130_fd_sc_hd__inv_2 _364_ (.A(\mem_bottom_ipin_3.DFFR_1_.Q ),
    .Y(_118_));
 sky130_fd_sc_hd__inv_2 _365_ (.A(\mem_bottom_ipin_3.DFFR_4_.Q ),
    .Y(_116_));
 sky130_fd_sc_hd__inv_2 _366_ (.A(\mem_bottom_ipin_3.DFFR_0_.Q ),
    .Y(_126_));
 sky130_fd_sc_hd__inv_2 _367_ (.A(\mem_bottom_ipin_3.DFFR_2_.Q ),
    .Y(_121_));
 sky130_fd_sc_hd__inv_2 _368_ (.A(\mem_bottom_ipin_3.DFFR_1_.Q ),
    .Y(_120_));
 sky130_fd_sc_hd__inv_2 _369_ (.A(\mem_bottom_ipin_2.DFFR_3_.Q ),
    .Y(_112_));
 sky130_fd_sc_hd__inv_2 _370_ (.A(\mem_bottom_ipin_2.DFFR_0_.Q ),
    .Y(_115_));
 sky130_fd_sc_hd__inv_2 _371_ (.A(\mem_bottom_ipin_2.DFFR_2_.Q ),
    .Y(_111_));
 sky130_fd_sc_hd__inv_2 _372_ (.A(\mem_bottom_ipin_2.DFFR_1_.Q ),
    .Y(_110_));
 sky130_fd_sc_hd__inv_2 _373_ (.A(\mem_bottom_ipin_2.DFFR_5_.Q ),
    .Y(_105_));
 sky130_fd_sc_hd__inv_2 _374_ (.A(\mem_bottom_ipin_2.DFFR_0_.Q ),
    .Y(_113_));
 sky130_fd_sc_hd__inv_2 _375_ (.A(\mem_bottom_ipin_2.DFFR_2_.Q ),
    .Y(_107_));
 sky130_fd_sc_hd__inv_2 _376_ (.A(\mem_bottom_ipin_2.DFFR_1_.Q ),
    .Y(_106_));
 sky130_fd_sc_hd__inv_2 _377_ (.A(\mem_bottom_ipin_2.DFFR_4_.Q ),
    .Y(_104_));
 sky130_fd_sc_hd__inv_2 _378_ (.A(\mem_bottom_ipin_2.DFFR_0_.Q ),
    .Y(_114_));
 sky130_fd_sc_hd__inv_2 _379_ (.A(\mem_bottom_ipin_2.DFFR_2_.Q ),
    .Y(_109_));
 sky130_fd_sc_hd__inv_2 _380_ (.A(\mem_bottom_ipin_2.DFFR_1_.Q ),
    .Y(_108_));
 sky130_fd_sc_hd__inv_2 _381_ (.A(\mem_bottom_ipin_1.DFFR_3_.Q ),
    .Y(_100_));
 sky130_fd_sc_hd__inv_2 _382_ (.A(\mem_bottom_ipin_1.DFFR_0_.Q ),
    .Y(_103_));
 sky130_fd_sc_hd__inv_2 _383_ (.A(\mem_bottom_ipin_1.DFFR_1_.Q ),
    .Y(_099_));
 sky130_fd_sc_hd__inv_2 _384_ (.A(\mem_bottom_ipin_1.DFFR_2_.Q ),
    .Y(_098_));
 sky130_fd_sc_hd__inv_2 _385_ (.A(\mem_bottom_ipin_1.DFFR_4_.Q ),
    .Y(_097_));
 sky130_fd_sc_hd__inv_2 _386_ (.A(\mem_bottom_ipin_1.DFFR_0_.Q ),
    .Y(_102_));
 sky130_fd_sc_hd__inv_2 _387_ (.A(\mem_bottom_ipin_1.DFFR_1_.Q ),
    .Y(_095_));
 sky130_fd_sc_hd__inv_2 _388_ (.A(\mem_bottom_ipin_1.DFFR_2_.Q ),
    .Y(_094_));
 sky130_fd_sc_hd__inv_2 _389_ (.A(\mem_bottom_ipin_1.DFFR_5_.Q ),
    .Y(_092_));
 sky130_fd_sc_hd__inv_2 _390_ (.A(\mem_bottom_ipin_1.DFFR_0_.Q ),
    .Y(_101_));
 sky130_fd_sc_hd__inv_2 _391_ (.A(\mem_bottom_ipin_1.DFFR_2_.Q ),
    .Y(_096_));
 sky130_fd_sc_hd__inv_2 _392_ (.A(\mem_bottom_ipin_1.DFFR_1_.Q ),
    .Y(_093_));
 sky130_fd_sc_hd__inv_2 _393_ (.A(\mem_bottom_ipin_0.DFFR_3_.Q ),
    .Y(_091_));
 sky130_fd_sc_hd__inv_2 _394_ (.A(\mem_bottom_ipin_0.DFFR_0_.Q ),
    .Y(_088_));
 sky130_fd_sc_hd__inv_2 _395_ (.A(\mem_bottom_ipin_0.DFFR_4_.Q ),
    .Y(_087_));
 sky130_fd_sc_hd__inv_2 _396_ (.A(\mem_bottom_ipin_0.DFFR_0_.Q ),
    .Y(_089_));
 sky130_fd_sc_hd__inv_2 _397_ (.A(\mem_bottom_ipin_0.DFFR_5_.Q ),
    .Y(_086_));
 sky130_fd_sc_hd__inv_2 _398_ (.A(\mem_bottom_ipin_0.DFFR_0_.Q ),
    .Y(_090_));
 sky130_fd_sc_hd__inv_2 _399_ (.A(\mem_bottom_ipin_0.DFFR_1_.Q ),
    .Y(_085_));
 sky130_fd_sc_hd__inv_2 _400_ (.A(\mem_bottom_ipin_0.DFFR_2_.Q ),
    .Y(_084_));
 sky130_fd_sc_hd__inv_2 _401_ (.A(\mem_bottom_ipin_0.DFFR_1_.Q ),
    .Y(_083_));
 sky130_fd_sc_hd__inv_2 _402_ (.A(\mem_bottom_ipin_0.DFFR_2_.Q ),
    .Y(_082_));
 sky130_fd_sc_hd__inv_2 _403_ (.A(\mem_bottom_ipin_0.DFFR_1_.Q ),
    .Y(_081_));
 sky130_fd_sc_hd__inv_2 _404_ (.A(\mem_bottom_ipin_0.DFFR_2_.Q ),
    .Y(_080_));
 sky130_fd_sc_hd__inv_2 _405_ (.A(net5),
    .Y(\mux_bottom_ipin_0.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _406_ (.A(net24),
    .Y(\mux_bottom_ipin_0.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _407_ (.A(net11),
    .Y(\mux_bottom_ipin_0.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _408_ (.A(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net84));
 sky130_fd_sc_hd__inv_2 _409_ (.A(net30),
    .Y(\mux_bottom_ipin_0.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _410_ (.A(net2),
    .Y(\mux_bottom_ipin_0.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _411_ (.A(net21),
    .Y(\mux_bottom_ipin_0.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _412_ (.A(net17),
    .Y(\mux_bottom_ipin_0.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _413_ (.A(net36),
    .Y(\mux_bottom_ipin_0.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _414_ (.A(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net85));
 sky130_fd_sc_hd__inv_2 _415_ (.A(net37),
    .Y(\mux_bottom_ipin_1.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _416_ (.A(net18),
    .Y(\mux_bottom_ipin_1.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _417_ (.A(net6),
    .Y(\mux_bottom_ipin_1.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _418_ (.A(net31),
    .Y(\mux_bottom_ipin_1.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _419_ (.A(net12),
    .Y(\mux_bottom_ipin_1.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _420_ (.A(net25),
    .Y(\mux_bottom_ipin_1.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _421_ (.A(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net86));
 sky130_fd_sc_hd__inv_2 _422_ (.A(net7),
    .Y(\mux_bottom_ipin_2.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _423_ (.A(net38),
    .Y(\mux_bottom_ipin_2.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _424_ (.A(net19),
    .Y(\mux_bottom_ipin_2.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _425_ (.A(net32),
    .Y(\mux_bottom_ipin_2.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _426_ (.A(net13),
    .Y(\mux_bottom_ipin_2.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _427_ (.A(net26),
    .Y(\mux_bottom_ipin_2.INVTX1_7_.out ));
 sky130_fd_sc_hd__clkinv_2 _428_ (.A(\mux_bottom_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net87));
 sky130_fd_sc_hd__inv_2 _429_ (.A(net8),
    .Y(\mux_bottom_ipin_3.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _430_ (.A(net39),
    .Y(\mux_bottom_ipin_3.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _431_ (.A(net20),
    .Y(\mux_bottom_ipin_3.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _432_ (.A(net33),
    .Y(\mux_bottom_ipin_3.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _433_ (.A(net14),
    .Y(\mux_bottom_ipin_3.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _434_ (.A(net27),
    .Y(\mux_bottom_ipin_3.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _435_ (.A(\mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net88));
 sky130_fd_sc_hd__inv_2 _436_ (.A(net9),
    .Y(\mux_bottom_ipin_4.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _437_ (.A(net22),
    .Y(\mux_bottom_ipin_4.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _438_ (.A(net3),
    .Y(\mux_bottom_ipin_4.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _439_ (.A(net34),
    .Y(\mux_bottom_ipin_4.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _440_ (.A(net15),
    .Y(\mux_bottom_ipin_4.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _441_ (.A(net28),
    .Y(\mux_bottom_ipin_4.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _442_ (.A(\mux_bottom_ipin_5.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net89));
 sky130_fd_sc_hd__inv_2 _443_ (.A(net10),
    .Y(\mux_bottom_ipin_5.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _444_ (.A(net23),
    .Y(\mux_bottom_ipin_5.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _445_ (.A(net4),
    .Y(\mux_bottom_ipin_5.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _446_ (.A(net35),
    .Y(\mux_bottom_ipin_5.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _447_ (.A(net16),
    .Y(\mux_bottom_ipin_5.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _448_ (.A(net29),
    .Y(\mux_bottom_ipin_5.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _449_ (.A(\mux_bottom_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net90));
 sky130_fd_sc_hd__inv_2 _450_ (.A(\mux_bottom_ipin_7.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net91));
 sky130_fd_sc_hd__inv_2 _451_ (.A(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net41));
 sky130_fd_sc_hd__inv_2 _452_ (.A(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net42));
 sky130_fd_sc_hd__inv_2 _453_ (.A(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net43));
 sky130_fd_sc_hd__inv_2 _454_ (.A(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net44));
 sky130_fd_sc_hd__buf_2 _455_ (.A(net40),
    .X(_072_));
 sky130_fd_sc_hd__buf_4 _456_ (.A(_072_),
    .X(_073_));
 sky130_fd_sc_hd__inv_2 _457_ (.A(_073_),
    .Y(_000_));
 sky130_fd_sc_hd__inv_2 _458_ (.A(_073_),
    .Y(_001_));
 sky130_fd_sc_hd__inv_2 _459_ (.A(_073_),
    .Y(_002_));
 sky130_fd_sc_hd__inv_2 _460_ (.A(_073_),
    .Y(_003_));
 sky130_fd_sc_hd__inv_2 _461_ (.A(_073_),
    .Y(_004_));
 sky130_fd_sc_hd__inv_2 _462_ (.A(_073_),
    .Y(_005_));
 sky130_fd_sc_hd__inv_2 _463_ (.A(_073_),
    .Y(_006_));
 sky130_fd_sc_hd__inv_2 _464_ (.A(_073_),
    .Y(_007_));
 sky130_fd_sc_hd__inv_2 _465_ (.A(_073_),
    .Y(_008_));
 sky130_fd_sc_hd__inv_2 _466_ (.A(_073_),
    .Y(_009_));
 sky130_fd_sc_hd__buf_4 _467_ (.A(_072_),
    .X(_074_));
 sky130_fd_sc_hd__inv_2 _468_ (.A(_074_),
    .Y(_010_));
 sky130_fd_sc_hd__inv_2 _469_ (.A(_074_),
    .Y(_011_));
 sky130_fd_sc_hd__inv_2 _470_ (.A(_074_),
    .Y(_012_));
 sky130_fd_sc_hd__inv_2 _471_ (.A(_074_),
    .Y(_013_));
 sky130_fd_sc_hd__inv_2 _472_ (.A(_074_),
    .Y(_014_));
 sky130_fd_sc_hd__inv_2 _473_ (.A(_074_),
    .Y(_015_));
 sky130_fd_sc_hd__inv_2 _474_ (.A(_074_),
    .Y(_016_));
 sky130_fd_sc_hd__inv_2 _475_ (.A(_074_),
    .Y(_017_));
 sky130_fd_sc_hd__inv_2 _476_ (.A(_074_),
    .Y(_018_));
 sky130_fd_sc_hd__inv_2 _477_ (.A(_074_),
    .Y(_019_));
 sky130_fd_sc_hd__buf_4 _478_ (.A(_072_),
    .X(_075_));
 sky130_fd_sc_hd__inv_2 _479_ (.A(_075_),
    .Y(_020_));
 sky130_fd_sc_hd__inv_2 _480_ (.A(_075_),
    .Y(_021_));
 sky130_fd_sc_hd__inv_2 _481_ (.A(_075_),
    .Y(_022_));
 sky130_fd_sc_hd__inv_2 _482_ (.A(_075_),
    .Y(_023_));
 sky130_fd_sc_hd__inv_2 _483_ (.A(_075_),
    .Y(_024_));
 sky130_fd_sc_hd__inv_2 _484_ (.A(_075_),
    .Y(_025_));
 sky130_fd_sc_hd__inv_2 _485_ (.A(_075_),
    .Y(_026_));
 sky130_fd_sc_hd__inv_2 _486_ (.A(_075_),
    .Y(_027_));
 sky130_fd_sc_hd__inv_2 _487_ (.A(_075_),
    .Y(_028_));
 sky130_fd_sc_hd__inv_2 _488_ (.A(_075_),
    .Y(_029_));
 sky130_fd_sc_hd__buf_4 _489_ (.A(_072_),
    .X(_076_));
 sky130_fd_sc_hd__inv_2 _490_ (.A(_076_),
    .Y(_030_));
 sky130_fd_sc_hd__inv_2 _491_ (.A(_076_),
    .Y(_031_));
 sky130_fd_sc_hd__inv_2 _492_ (.A(_076_),
    .Y(_032_));
 sky130_fd_sc_hd__inv_2 _493_ (.A(_076_),
    .Y(_033_));
 sky130_fd_sc_hd__inv_2 _494_ (.A(_076_),
    .Y(_034_));
 sky130_fd_sc_hd__inv_2 _495_ (.A(_076_),
    .Y(_035_));
 sky130_fd_sc_hd__inv_2 _496_ (.A(_076_),
    .Y(_036_));
 sky130_fd_sc_hd__inv_2 _497_ (.A(_076_),
    .Y(_037_));
 sky130_fd_sc_hd__inv_2 _498_ (.A(_076_),
    .Y(_038_));
 sky130_fd_sc_hd__inv_2 _499_ (.A(_076_),
    .Y(_039_));
 sky130_fd_sc_hd__buf_4 _500_ (.A(_072_),
    .X(_077_));
 sky130_fd_sc_hd__inv_2 _501_ (.A(_077_),
    .Y(_040_));
 sky130_fd_sc_hd__inv_2 _502_ (.A(_077_),
    .Y(_041_));
 sky130_fd_sc_hd__inv_2 _503_ (.A(_077_),
    .Y(_042_));
 sky130_fd_sc_hd__inv_2 _504_ (.A(_077_),
    .Y(_043_));
 sky130_fd_sc_hd__inv_2 _505_ (.A(_077_),
    .Y(_044_));
 sky130_fd_sc_hd__inv_2 _506_ (.A(_077_),
    .Y(_045_));
 sky130_fd_sc_hd__inv_2 _507_ (.A(_077_),
    .Y(_046_));
 sky130_fd_sc_hd__inv_2 _508_ (.A(_077_),
    .Y(_047_));
 sky130_fd_sc_hd__inv_2 _509_ (.A(_077_),
    .Y(_048_));
 sky130_fd_sc_hd__dfrtp_1 _510_ (.CLK(clknet_3_1__leaf_prog_clk),
    .D(\mem_bottom_ipin_0.DFFR_4_.Q ),
    .RESET_B(_000_),
    .Q(\mem_bottom_ipin_0.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _511_ (.CLK(clknet_3_1__leaf_prog_clk),
    .D(\mem_bottom_ipin_0.DFFR_3_.Q ),
    .RESET_B(_001_),
    .Q(\mem_bottom_ipin_0.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _512_ (.CLK(clknet_3_2__leaf_prog_clk),
    .D(\mem_bottom_ipin_0.DFFR_2_.Q ),
    .RESET_B(_002_),
    .Q(\mem_bottom_ipin_0.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _513_ (.CLK(clknet_3_2__leaf_prog_clk),
    .D(\mem_bottom_ipin_0.DFFR_1_.Q ),
    .RESET_B(_003_),
    .Q(\mem_bottom_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _514_ (.CLK(clknet_3_3__leaf_prog_clk),
    .D(\mem_bottom_ipin_0.DFFR_0_.Q ),
    .RESET_B(_004_),
    .Q(\mem_bottom_ipin_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _515_ (.CLK(clknet_3_2__leaf_prog_clk),
    .D(net1),
    .RESET_B(_005_),
    .Q(\mem_bottom_ipin_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _516_ (.CLK(clknet_3_0__leaf_prog_clk),
    .D(\mem_bottom_ipin_1.DFFR_4_.Q ),
    .RESET_B(_006_),
    .Q(\mem_bottom_ipin_1.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _517_ (.CLK(clknet_3_0__leaf_prog_clk),
    .D(\mem_bottom_ipin_1.DFFR_3_.Q ),
    .RESET_B(_007_),
    .Q(\mem_bottom_ipin_1.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _518_ (.CLK(clknet_3_2__leaf_prog_clk),
    .D(\mem_bottom_ipin_1.DFFR_2_.Q ),
    .RESET_B(_008_),
    .Q(\mem_bottom_ipin_1.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _519_ (.CLK(clknet_3_6__leaf_prog_clk),
    .D(\mem_bottom_ipin_1.DFFR_1_.Q ),
    .RESET_B(_009_),
    .Q(\mem_bottom_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _520_ (.CLK(clknet_3_4__leaf_prog_clk),
    .D(\mem_bottom_ipin_1.DFFR_0_.Q ),
    .RESET_B(_010_),
    .Q(\mem_bottom_ipin_1.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _521_ (.CLK(clknet_3_2__leaf_prog_clk),
    .D(\mem_bottom_ipin_0.DFFR_5_.Q ),
    .RESET_B(_011_),
    .Q(\mem_bottom_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _522_ (.CLK(clknet_3_4__leaf_prog_clk),
    .D(\mem_bottom_ipin_2.DFFR_4_.Q ),
    .RESET_B(_012_),
    .Q(\mem_bottom_ipin_2.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _523_ (.CLK(clknet_3_5__leaf_prog_clk),
    .D(\mem_bottom_ipin_2.DFFR_3_.Q ),
    .RESET_B(_013_),
    .Q(\mem_bottom_ipin_2.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _524_ (.CLK(clknet_3_7__leaf_prog_clk),
    .D(\mem_bottom_ipin_2.DFFR_2_.Q ),
    .RESET_B(_014_),
    .Q(\mem_bottom_ipin_2.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _525_ (.CLK(clknet_3_7__leaf_prog_clk),
    .D(\mem_bottom_ipin_2.DFFR_1_.Q ),
    .RESET_B(_015_),
    .Q(\mem_bottom_ipin_2.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _526_ (.CLK(clknet_3_6__leaf_prog_clk),
    .D(\mem_bottom_ipin_2.DFFR_0_.Q ),
    .RESET_B(_016_),
    .Q(\mem_bottom_ipin_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _527_ (.CLK(clknet_3_1__leaf_prog_clk),
    .D(\mem_bottom_ipin_1.DFFR_5_.Q ),
    .RESET_B(_017_),
    .Q(\mem_bottom_ipin_2.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _528_ (.CLK(clknet_3_5__leaf_prog_clk),
    .D(\mem_bottom_ipin_3.DFFR_4_.Q ),
    .RESET_B(_018_),
    .Q(\mem_bottom_ipin_3.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _529_ (.CLK(clknet_3_6__leaf_prog_clk),
    .D(\mem_bottom_ipin_3.DFFR_3_.Q ),
    .RESET_B(_019_),
    .Q(\mem_bottom_ipin_3.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _530_ (.CLK(clknet_3_6__leaf_prog_clk),
    .D(\mem_bottom_ipin_3.DFFR_2_.Q ),
    .RESET_B(_020_),
    .Q(\mem_bottom_ipin_3.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _531_ (.CLK(clknet_3_7__leaf_prog_clk),
    .D(\mem_bottom_ipin_3.DFFR_1_.Q ),
    .RESET_B(_021_),
    .Q(\mem_bottom_ipin_3.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _532_ (.CLK(clknet_3_7__leaf_prog_clk),
    .D(\mem_bottom_ipin_3.DFFR_0_.Q ),
    .RESET_B(_022_),
    .Q(\mem_bottom_ipin_3.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _533_ (.CLK(clknet_3_6__leaf_prog_clk),
    .D(\mem_bottom_ipin_2.DFFR_5_.Q ),
    .RESET_B(_023_),
    .Q(\mem_bottom_ipin_3.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _534_ (.CLK(clknet_3_7__leaf_prog_clk),
    .D(\mem_bottom_ipin_4.DFFR_4_.Q ),
    .RESET_B(_024_),
    .Q(\mem_bottom_ipin_4.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _535_ (.CLK(clknet_3_5__leaf_prog_clk),
    .D(\mem_bottom_ipin_4.DFFR_3_.Q ),
    .RESET_B(_025_),
    .Q(\mem_bottom_ipin_4.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _536_ (.CLK(clknet_3_0__leaf_prog_clk),
    .D(\mem_bottom_ipin_4.DFFR_2_.Q ),
    .RESET_B(_026_),
    .Q(\mem_bottom_ipin_4.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _537_ (.CLK(clknet_3_6__leaf_prog_clk),
    .D(\mem_bottom_ipin_4.DFFR_1_.Q ),
    .RESET_B(_027_),
    .Q(\mem_bottom_ipin_4.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _538_ (.CLK(clknet_3_3__leaf_prog_clk),
    .D(\mem_bottom_ipin_4.DFFR_0_.Q ),
    .RESET_B(_028_),
    .Q(\mem_bottom_ipin_4.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _539_ (.CLK(clknet_3_6__leaf_prog_clk),
    .D(\mem_bottom_ipin_3.DFFR_5_.Q ),
    .RESET_B(_029_),
    .Q(\mem_bottom_ipin_4.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _540_ (.CLK(clknet_3_5__leaf_prog_clk),
    .D(\mem_bottom_ipin_5.DFFR_4_.Q ),
    .RESET_B(_030_),
    .Q(\mem_bottom_ipin_5.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _541_ (.CLK(clknet_3_5__leaf_prog_clk),
    .D(\mem_bottom_ipin_5.DFFR_3_.Q ),
    .RESET_B(_031_),
    .Q(\mem_bottom_ipin_5.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _542_ (.CLK(clknet_3_7__leaf_prog_clk),
    .D(\mem_bottom_ipin_5.DFFR_2_.Q ),
    .RESET_B(_032_),
    .Q(\mem_bottom_ipin_5.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _543_ (.CLK(clknet_3_4__leaf_prog_clk),
    .D(\mem_bottom_ipin_5.DFFR_1_.Q ),
    .RESET_B(_033_),
    .Q(\mem_bottom_ipin_5.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _544_ (.CLK(clknet_3_7__leaf_prog_clk),
    .D(\mem_bottom_ipin_5.DFFR_0_.Q ),
    .RESET_B(_034_),
    .Q(\mem_bottom_ipin_5.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _545_ (.CLK(clknet_3_4__leaf_prog_clk),
    .D(\mem_bottom_ipin_4.DFFR_5_.Q ),
    .RESET_B(_035_),
    .Q(\mem_bottom_ipin_5.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _546_ (.CLK(clknet_3_0__leaf_prog_clk),
    .D(\mem_bottom_ipin_6.DFFR_4_.Q ),
    .RESET_B(_036_),
    .Q(\mem_bottom_ipin_6.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _547_ (.CLK(clknet_3_0__leaf_prog_clk),
    .D(\mem_bottom_ipin_6.DFFR_3_.Q ),
    .RESET_B(_037_),
    .Q(\mem_bottom_ipin_6.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _548_ (.CLK(clknet_3_3__leaf_prog_clk),
    .D(\mem_bottom_ipin_6.DFFR_2_.Q ),
    .RESET_B(_038_),
    .Q(\mem_bottom_ipin_6.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _549_ (.CLK(clknet_3_2__leaf_prog_clk),
    .D(\mem_bottom_ipin_6.DFFR_1_.Q ),
    .RESET_B(_039_),
    .Q(\mem_bottom_ipin_6.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _550_ (.CLK(clknet_3_4__leaf_prog_clk),
    .D(\mem_bottom_ipin_6.DFFR_0_.Q ),
    .RESET_B(_040_),
    .Q(\mem_bottom_ipin_6.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _551_ (.CLK(clknet_3_5__leaf_prog_clk),
    .D(\mem_bottom_ipin_5.DFFR_5_.Q ),
    .RESET_B(_041_),
    .Q(\mem_bottom_ipin_6.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _552_ (.CLK(clknet_3_1__leaf_prog_clk),
    .D(\mem_bottom_ipin_7.DFFR_4_.Q ),
    .RESET_B(_042_),
    .Q(\mem_bottom_ipin_7.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _553_ (.CLK(clknet_3_3__leaf_prog_clk),
    .D(\mem_bottom_ipin_7.DFFR_3_.Q ),
    .RESET_B(_043_),
    .Q(\mem_bottom_ipin_7.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _554_ (.CLK(clknet_3_1__leaf_prog_clk),
    .D(\mem_bottom_ipin_7.DFFR_2_.Q ),
    .RESET_B(_044_),
    .Q(\mem_bottom_ipin_7.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _555_ (.CLK(clknet_3_4__leaf_prog_clk),
    .D(\mem_bottom_ipin_7.DFFR_1_.Q ),
    .RESET_B(_045_),
    .Q(\mem_bottom_ipin_7.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _556_ (.CLK(clknet_3_3__leaf_prog_clk),
    .D(\mem_bottom_ipin_7.DFFR_0_.Q ),
    .RESET_B(_046_),
    .Q(\mem_bottom_ipin_7.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _557_ (.CLK(clknet_3_3__leaf_prog_clk),
    .D(\mem_bottom_ipin_6.DFFR_5_.Q ),
    .RESET_B(_047_),
    .Q(\mem_bottom_ipin_7.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _558_ (.CLK(clknet_3_4__leaf_prog_clk),
    .D(\mem_top_ipin_0.DFFR_4_.Q ),
    .RESET_B(_048_),
    .Q(\mem_top_ipin_0.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _559_ (.CLK(clknet_3_1__leaf_prog_clk),
    .D(\mem_top_ipin_0.DFFR_3_.Q ),
    .RESET_B(_049_),
    .Q(\mem_top_ipin_0.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _560_ (.CLK(clknet_3_5__leaf_prog_clk),
    .D(\mem_top_ipin_0.DFFR_2_.Q ),
    .RESET_B(_050_),
    .Q(\mem_top_ipin_0.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _561_ (.CLK(clknet_3_7__leaf_prog_clk),
    .D(\mem_top_ipin_0.DFFR_1_.Q ),
    .RESET_B(_051_),
    .Q(\mem_top_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _562_ (.CLK(clknet_3_6__leaf_prog_clk),
    .D(\mem_top_ipin_0.DFFR_0_.Q ),
    .RESET_B(_052_),
    .Q(\mem_top_ipin_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _563_ (.CLK(clknet_3_4__leaf_prog_clk),
    .D(\mem_bottom_ipin_7.DFFR_5_.Q ),
    .RESET_B(_053_),
    .Q(\mem_top_ipin_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _564_ (.CLK(clknet_3_5__leaf_prog_clk),
    .D(\mem_top_ipin_1.DFFR_4_.Q ),
    .RESET_B(_054_),
    .Q(\mem_top_ipin_1.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _565_ (.CLK(clknet_3_4__leaf_prog_clk),
    .D(\mem_top_ipin_1.DFFR_3_.Q ),
    .RESET_B(_055_),
    .Q(\mem_top_ipin_1.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _566_ (.CLK(clknet_3_1__leaf_prog_clk),
    .D(\mem_top_ipin_1.DFFR_2_.Q ),
    .RESET_B(_056_),
    .Q(\mem_top_ipin_1.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _567_ (.CLK(clknet_3_3__leaf_prog_clk),
    .D(\mem_top_ipin_1.DFFR_1_.Q ),
    .RESET_B(_057_),
    .Q(\mem_top_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _568_ (.CLK(clknet_3_1__leaf_prog_clk),
    .D(\mem_top_ipin_1.DFFR_0_.Q ),
    .RESET_B(_058_),
    .Q(\mem_top_ipin_1.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _569_ (.CLK(clknet_3_5__leaf_prog_clk),
    .D(\mem_top_ipin_0.DFFR_5_.Q ),
    .RESET_B(_059_),
    .Q(\mem_top_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _570_ (.CLK(clknet_3_0__leaf_prog_clk),
    .D(\mem_top_ipin_2.DFFR_4_.Q ),
    .RESET_B(_060_),
    .Q(\mem_top_ipin_2.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _571_ (.CLK(clknet_3_0__leaf_prog_clk),
    .D(\mem_top_ipin_2.DFFR_3_.Q ),
    .RESET_B(_061_),
    .Q(\mem_top_ipin_2.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _572_ (.CLK(clknet_3_0__leaf_prog_clk),
    .D(\mem_top_ipin_2.DFFR_2_.Q ),
    .RESET_B(_062_),
    .Q(\mem_top_ipin_2.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _573_ (.CLK(clknet_3_2__leaf_prog_clk),
    .D(\mem_top_ipin_2.DFFR_1_.Q ),
    .RESET_B(_063_),
    .Q(\mem_top_ipin_2.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _574_ (.CLK(clknet_3_2__leaf_prog_clk),
    .D(\mem_top_ipin_2.DFFR_0_.Q ),
    .RESET_B(_064_),
    .Q(\mem_top_ipin_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _575_ (.CLK(clknet_3_3__leaf_prog_clk),
    .D(\mem_top_ipin_1.DFFR_5_.Q ),
    .RESET_B(_065_),
    .Q(\mem_top_ipin_2.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _576_ (.CLK(clknet_3_2__leaf_prog_clk),
    .D(\mem_top_ipin_3.DFFR_4_.Q ),
    .RESET_B(_066_),
    .Q(net45));
 sky130_fd_sc_hd__dfrtp_1 _577_ (.CLK(clknet_3_0__leaf_prog_clk),
    .D(\mem_top_ipin_3.DFFR_3_.Q ),
    .RESET_B(_067_),
    .Q(\mem_top_ipin_3.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _578_ (.CLK(clknet_3_2__leaf_prog_clk),
    .D(\mem_top_ipin_3.DFFR_2_.Q ),
    .RESET_B(_068_),
    .Q(\mem_top_ipin_3.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _579_ (.CLK(clknet_3_3__leaf_prog_clk),
    .D(\mem_top_ipin_3.DFFR_1_.Q ),
    .RESET_B(_069_),
    .Q(\mem_top_ipin_3.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _580_ (.CLK(clknet_3_0__leaf_prog_clk),
    .D(\mem_top_ipin_3.DFFR_0_.Q ),
    .RESET_B(_070_),
    .Q(\mem_top_ipin_3.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _581_ (.CLK(clknet_3_1__leaf_prog_clk),
    .D(\mem_top_ipin_2.DFFR_5_.Q ),
    .RESET_B(_071_),
    .Q(\mem_top_ipin_3.DFFR_0_.Q ));
 sky130_fd_sc_hd__conb_1 _648__93 (.HI(net93));
 sky130_fd_sc_hd__conb_1 _659__94 (.HI(net94));
 sky130_fd_sc_hd__conb_1 _671__95 (.HI(net95));
 sky130_fd_sc_hd__conb_1 _683__96 (.HI(net96));
 sky130_fd_sc_hd__conb_1 _695__97 (.HI(net97));
 sky130_fd_sc_hd__conb_1 _707__98 (.HI(net98));
 sky130_fd_sc_hd__conb_1 _719__99 (.HI(net99));
 sky130_fd_sc_hd__conb_1 _731__100 (.HI(net100));
 sky130_fd_sc_hd__conb_1 _743__101 (.HI(net101));
 sky130_fd_sc_hd__conb_1 _755__102 (.HI(net102));
 sky130_fd_sc_hd__conb_1 _767__103 (.HI(net103));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_prog_clk (.A(prog_clk),
    .X(clknet_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_1 _594_ (.A(net30),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 _595_ (.A(net29),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 _596_ (.A(net28),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 _597_ (.A(net27),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 _598_ (.A(net26),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 _599_ (.A(net25),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 _600_ (.A(net24),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 _601_ (.A(net23),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 _602_ (.A(net22),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 _603_ (.A(net39),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 _604_ (.A(net38),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 _605_ (.A(net37),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 _606_ (.A(net36),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 _607_ (.A(net35),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 _608_ (.A(net34),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 _609_ (.A(net33),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 _610_ (.A(net32),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 _611_ (.A(net31),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 _612_ (.A(net21),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 _613_ (.A(net11),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 _614_ (.A(net10),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 _615_ (.A(net9),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 _616_ (.A(net8),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 _617_ (.A(net7),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 _618_ (.A(net6),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 _619_ (.A(net5),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 _620_ (.A(net4),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 _621_ (.A(net3),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 _622_ (.A(net20),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 _623_ (.A(net19),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 _624_ (.A(net18),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 _625_ (.A(net17),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 _626_ (.A(net16),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 _627_ (.A(net15),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 _628_ (.A(net14),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 _629_ (.A(net13),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 _630_ (.A(net12),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 _631_ (.A(net2),
    .X(net65));
 sky130_fd_sc_hd__ebufn_2 _632_ (.A(\mux_bottom_ipin_0.INVTX1_2_.out ),
    .TE_B(_080_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _633_ (.A(\mux_bottom_ipin_0.INVTX1_1_.out ),
    .TE_B(_081_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _634_ (.A(\mux_bottom_ipin_0.INVTX1_5_.out ),
    .TE_B(_082_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _635_ (.A(\mux_bottom_ipin_0.INVTX1_4_.out ),
    .TE_B(_083_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _636_ (.A(net92),
    .TE_B(_084_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _637_ (.A(\mux_bottom_ipin_0.INVTX1_7_.out ),
    .TE_B(_085_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_4 _638_ (.A(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_086_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_4 _639_ (.A(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_087_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _640_ (.A(\mux_bottom_ipin_0.INVTX1_0_.out ),
    .TE_B(_088_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _641_ (.A(\mux_bottom_ipin_0.INVTX1_3_.out ),
    .TE_B(_089_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _642_ (.A(\mux_bottom_ipin_0.INVTX1_6_.out ),
    .TE_B(_090_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_4 _643_ (.A(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_091_),
    .Z(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _644_ (.A(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_092_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _645_ (.A(\mux_bottom_ipin_1.INVTX1_7_.out ),
    .TE_B(_093_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _646_ (.A(\mux_bottom_ipin_1.INVTX1_5_.out ),
    .TE_B(_094_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _647_ (.A(\mux_bottom_ipin_1.INVTX1_4_.out ),
    .TE_B(_095_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _648_ (.A(net93),
    .TE_B(_096_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _649_ (.A(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_097_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _650_ (.A(\mux_bottom_ipin_1.INVTX1_2_.out ),
    .TE_B(_098_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _651_ (.A(\mux_bottom_ipin_0.INVTX1_1_.out ),
    .TE_B(_099_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _652_ (.A(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_100_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _653_ (.A(\mux_bottom_ipin_1.INVTX1_6_.out ),
    .TE_B(_101_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _654_ (.A(\mux_bottom_ipin_1.INVTX1_3_.out ),
    .TE_B(_102_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _655_ (.A(\mux_bottom_ipin_0.INVTX1_0_.out ),
    .TE_B(_103_),
    .Z(\mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _656_ (.A(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_104_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _657_ (.A(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_105_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _658_ (.A(\mux_bottom_ipin_2.INVTX1_7_.out ),
    .TE_B(_106_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _659_ (.A(net94),
    .TE_B(_107_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _660_ (.A(\mux_bottom_ipin_2.INVTX1_4_.out ),
    .TE_B(_108_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _661_ (.A(\mux_bottom_ipin_2.INVTX1_5_.out ),
    .TE_B(_109_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_1 _662_ (.A(\mux_bottom_ipin_1.INVTX1_3_.out ),
    .TE_B(_110_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_1 _663_ (.A(\mux_bottom_ipin_2.INVTX1_2_.out ),
    .TE_B(_111_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _664_ (.A(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_112_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _665_ (.A(\mux_bottom_ipin_2.INVTX1_6_.out ),
    .TE_B(_113_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _666_ (.A(\mux_bottom_ipin_2.INVTX1_3_.out ),
    .TE_B(_114_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_1 _667_ (.A(\mux_bottom_ipin_1.INVTX1_2_.out ),
    .TE_B(_115_),
    .Z(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_4 _668_ (.A(\mux_bottom_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_116_),
    .Z(\mux_bottom_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_4 _669_ (.A(\mux_bottom_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_117_),
    .Z(\mux_bottom_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _670_ (.A(\mux_bottom_ipin_3.INVTX1_7_.out ),
    .TE_B(_118_),
    .Z(\mux_bottom_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _671_ (.A(net95),
    .TE_B(_119_),
    .Z(\mux_bottom_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _672_ (.A(\mux_bottom_ipin_3.INVTX1_4_.out ),
    .TE_B(_120_),
    .Z(\mux_bottom_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _673_ (.A(\mux_bottom_ipin_3.INVTX1_5_.out ),
    .TE_B(_121_),
    .Z(\mux_bottom_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _674_ (.A(\mux_bottom_ipin_2.INVTX1_3_.out ),
    .TE_B(_122_),
    .Z(\mux_bottom_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _675_ (.A(\mux_bottom_ipin_3.INVTX1_2_.out ),
    .TE_B(_123_),
    .Z(\mux_bottom_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_4 _676_ (.A(\mux_bottom_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_124_),
    .Z(\mux_bottom_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _677_ (.A(\mux_bottom_ipin_3.INVTX1_6_.out ),
    .TE_B(_125_),
    .Z(\mux_bottom_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _678_ (.A(\mux_bottom_ipin_3.INVTX1_3_.out ),
    .TE_B(_126_),
    .Z(\mux_bottom_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _679_ (.A(\mux_bottom_ipin_2.INVTX1_2_.out ),
    .TE_B(_127_),
    .Z(\mux_bottom_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _680_ (.A(\mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_128_),
    .Z(\mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _681_ (.A(\mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_129_),
    .Z(\mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _682_ (.A(\mux_bottom_ipin_4.INVTX1_7_.out ),
    .TE_B(_130_),
    .Z(\mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _683_ (.A(net96),
    .TE_B(_131_),
    .Z(\mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _684_ (.A(\mux_bottom_ipin_4.INVTX1_4_.out ),
    .TE_B(_132_),
    .Z(\mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _685_ (.A(\mux_bottom_ipin_4.INVTX1_5_.out ),
    .TE_B(_133_),
    .Z(\mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _686_ (.A(\mux_bottom_ipin_3.INVTX1_3_.out ),
    .TE_B(_134_),
    .Z(\mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _687_ (.A(\mux_bottom_ipin_4.INVTX1_2_.out ),
    .TE_B(_135_),
    .Z(\mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _688_ (.A(\mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_136_),
    .Z(\mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _689_ (.A(\mux_bottom_ipin_4.INVTX1_6_.out ),
    .TE_B(_137_),
    .Z(\mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _690_ (.A(\mux_bottom_ipin_4.INVTX1_3_.out ),
    .TE_B(_138_),
    .Z(\mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _691_ (.A(\mux_bottom_ipin_3.INVTX1_2_.out ),
    .TE_B(_139_),
    .Z(\mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _692_ (.A(\mux_bottom_ipin_5.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_140_),
    .Z(\mux_bottom_ipin_5.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _693_ (.A(\mux_bottom_ipin_5.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_141_),
    .Z(\mux_bottom_ipin_5.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _694_ (.A(\mux_bottom_ipin_5.INVTX1_7_.out ),
    .TE_B(_142_),
    .Z(\mux_bottom_ipin_5.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _695_ (.A(net97),
    .TE_B(_143_),
    .Z(\mux_bottom_ipin_5.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _696_ (.A(\mux_bottom_ipin_5.INVTX1_4_.out ),
    .TE_B(_144_),
    .Z(\mux_bottom_ipin_5.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _697_ (.A(\mux_bottom_ipin_5.INVTX1_5_.out ),
    .TE_B(_145_),
    .Z(\mux_bottom_ipin_5.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _698_ (.A(\mux_bottom_ipin_4.INVTX1_3_.out ),
    .TE_B(_146_),
    .Z(\mux_bottom_ipin_5.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _699_ (.A(\mux_bottom_ipin_5.INVTX1_2_.out ),
    .TE_B(_147_),
    .Z(\mux_bottom_ipin_5.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _700_ (.A(\mux_bottom_ipin_5.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_148_),
    .Z(\mux_bottom_ipin_5.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _701_ (.A(\mux_bottom_ipin_5.INVTX1_6_.out ),
    .TE_B(_149_),
    .Z(\mux_bottom_ipin_5.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _702_ (.A(\mux_bottom_ipin_5.INVTX1_3_.out ),
    .TE_B(_150_),
    .Z(\mux_bottom_ipin_5.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _703_ (.A(\mux_bottom_ipin_4.INVTX1_2_.out ),
    .TE_B(_151_),
    .Z(\mux_bottom_ipin_5.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _704_ (.A(\mux_bottom_ipin_6.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_152_),
    .Z(\mux_bottom_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _705_ (.A(\mux_bottom_ipin_6.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_153_),
    .Z(\mux_bottom_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _706_ (.A(\mux_bottom_ipin_0.INVTX1_7_.out ),
    .TE_B(_154_),
    .Z(\mux_bottom_ipin_6.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _707_ (.A(net98),
    .TE_B(_155_),
    .Z(\mux_bottom_ipin_6.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _708_ (.A(\mux_bottom_ipin_0.INVTX1_4_.out ),
    .TE_B(_156_),
    .Z(\mux_bottom_ipin_6.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _709_ (.A(\mux_bottom_ipin_0.INVTX1_5_.out ),
    .TE_B(_157_),
    .Z(\mux_bottom_ipin_6.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _710_ (.A(\mux_bottom_ipin_5.INVTX1_3_.out ),
    .TE_B(_158_),
    .Z(\mux_bottom_ipin_6.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _711_ (.A(\mux_bottom_ipin_0.INVTX1_2_.out ),
    .TE_B(_159_),
    .Z(\mux_bottom_ipin_6.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _712_ (.A(\mux_bottom_ipin_6.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_160_),
    .Z(\mux_bottom_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _713_ (.A(\mux_bottom_ipin_0.INVTX1_6_.out ),
    .TE_B(_161_),
    .Z(\mux_bottom_ipin_6.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _714_ (.A(\mux_bottom_ipin_0.INVTX1_3_.out ),
    .TE_B(_162_),
    .Z(\mux_bottom_ipin_6.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _715_ (.A(\mux_bottom_ipin_5.INVTX1_2_.out ),
    .TE_B(_163_),
    .Z(\mux_bottom_ipin_6.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _716_ (.A(\mux_bottom_ipin_7.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_164_),
    .Z(\mux_bottom_ipin_7.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _717_ (.A(\mux_bottom_ipin_7.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_165_),
    .Z(\mux_bottom_ipin_7.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _718_ (.A(\mux_bottom_ipin_1.INVTX1_7_.out ),
    .TE_B(_166_),
    .Z(\mux_bottom_ipin_7.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _719_ (.A(net99),
    .TE_B(_167_),
    .Z(\mux_bottom_ipin_7.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _720_ (.A(\mux_bottom_ipin_1.INVTX1_4_.out ),
    .TE_B(_168_),
    .Z(\mux_bottom_ipin_7.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _721_ (.A(\mux_bottom_ipin_1.INVTX1_5_.out ),
    .TE_B(_169_),
    .Z(\mux_bottom_ipin_7.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _722_ (.A(\mux_bottom_ipin_0.INVTX1_1_.out ),
    .TE_B(_170_),
    .Z(\mux_bottom_ipin_7.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _723_ (.A(\mux_bottom_ipin_0.INVTX1_2_.out ),
    .TE_B(_171_),
    .Z(\mux_bottom_ipin_7.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _724_ (.A(\mux_bottom_ipin_7.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_172_),
    .Z(\mux_bottom_ipin_7.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _725_ (.A(\mux_bottom_ipin_1.INVTX1_6_.out ),
    .TE_B(_173_),
    .Z(\mux_bottom_ipin_7.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _726_ (.A(\mux_bottom_ipin_0.INVTX1_3_.out ),
    .TE_B(_174_),
    .Z(\mux_bottom_ipin_7.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _727_ (.A(\mux_bottom_ipin_0.INVTX1_0_.out ),
    .TE_B(_175_),
    .Z(\mux_bottom_ipin_7.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _728_ (.A(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_176_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _729_ (.A(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_177_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _730_ (.A(\mux_bottom_ipin_2.INVTX1_7_.out ),
    .TE_B(_178_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _731_ (.A(net100),
    .TE_B(_179_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _732_ (.A(\mux_bottom_ipin_2.INVTX1_4_.out ),
    .TE_B(_180_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _733_ (.A(\mux_bottom_ipin_2.INVTX1_5_.out ),
    .TE_B(_181_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _734_ (.A(\mux_bottom_ipin_1.INVTX1_3_.out ),
    .TE_B(_182_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _735_ (.A(\mux_bottom_ipin_1.INVTX1_4_.out ),
    .TE_B(_183_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _736_ (.A(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_184_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _737_ (.A(\mux_bottom_ipin_2.INVTX1_6_.out ),
    .TE_B(_185_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _738_ (.A(\mux_bottom_ipin_1.INVTX1_5_.out ),
    .TE_B(_186_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _739_ (.A(\mux_bottom_ipin_1.INVTX1_2_.out ),
    .TE_B(_187_),
    .Z(\mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _740_ (.A(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_188_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _741_ (.A(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_189_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _742_ (.A(\mux_bottom_ipin_3.INVTX1_7_.out ),
    .TE_B(_190_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _743_ (.A(net101),
    .TE_B(_191_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _744_ (.A(\mux_bottom_ipin_3.INVTX1_4_.out ),
    .TE_B(_192_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _745_ (.A(\mux_bottom_ipin_3.INVTX1_5_.out ),
    .TE_B(_193_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _746_ (.A(\mux_bottom_ipin_2.INVTX1_3_.out ),
    .TE_B(_194_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _747_ (.A(\mux_bottom_ipin_2.INVTX1_4_.out ),
    .TE_B(_195_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _748_ (.A(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_196_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _749_ (.A(\mux_bottom_ipin_3.INVTX1_6_.out ),
    .TE_B(_197_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _750_ (.A(\mux_bottom_ipin_2.INVTX1_5_.out ),
    .TE_B(_198_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _751_ (.A(\mux_bottom_ipin_2.INVTX1_2_.out ),
    .TE_B(_199_),
    .Z(\mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _752_ (.A(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_200_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _753_ (.A(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_201_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _754_ (.A(\mux_bottom_ipin_4.INVTX1_7_.out ),
    .TE_B(_202_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _755_ (.A(net102),
    .TE_B(_203_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _756_ (.A(\mux_bottom_ipin_4.INVTX1_4_.out ),
    .TE_B(_204_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _757_ (.A(\mux_bottom_ipin_4.INVTX1_5_.out ),
    .TE_B(_205_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _758_ (.A(\mux_bottom_ipin_3.INVTX1_3_.out ),
    .TE_B(_206_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _759_ (.A(\mux_bottom_ipin_3.INVTX1_4_.out ),
    .TE_B(_207_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _760_ (.A(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_208_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _761_ (.A(\mux_bottom_ipin_4.INVTX1_6_.out ),
    .TE_B(_209_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _762_ (.A(\mux_bottom_ipin_3.INVTX1_5_.out ),
    .TE_B(_210_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _763_ (.A(\mux_bottom_ipin_3.INVTX1_2_.out ),
    .TE_B(_211_),
    .Z(\mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _764_ (.A(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_212_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _765_ (.A(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_213_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _766_ (.A(\mux_bottom_ipin_5.INVTX1_7_.out ),
    .TE_B(_214_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _767_ (.A(net103),
    .TE_B(_215_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _768_ (.A(\mux_bottom_ipin_5.INVTX1_4_.out ),
    .TE_B(_216_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _769_ (.A(\mux_bottom_ipin_5.INVTX1_5_.out ),
    .TE_B(_217_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _770_ (.A(\mux_bottom_ipin_4.INVTX1_3_.out ),
    .TE_B(_218_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _771_ (.A(\mux_bottom_ipin_4.INVTX1_4_.out ),
    .TE_B(_219_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _772_ (.A(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_220_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _773_ (.A(\mux_bottom_ipin_5.INVTX1_6_.out ),
    .TE_B(_221_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _774_ (.A(\mux_bottom_ipin_4.INVTX1_5_.out ),
    .TE_B(_222_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _775_ (.A(\mux_bottom_ipin_4.INVTX1_2_.out ),
    .TE_B(_223_),
    .Z(\mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(ccff_head),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(chanx_left_in[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(chanx_left_in[10]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(chanx_left_in[11]),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(chanx_left_in[12]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(chanx_left_in[13]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(chanx_left_in[14]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(chanx_left_in[15]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(chanx_left_in[16]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(chanx_left_in[17]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(chanx_left_in[18]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(chanx_left_in[1]),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(chanx_left_in[2]),
    .X(net13));
 sky130_fd_sc_hd__dlymetal6s2s_1 input14 (.A(chanx_left_in[3]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(chanx_left_in[4]),
    .X(net15));
 sky130_fd_sc_hd__dlymetal6s2s_1 input16 (.A(chanx_left_in[5]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(chanx_left_in[6]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(chanx_left_in[7]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(chanx_left_in[8]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(chanx_left_in[9]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(chanx_right_in[0]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(chanx_right_in[10]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(chanx_right_in[11]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(chanx_right_in[12]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(chanx_right_in[13]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(chanx_right_in[14]),
    .X(net26));
 sky130_fd_sc_hd__dlymetal6s2s_1 input27 (.A(chanx_right_in[15]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(chanx_right_in[16]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(chanx_right_in[17]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(chanx_right_in[18]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(chanx_right_in[1]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(chanx_right_in[2]),
    .X(net32));
 sky130_fd_sc_hd__dlymetal6s2s_1 input33 (.A(chanx_right_in[3]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(chanx_right_in[4]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(chanx_right_in[5]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(chanx_right_in[6]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(chanx_right_in[7]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(chanx_right_in[8]),
    .X(net38));
 sky130_fd_sc_hd__dlymetal6s2s_1 input39 (.A(chanx_right_in[9]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(pReset),
    .X(net40));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .X(bottom_grid_top_width_0_height_0_subtile_0__pin_clk_0_));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(ccff_tail));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .X(chanx_left_out[0]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .X(chanx_left_out[10]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(chanx_left_out[11]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .X(chanx_left_out[12]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .X(chanx_left_out[13]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(chanx_left_out[14]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .X(chanx_left_out[15]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(chanx_left_out[16]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net54),
    .X(chanx_left_out[17]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .X(chanx_left_out[18]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(chanx_left_out[1]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(chanx_left_out[2]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net58),
    .X(chanx_left_out[3]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(chanx_left_out[4]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(chanx_left_out[5]));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(chanx_left_out[6]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(chanx_left_out[7]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(chanx_left_out[8]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(chanx_left_out[9]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(chanx_right_out[0]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(chanx_right_out[10]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(chanx_right_out[11]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(chanx_right_out[12]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(chanx_right_out[13]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(chanx_right_out[14]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(chanx_right_out[15]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(chanx_right_out[16]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(chanx_right_out[17]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(chanx_right_out[18]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(chanx_right_out[1]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(chanx_right_out[2]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(chanx_right_out[3]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(chanx_right_out[4]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(chanx_right_out[5]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(chanx_right_out[6]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(chanx_right_out[7]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(chanx_right_out[8]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(chanx_right_out[9]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .X(top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_));
 sky130_fd_sc_hd__conb_1 _636__92 (.HI(net92));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_3_0__leaf_prog_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_3_1__leaf_prog_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_3_2__leaf_prog_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_3_3__leaf_prog_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_3_4__leaf_prog_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_3_5__leaf_prog_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_3_6__leaf_prog_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_3_7__leaf_prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__499__A (.DIODE(_076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__498__A (.DIODE(_076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__497__A (.DIODE(_076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__496__A (.DIODE(_076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__495__A (.DIODE(_076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__494__A (.DIODE(_076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__493__A (.DIODE(_076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__492__A (.DIODE(_076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__491__A (.DIODE(_076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__490__A (.DIODE(_076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__247__A (.DIODE(_078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__246__A (.DIODE(_078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__245__A (.DIODE(_078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__244__A (.DIODE(_078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__243__A (.DIODE(_078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__242__A (.DIODE(_078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__241__A (.DIODE(_078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__240__A (.DIODE(_078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__239__A (.DIODE(_078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__238__A (.DIODE(_078_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7__f_prog_clk_A (.DIODE(clknet_0_prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6__f_prog_clk_A (.DIODE(clknet_0_prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5__f_prog_clk_A (.DIODE(clknet_0_prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4__f_prog_clk_A (.DIODE(clknet_0_prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3__f_prog_clk_A (.DIODE(clknet_0_prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2__f_prog_clk_A (.DIODE(clknet_0_prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1__f_prog_clk_A (.DIODE(clknet_0_prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0__f_prog_clk_A (.DIODE(clknet_0_prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(ccff_head));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(chanx_left_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(chanx_left_in[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(chanx_left_in[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(chanx_left_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(chanx_left_in[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(chanx_left_in[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(chanx_left_in[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(chanx_left_in[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(chanx_left_in[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(chanx_left_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(chanx_left_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(chanx_left_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(chanx_left_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(chanx_left_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(chanx_left_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(chanx_left_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(chanx_left_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(chanx_left_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(chanx_left_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(chanx_right_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(chanx_right_in[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(chanx_right_in[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(chanx_right_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(chanx_right_in[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(chanx_right_in[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(chanx_right_in[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(chanx_right_in[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(chanx_right_in[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(chanx_right_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(chanx_right_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(chanx_right_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(chanx_right_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(chanx_right_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(chanx_right_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(chanx_right_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(chanx_right_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(chanx_right_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(chanx_right_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__514__D (.DIODE(\mem_bottom_ipin_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__398__A (.DIODE(\mem_bottom_ipin_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__396__A (.DIODE(\mem_bottom_ipin_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__394__A (.DIODE(\mem_bottom_ipin_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__512__D (.DIODE(\mem_bottom_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__404__A (.DIODE(\mem_bottom_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__402__A (.DIODE(\mem_bottom_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__400__A (.DIODE(\mem_bottom_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__520__D (.DIODE(\mem_bottom_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__390__A (.DIODE(\mem_bottom_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__386__A (.DIODE(\mem_bottom_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__382__A (.DIODE(\mem_bottom_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__518__D (.DIODE(\mem_bottom_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__391__A (.DIODE(\mem_bottom_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__388__A (.DIODE(\mem_bottom_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__384__A (.DIODE(\mem_bottom_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__527__D (.DIODE(\mem_bottom_ipin_1.DFFR_5_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__389__A (.DIODE(\mem_bottom_ipin_1.DFFR_5_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__526__D (.DIODE(\mem_bottom_ipin_2.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__378__A (.DIODE(\mem_bottom_ipin_2.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__374__A (.DIODE(\mem_bottom_ipin_2.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__370__A (.DIODE(\mem_bottom_ipin_2.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__530__D (.DIODE(\mem_bottom_ipin_3.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__367__A (.DIODE(\mem_bottom_ipin_3.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__363__A (.DIODE(\mem_bottom_ipin_3.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__359__A (.DIODE(\mem_bottom_ipin_3.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__538__D (.DIODE(\mem_bottom_ipin_4.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__354__A (.DIODE(\mem_bottom_ipin_4.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__350__A (.DIODE(\mem_bottom_ipin_4.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__346__A (.DIODE(\mem_bottom_ipin_4.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__537__D (.DIODE(\mem_bottom_ipin_4.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__356__A (.DIODE(\mem_bottom_ipin_4.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__352__A (.DIODE(\mem_bottom_ipin_4.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__348__A (.DIODE(\mem_bottom_ipin_4.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__536__D (.DIODE(\mem_bottom_ipin_4.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__355__A (.DIODE(\mem_bottom_ipin_4.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__351__A (.DIODE(\mem_bottom_ipin_4.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__347__A (.DIODE(\mem_bottom_ipin_4.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__544__D (.DIODE(\mem_bottom_ipin_5.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__342__A (.DIODE(\mem_bottom_ipin_5.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__338__A (.DIODE(\mem_bottom_ipin_5.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__334__A (.DIODE(\mem_bottom_ipin_5.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__543__D (.DIODE(\mem_bottom_ipin_5.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__344__A (.DIODE(\mem_bottom_ipin_5.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__340__A (.DIODE(\mem_bottom_ipin_5.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__336__A (.DIODE(\mem_bottom_ipin_5.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__542__D (.DIODE(\mem_bottom_ipin_5.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__343__A (.DIODE(\mem_bottom_ipin_5.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__339__A (.DIODE(\mem_bottom_ipin_5.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__335__A (.DIODE(\mem_bottom_ipin_5.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__550__D (.DIODE(\mem_bottom_ipin_6.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__330__A (.DIODE(\mem_bottom_ipin_6.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__326__A (.DIODE(\mem_bottom_ipin_6.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__322__A (.DIODE(\mem_bottom_ipin_6.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__549__D (.DIODE(\mem_bottom_ipin_6.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__332__A (.DIODE(\mem_bottom_ipin_6.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__328__A (.DIODE(\mem_bottom_ipin_6.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__324__A (.DIODE(\mem_bottom_ipin_6.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__555__D (.DIODE(\mem_bottom_ipin_7.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__320__A (.DIODE(\mem_bottom_ipin_7.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__316__A (.DIODE(\mem_bottom_ipin_7.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__312__A (.DIODE(\mem_bottom_ipin_7.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__568__D (.DIODE(\mem_top_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__294__A (.DIODE(\mem_top_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__290__A (.DIODE(\mem_top_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__286__A (.DIODE(\mem_top_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__567__D (.DIODE(\mem_top_ipin_1.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__296__A (.DIODE(\mem_top_ipin_1.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__292__A (.DIODE(\mem_top_ipin_1.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__288__A (.DIODE(\mem_top_ipin_1.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__566__D (.DIODE(\mem_top_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__295__A (.DIODE(\mem_top_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__291__A (.DIODE(\mem_top_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__287__A (.DIODE(\mem_top_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__574__D (.DIODE(\mem_top_ipin_2.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__282__A (.DIODE(\mem_top_ipin_2.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__278__A (.DIODE(\mem_top_ipin_2.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__274__A (.DIODE(\mem_top_ipin_2.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__573__D (.DIODE(\mem_top_ipin_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__284__A (.DIODE(\mem_top_ipin_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__280__A (.DIODE(\mem_top_ipin_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__276__A (.DIODE(\mem_top_ipin_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__572__D (.DIODE(\mem_top_ipin_2.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__283__A (.DIODE(\mem_top_ipin_2.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__279__A (.DIODE(\mem_top_ipin_2.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__275__A (.DIODE(\mem_top_ipin_2.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__580__D (.DIODE(\mem_top_ipin_3.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__270__A (.DIODE(\mem_top_ipin_3.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__266__A (.DIODE(\mem_top_ipin_3.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__262__A (.DIODE(\mem_top_ipin_3.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__579__D (.DIODE(\mem_top_ipin_3.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__272__A (.DIODE(\mem_top_ipin_3.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__268__A (.DIODE(\mem_top_ipin_3.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__264__A (.DIODE(\mem_top_ipin_3.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__408__A (.DIODE(\mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__746__A (.DIODE(\mux_bottom_ipin_2.INVTX1_3_.out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__674__A (.DIODE(\mux_bottom_ipin_2.INVTX1_3_.out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__666__A (.DIODE(\mux_bottom_ipin_2.INVTX1_3_.out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__421__A (.DIODE(\mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__428__A (.DIODE(\mux_bottom_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__688__A (.DIODE(\mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__680__A (.DIODE(\mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__681__A (.DIODE(\mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__693__A (.DIODE(\mux_bottom_ipin_5.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__712__A (.DIODE(\mux_bottom_ipin_6.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(pReset));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_prog_clk_A (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__515__D (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__631__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__410__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__621__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__438__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__620__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__445__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__619__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__405__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__616__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__429__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__615__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__436__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__630__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__419__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__629__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__426__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__628__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__433__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__627__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__440__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__625__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__412__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__624__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__416__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__623__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__424__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__622__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__431__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__612__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__411__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__602__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__437__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__601__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__444__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__600__A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__406__A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__599__A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__420__A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__596__A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__441__A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__595__A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__448__A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__611__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__418__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__609__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__432__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__608__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__439__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__607__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__446__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__606__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__413__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__604__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__423__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_output45_A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__265__A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_output46_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_output49_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_output50_A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_output56_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_output58_A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_output59_A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net83));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_384 ();
endmodule

