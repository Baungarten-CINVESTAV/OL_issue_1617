* NGSPICE file created from sb_4__0_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

.subckt sb_4__0_ ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11]
+ chanx_left_in[12] chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16]
+ chanx_left_in[17] chanx_left_in[18] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3]
+ chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8]
+ chanx_left_in[9] chanx_left_out[0] chanx_left_out[10] chanx_left_out[11] chanx_left_out[12]
+ chanx_left_out[13] chanx_left_out[14] chanx_left_out[15] chanx_left_out[16] chanx_left_out[17]
+ chanx_left_out[18] chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4]
+ chanx_left_out[5] chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_left_out[9]
+ chany_top_in[0] chany_top_in[10] chany_top_in[11] chany_top_in[12] chany_top_in[13]
+ chany_top_in[14] chany_top_in[15] chany_top_in[16] chany_top_in[17] chany_top_in[18]
+ chany_top_in[1] chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5]
+ chany_top_in[6] chany_top_in[7] chany_top_in[8] chany_top_in[9] chany_top_out[0]
+ chany_top_out[10] chany_top_out[11] chany_top_out[12] chany_top_out[13] chany_top_out[14]
+ chany_top_out[15] chany_top_out[16] chany_top_out[17] chany_top_out[18] chany_top_out[1]
+ chany_top_out[2] chany_top_out[3] chany_top_out[4] chany_top_out[5] chany_top_out[6]
+ chany_top_out[7] chany_top_out[8] chany_top_out[9] left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
+ left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_ left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
+ left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_ left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_
+ left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_ left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_
+ left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_ left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
+ left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_ pReset prog_clk top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_ top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
+ top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_ top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
+ top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_ top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_
+ top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_ top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_
+ top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_ vccd1 vssd1 vssd1_uq0
+ vccd1_uq0
XFILLER_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0419_ _0076_ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0770_ net20 vssd1 vssd1 vccd1 vccd1 mux_top_track_20.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XFILLER_5_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1184_ mux_top_track_24.mux_2level_tapbuf_basis_input2_mem1_0_out _0324_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input2_mem1_1_out sky130_fd_sc_hd__ebufn_1
XFILLER_20_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0899_ clknet_3_0__leaf_prog_clk mem_top_track_6.DFFR_1_.Q _0064_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_8.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0822_ _0176_ vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__inv_2
XFILLER_21_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0684_ _0165_ vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__clkbuf_1
X_0753_ net43 vssd1 vssd1 vccd1 vccd1 mux_left_track_11.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1236_ mux_left_track_35.mux_2level_tapbuf_basis_input2_mem1_0_out _0376_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_35.mux_2level_tapbuf_basis_input2_mem1_1_out sky130_fd_sc_hd__ebufn_2
XFILLER_64_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1098_ mux_top_track_16.INVTX1_1_.out _0238_ vssd1 vssd1 vccd1 vccd1 mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1167_ mux_left_track_19.INVTX1_0_.out _0307_ vssd1 vssd1 vccd1 vccd1 mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_12_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1178__123 vssd1 vssd1 vccd1 vccd1 net123 _1178__123/LO sky130_fd_sc_hd__conb_1
XFILLER_62_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1226__135 vssd1 vssd1 vccd1 vccd1 net135 _1226__135/LO sky130_fd_sc_hd__conb_1
XFILLER_34_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1021_ mux_left_track_3.out vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__clkbuf_1
X_0805_ net32 vssd1 vssd1 vccd1 vccd1 mux_left_track_35.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0736_ mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_2_out vssd1 vssd1 vccd1
+ vccd1 mux_top_track_18.out sky130_fd_sc_hd__inv_2
X_0598_ _0136_ vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__clkbuf_1
X_0667_ mem_top_track_10.DFFR_0_.D vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__inv_2
XFILLER_44_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1219_ mux_left_track_27.INVTX1_1_.out _0359_ vssd1 vssd1 vccd1 vccd1 mux_left_track_27.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0521_ mem_left_track_37.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_5 mux_top_track_34.INVTX1_1_.out vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0452_ mem_left_track_23.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__inv_2
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1004_ mux_left_track_37.out vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__clkbuf_1
X_0719_ mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_2_out vssd1 vssd1 vccd1
+ vccd1 mux_top_track_6.out sky130_fd_sc_hd__inv_2
XFILLER_57_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 chanx_left_out[11] sky130_fd_sc_hd__buf_2
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 chanx_left_out[4] sky130_fd_sc_hd__buf_2
XFILLER_63_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 chany_top_out[14] sky130_fd_sc_hd__buf_2
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 chany_top_out[7] sky130_fd_sc_hd__buf_2
XFILLER_31_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0504_ mem_top_track_22.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__clkbuf_1
X_0435_ mem_left_track_29.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__inv_2
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0418_ mem_left_track_35.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1183_ mux_top_track_24.INVTX1_1_.out _0323_ vssd1 vssd1 vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0898_ clknet_3_1__leaf_prog_clk mem_top_track_8.DFFR_0_.Q _0063_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_10.DFFR_0_.D sky130_fd_sc_hd__dfrtp_2
XFILLER_2_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0821_ _0176_ vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__inv_2
XFILLER_9_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0752_ mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_2_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_11.out sky130_fd_sc_hd__inv_2
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0683_ mem_top_track_6.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1235_ mux_left_track_15.INVTX1_2_.out _0375_ vssd1 vssd1 vccd1 vccd1 mux_left_track_35.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1166_ mux_left_track_17.INVTX1_2_.out _0306_ vssd1 vssd1 vccd1 vccd1 mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
X_1097_ net109 _0237_ vssd1 vssd1 vccd1 vccd1 mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_47_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1020_ mux_left_track_5.out vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__clkbuf_1
XFILLER_22_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0804_ mux_left_track_35.mux_2level_tapbuf_basis_input2_mem1_1_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_35.out sky130_fd_sc_hd__inv_2
X_0735_ net4 vssd1 vssd1 vccd1 vccd1 mux_top_track_16.INVTX1_2_.out sky130_fd_sc_hd__inv_2
XFILLER_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0666_ _0159_ vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__clkbuf_1
X_0597_ mem_left_track_3.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__clkbuf_1
X_1149_ mux_left_track_13.INVTX1_0_.out _0289_ vssd1 vssd1 vccd1 vccd1 mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_29_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1218_ net133 _0358_ vssd1 vssd1 vccd1 vccd1 mux_left_track_27.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_52_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0520_ mem_left_track_37.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__inv_2
XFILLER_3_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0451_ _0087_ vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0718_ net10 vssd1 vssd1 vccd1 vccd1 mux_top_track_4.INVTX1_2_.out sky130_fd_sc_hd__inv_2
XFILLER_57_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0649_ mem_top_track_12.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__inv_2
XFILLER_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 chany_top_out[8] sky130_fd_sc_hd__buf_2
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 chanx_left_out[5] sky130_fd_sc_hd__buf_2
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 chanx_left_out[12] sky130_fd_sc_hd__buf_2
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 chany_top_out[15] sky130_fd_sc_hd__buf_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0503_ mem_top_track_22.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__inv_2
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0434_ mem_left_track_29.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__inv_2
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0417_ mem_left_track_35.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__inv_2
XFILLER_35_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1182_ net124 _0322_ vssd1 vssd1 vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_32_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0897_ clknet_3_1__leaf_prog_clk mem_top_track_4.DFFR_1_.Q _0062_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_6.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0751_ net27 vssd1 vssd1 vccd1 vccd1 mux_left_track_9.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0820_ _0176_ vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__inv_2
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0682_ mem_top_track_6.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__inv_2
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1096_ mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_1_out _0236_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
X_1234_ net137 _0374_ vssd1 vssd1 vccd1 vccd1 mux_left_track_35.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1165_ mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_0_out _0305_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
XFILLER_20_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0949_ clknet_3_2__leaf_prog_clk mem_top_track_32.DFFR_1_.Q _0038_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_34.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0665_ mem_top_track_10.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__clkbuf_1
X_0734_ net60 vssd1 vssd1 vccd1 vccd1 mux_top_track_16.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_0803_ net33 vssd1 vssd1 vccd1 vccd1 mux_left_track_33.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0596_ mem_left_track_3.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__inv_2
XFILLER_52_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1217_ mux_left_track_25.INVTX1_0_.out _0357_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1148_ mux_left_track_13.INVTX1_2_.out _0288_ vssd1 vssd1 vccd1 vccd1 mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
X_1079_ net106 _0219_ vssd1 vssd1 vccd1 vccd1 mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0450_ mem_left_track_25.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0717_ mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_2_out vssd1 vssd1 vccd1
+ vccd1 mux_top_track_4.out sky130_fd_sc_hd__inv_2
X_0648_ _0153_ vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0579_ mem_left_track_7.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 chany_top_out[9] sky130_fd_sc_hd__buf_2
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 chanx_left_out[6] sky130_fd_sc_hd__buf_2
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 chany_top_out[16] sky130_fd_sc_hd__buf_2
XFILLER_0_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 chanx_left_out[13] sky130_fd_sc_hd__buf_2
XFILLER_63_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1198__128 vssd1 vssd1 vccd1 vccd1 net128 _1198__128/LO sky130_fd_sc_hd__conb_1
X_0502_ mem_top_track_22.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__inv_2
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0433_ _0081_ vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__clkbuf_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1061__103 vssd1 vssd1 vccd1 vccd1 net103 _1061__103/LO sky130_fd_sc_hd__conb_1
X_0416_ mem_left_track_35.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__inv_2
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1181_ mux_top_track_2.INVTX1_1_.out _0321_ vssd1 vssd1 vccd1 vccd1 mux_top_track_22.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0965_ clknet_3_4__leaf_prog_clk mem_left_track_33.DFFR_1_.Q _0054_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_35.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_1
X_0896_ clknet_3_0__leaf_prog_clk mem_top_track_6.DFFR_0_.Q _0061_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_6.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0681_ _0164_ vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__clkbuf_1
X_0750_ mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_2_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_9.out sky130_fd_sc_hd__inv_2
XFILLER_56_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1233_ mux_left_track_33.INVTX1_0_.out _0373_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1164_ mux_left_track_1.INVTX1_1_.out _0304_ vssd1 vssd1 vccd1 vccd1 mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1095_ mux_top_track_14.INVTX1_1_.out _0235_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_20_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0948_ clknet_3_7__leaf_prog_clk mem_top_track_34.DFFR_0_.Q _0037_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_34.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
X_0879_ _0181_ vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__inv_2
XFILLER_47_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0802_ mux_left_track_33.mux_2level_tapbuf_basis_input2_mem1_1_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_33.out sky130_fd_sc_hd__inv_2
X_0733_ mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_2_out vssd1 vssd1 vccd1
+ vccd1 mux_top_track_16.out sky130_fd_sc_hd__inv_2
X_0664_ mem_top_track_10.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__inv_2
XFILLER_37_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0595_ mem_left_track_3.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__inv_2
X_1216_ mux_left_track_25.mux_2level_tapbuf_basis_input2_mem1_0_out _0356_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input2_mem1_1_out sky130_fd_sc_hd__ebufn_2
XFILLER_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1147_ mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_0_out _0287_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_1
X_1078_ mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_1_out _0218_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0578_ mem_left_track_7.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__inv_2
X_0716_ net11 vssd1 vssd1 vccd1 vccd1 mux_top_track_2.INVTX1_2_.out sky130_fd_sc_hd__inv_2
X_0647_ mem_top_track_14.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 chanx_left_out[7] sky130_fd_sc_hd__buf_2
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 chanx_left_out[14] sky130_fd_sc_hd__buf_2
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 chany_top_out[17] sky130_fd_sc_hd__buf_2
XFILLER_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0432_ mem_left_track_31.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__clkbuf_1
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0501_ _0104_ vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1091__108 vssd1 vssd1 vccd1 vccd1 net108 _1091__108/LO sky130_fd_sc_hd__conb_1
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1180_ mux_top_track_22.mux_2level_tapbuf_basis_input2_mem1_0_out _0320_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_22.mux_2level_tapbuf_basis_input2_mem1_1_out sky130_fd_sc_hd__ebufn_2
XFILLER_32_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0964_ clknet_3_4__leaf_prog_clk mem_left_track_35.DFFR_0_.Q _0053_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_35.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_2
X_0895_ clknet_3_6__leaf_prog_clk mem_top_track_2.DFFR_1_.Q _0060_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_4.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0680_ mem_top_track_6.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__clkbuf_1
X_1232_ mux_left_track_33.mux_2level_tapbuf_basis_input2_mem1_0_out _0372_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input2_mem1_1_out sky130_fd_sc_hd__ebufn_2
XFILLER_1_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1094_ mux_top_track_16.INVTX1_2_.out _0234_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
X_1163_ net120 _0303_ vssd1 vssd1 vccd1 vccd1 mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_20_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0947_ clknet_3_0__leaf_prog_clk mem_top_track_30.DFFR_1_.Q _0036_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_32.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0878_ _0181_ vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__inv_2
XFILLER_43_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0801_ net34 vssd1 vssd1 vccd1 vccd1 mux_left_track_31.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0594_ _0135_ vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0663_ _0158_ vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__clkbuf_1
X_0732_ net5 vssd1 vssd1 vccd1 vccd1 mux_top_track_14.INVTX1_2_.out sky130_fd_sc_hd__inv_2
X_1146_ mux_left_track_11.INVTX1_2_.out _0286_ vssd1 vssd1 vccd1 vccd1 mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1215_ mux_left_track_25.INVTX1_1_.out _0355_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_25_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1077_ mux_top_track_10.INVTX1_0_.out _0217_ vssd1 vssd1 vccd1 vccd1 mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_25_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0715_ mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_2_out vssd1 vssd1 vccd1
+ vccd1 mux_top_track_2.out sky130_fd_sc_hd__inv_2
X_0577_ mem_left_track_7.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__inv_2
X_0646_ mem_top_track_14.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__inv_2
X_1129_ mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_0_out _0269_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 chanx_left_out[15] sky130_fd_sc_hd__buf_2
XFILLER_56_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 chanx_left_out[8] sky130_fd_sc_hd__buf_2
XFILLER_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0431_ _0080_ vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__clkbuf_1
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0500_ mem_top_track_24.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0629_ mem_top_track_18.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0963_ clknet_3_5__leaf_prog_clk mem_left_track_31.DFFR_1_.Q _0052_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_33.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_1
X_0894_ clknet_3_1__leaf_prog_clk mem_top_track_4.DFFR_0_.Q _0059_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_4.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_2
XFILLER_4_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1231_ mux_left_track_13.INVTX1_2_.out _0371_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1162_ mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_1_out _0302_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
XFILLER_64_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1093_ mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_0_out _0233_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
XFILLER_20_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0946_ clknet_3_0__leaf_prog_clk mem_top_track_32.DFFR_0_.Q _0035_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_32.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_2
X_0877_ _0181_ vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__inv_2
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1115__112 vssd1 vssd1 vccd1 vccd1 net112 _1115__112/LO sky130_fd_sc_hd__conb_1
XFILLER_18_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0800_ mux_left_track_31.mux_2level_tapbuf_basis_input2_mem1_1_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_31.out sky130_fd_sc_hd__inv_2
X_0731_ net59 vssd1 vssd1 vccd1 vccd1 mux_top_track_14.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_0593_ mem_left_track_5.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0662_ mem_top_track_10.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1145_ net117 _0285_ vssd1 vssd1 vccd1 vccd1 mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_25_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1214_ net132 _0354_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1076_ mux_top_track_10.INVTX1_2_.out _0216_ vssd1 vssd1 vccd1 vccd1 mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
X_0929_ clknet_3_7__leaf_prog_clk mem_left_track_15.DFFR_1_.Q _0018_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_17.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_48 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0714_ net53 vssd1 vssd1 vccd1 vccd1 mux_top_track_2.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_0645_ _0152_ vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__clkbuf_1
X_0576_ _0129_ vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__clkbuf_1
X_1128_ mux_left_track_25.INVTX1_1_.out _0268_ vssd1 vssd1 vccd1 vccd1 mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1059_ mux_top_track_2.INVTX1_1_.out _0199_ vssd1 vssd1 vccd1 vccd1 mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 chanx_left_out[16] sky130_fd_sc_hd__buf_2
XFILLER_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0430_ mem_left_track_31.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__clkbuf_1
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0628_ mem_top_track_18.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__inv_2
XFILLER_26_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0559_ mem_left_track_11.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__inv_2
XFILLER_13_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0962_ clknet_3_5__leaf_prog_clk mem_left_track_33.DFFR_0_.Q _0051_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_33.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
X_0893_ clknet_3_6__leaf_prog_clk mem_top_track_0.DFFR_1_.Q _0058_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_2.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_2
XFILLER_4_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1230_ net136 _0370_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1092_ mux_top_track_16.INVTX1_1_.out _0232_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1161_ mux_left_track_17.INVTX1_0_.out _0301_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_20_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0945_ clknet_3_0__leaf_prog_clk mem_top_track_28.DFFR_1_.Q _0034_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_30.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_2
X_0876_ _0181_ vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__inv_2
XFILLER_9_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0661_ _0157_ vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__clkbuf_1
X_0730_ mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_2_out vssd1 vssd1 vccd1
+ vccd1 mux_top_track_14.out sky130_fd_sc_hd__inv_2
XFILLER_10_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0592_ mem_left_track_5.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__inv_2
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1213_ mux_left_track_23.INVTX1_0_.out _0353_ vssd1 vssd1 vccd1 vccd1 mux_left_track_23.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1144_ mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_1_out _0284_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_1
XFILLER_37_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1075_ mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_0_out _0215_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
XFILLER_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1145__117 vssd1 vssd1 vccd1 vccd1 net117 _1145__117/LO sky130_fd_sc_hd__conb_1
XFILLER_33_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0859_ _0179_ vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__inv_2
X_0928_ clknet_3_3__leaf_prog_clk mem_left_track_17.DFFR_0_.Q _0017_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_17.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0713_ net2 vssd1 vssd1 vccd1 vccd1 mux_top_track_0.INVTX1_2_.out sky130_fd_sc_hd__inv_2
X_0644_ mem_top_track_14.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__clkbuf_1
X_0575_ mem_left_track_9.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__clkbuf_1
X_1058_ mux_top_track_4.INVTX1_2_.out _0198_ vssd1 vssd1 vccd1 vccd1 mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
X_1127_ net114 _0267_ vssd1 vssd1 vccd1 vccd1 mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_25_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0558_ _0123_ vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__clkbuf_1
X_0627_ _0146_ vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0489_ _0100_ vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0961_ clknet_3_5__leaf_prog_clk mem_left_track_29.DFFR_1_.Q _0050_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_31.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_2
XFILLER_17_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0892_ clknet_3_6__leaf_prog_clk mem_top_track_2.DFFR_0_.Q _0057_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_2.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_55_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1091_ net108 _0231_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
X_1160_ mux_left_track_17.INVTX1_2_.out _0300_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0944_ clknet_3_2__leaf_prog_clk mem_top_track_30.DFFR_0_.Q _0033_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_30.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
X_0875_ _0181_ vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__inv_2
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0591_ _0134_ vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__clkbuf_1
X_0660_ mem_top_track_10.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1212_ mux_left_track_23.mux_2level_tapbuf_basis_input2_mem1_0_out _0352_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_23.mux_2level_tapbuf_basis_input2_mem1_1_out sky130_fd_sc_hd__ebufn_2
X_1074_ mux_top_track_10.INVTX1_1_.out _0214_ vssd1 vssd1 vccd1 vccd1 mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_1_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1143_ mux_left_track_11.INVTX1_0_.out _0283_ vssd1 vssd1 vccd1 vccd1 mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0927_ clknet_3_4__leaf_prog_clk mem_left_track_13.DFFR_1_.Q _0016_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_15.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
X_0789_ mux_left_track_23.mux_2level_tapbuf_basis_input2_mem1_1_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_23.out sky130_fd_sc_hd__inv_2
X_0858_ _0179_ vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__inv_2
XFILLER_28_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0712_ mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_2_out vssd1 vssd1 vccd1
+ vccd1 mux_top_track_0.out sky130_fd_sc_hd__inv_2
X_0643_ _0151_ vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__clkbuf_1
X_0574_ mem_left_track_9.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__inv_2
X_1126_ mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_1_out _0266_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
XFILLER_33_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1057_ mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_0_out _0197_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
XFILLER_15_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1174__122 vssd1 vssd1 vccd1 vccd1 net122 _1174__122/LO sky130_fd_sc_hd__conb_1
XFILLER_62_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1222__134 vssd1 vssd1 vccd1 vccd1 net134 _1222__134/LO sky130_fd_sc_hd__conb_1
XFILLER_7_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0557_ mem_left_track_13.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__clkbuf_1
X_0626_ mem_top_track_18.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__clkbuf_1
X_0488_ mem_top_track_28.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__clkbuf_1
X_1109_ net111 _0249_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0609_ _0140_ vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0960_ clknet_3_5__leaf_prog_clk mem_left_track_31.DFFR_0_.Q _0049_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_31.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_2
X_0891_ clknet_3_7__leaf_prog_clk net1 _0056_ vssd1 vssd1 vccd1 vccd1 mem_top_track_0.DFFR_0_.Q
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_4_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1090_ mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_1_out _0230_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
XFILLER_20_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0943_ clknet_3_5__leaf_prog_clk mem_top_track_26.DFFR_1_.Q _0032_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_28.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_2
X_0874_ _0181_ vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__inv_2
XFILLER_9_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0590_ mem_left_track_5.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1142_ mux_left_track_11.INVTX1_2_.out _0282_ vssd1 vssd1 vccd1 vccd1 mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
X_1211_ mux_left_track_23.INVTX1_1_.out _0351_ vssd1 vssd1 vccd1 vccd1 mux_left_track_23.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1073_ net105 _0213_ vssd1 vssd1 vccd1 vccd1 mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
X_0926_ clknet_3_4__leaf_prog_clk mem_left_track_15.DFFR_0_.Q _0015_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_15.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_2
X_0857_ _0179_ vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__inv_2
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0788_ net39 vssd1 vssd1 vccd1 vccd1 mux_left_track_21.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_56_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0711_ net52 vssd1 vssd1 vccd1 vccd1 mux_top_track_0.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0573_ _0128_ vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__clkbuf_1
X_0642_ mem_top_track_14.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__clkbuf_1
X_1125_ mux_left_track_5.INVTX1_0_.out _0265_ vssd1 vssd1 vccd1 vccd1 mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_38_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1056_ mux_top_track_24.INVTX1_0_.out _0196_ vssd1 vssd1 vccd1 vccd1 mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_0909_ clknet_3_0__leaf_prog_clk mem_top_track_16.DFFR_1_.Q _0074_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_18.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_48_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0625_ _0145_ vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0487_ _0099_ vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__clkbuf_1
X_0556_ mem_left_track_13.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__inv_2
XFILLER_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1039_ mux_top_track_4.out vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__clkbuf_1
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1108_ mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_1_out _0248_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
XFILLER_44_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0608_ mem_left_track_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__clkbuf_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0539_ mem_left_track_17.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0890_ clknet_3_6__leaf_prog_clk mem_top_track_0.DFFR_0_.Q _0055_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_0.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_55_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1067__104 vssd1 vssd1 vccd1 vccd1 net104 _1067__104/LO sky130_fd_sc_hd__conb_1
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0873_ net50 vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__buf_4
X_0942_ clknet_3_5__leaf_prog_clk mem_top_track_28.DFFR_0_.Q _0031_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_28.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_2
XFILLER_9_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1072_ mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_1_out _0212_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
XFILLER_1_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1210_ net131 _0350_ vssd1 vssd1 vccd1 vccd1 mux_left_track_23.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1141_ mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_0_out _0281_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
XFILLER_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0787_ mux_left_track_21.mux_2level_tapbuf_basis_input2_mem1_1_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_21.out sky130_fd_sc_hd__inv_2
X_0856_ _0179_ vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__inv_2
X_0925_ clknet_3_3__leaf_prog_clk mem_left_track_11.DFFR_1_.Q _0014_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_13.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0710_ net51 vssd1 vssd1 vccd1 vccd1 mux_top_track_0.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0641_ mem_top_track_14.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__inv_2
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0572_ mem_left_track_11.DFFR_0_.D vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1124_ mux_left_track_25.INVTX1_1_.out _0264_ vssd1 vssd1 vccd1 vccd1 mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
X_1055_ net102 _0195_ vssd1 vssd1 vccd1 vccd1 mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_33_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0908_ clknet_3_4__leaf_prog_clk mem_top_track_18.DFFR_0_.Q _0073_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_18.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0839_ _0177_ vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__inv_2
XFILLER_56_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0624_ mem_top_track_18.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0145_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0555_ _0122_ vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__clkbuf_1
X_0486_ mem_top_track_28.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__clkbuf_1
X_1038_ mux_top_track_6.out vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__clkbuf_1
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1107_ mux_top_track_0.INVTX1_0_.out _0247_ vssd1 vssd1 vccd1 vccd1 mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0538_ mem_left_track_17.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__inv_2
X_0607_ _0139_ vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0469_ _0093_ vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1194__127 vssd1 vssd1 vccd1 vccd1 net127 _1194__127/LO sky130_fd_sc_hd__conb_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0941_ clknet_3_7__leaf_prog_clk mem_top_track_24.DFFR_1_.Q _0030_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_26.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0872_ _0180_ vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__inv_2
XFILLER_9_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1097__109 vssd1 vssd1 vccd1 vccd1 net109 _1097__109/LO sky130_fd_sc_hd__conb_1
XFILLER_24_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1071_ mux_top_track_26.INVTX1_0_.out _0211_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_1_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1140_ mux_left_track_11.INVTX1_1_.out _0280_ vssd1 vssd1 vccd1 vccd1 mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0924_ clknet_3_5__leaf_prog_clk mem_left_track_13.DFFR_0_.Q _0013_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_13.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_2
X_0855_ _0179_ vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__inv_2
X_0786_ net13 vssd1 vssd1 vccd1 vccd1 mux_top_track_34.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XFILLER_28_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0571_ _0127_ vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__clkbuf_1
X_0640_ mem_top_track_14.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__inv_2
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1123_ mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_0_out _0263_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
X_1054_ mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_1_out _0194_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
XFILLER_18_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0907_ clknet_3_2__leaf_prog_clk mem_top_track_14.DFFR_1_.Q _0072_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_16.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_2
X_0838_ _0177_ vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__inv_2
X_0769_ mux_top_track_20.mux_2level_tapbuf_basis_input2_mem1_1_out vssd1 vssd1 vccd1
+ vccd1 mux_top_track_20.out sky130_fd_sc_hd__inv_2
XFILLER_56_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0554_ mem_left_track_13.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__clkbuf_1
X_0623_ mem_top_track_18.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__inv_2
XFILLER_7_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0485_ mem_top_track_28.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__inv_2
X_1106_ mux_top_track_36.INVTX1_2_.out _0246_ vssd1 vssd1 vccd1 vccd1 mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1037_ mux_top_track_8.out vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0606_ mem_left_track_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__clkbuf_1
X_0537_ _0116_ vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__clkbuf_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0468_ mem_top_track_34.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0940_ clknet_3_5__leaf_prog_clk mem_top_track_26.DFFR_0_.Q _0029_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_26.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_13_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0871_ _0180_ vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__inv_2
XFILLER_9_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1070_ mux_top_track_8.INVTX1_2_.out _0210_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0854_ _0179_ vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__inv_2
X_0923_ clknet_3_3__leaf_prog_clk mem_left_track_11.DFFR_0_.D _0012_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_11.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
X_0785_ mux_top_track_34.mux_2level_tapbuf_basis_input2_mem1_1_out vssd1 vssd1 vccd1
+ vccd1 mux_top_track_34.out sky130_fd_sc_hd__inv_2
XFILLER_61_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1199_ mux_top_track_32.INVTX1_1_.out _0339_ vssd1 vssd1 vccd1 vccd1 mux_top_track_32.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_24_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0570_ mem_left_track_9.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__clkbuf_1
X_1122_ mux_left_track_23.INVTX1_1_.out _0262_ vssd1 vssd1 vccd1 vccd1 mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1053_ mux_top_track_0.INVTX1_1_.out _0193_ vssd1 vssd1 vccd1 vccd1 mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_0906_ clknet_3_0__leaf_prog_clk mem_top_track_16.DFFR_0_.Q _0071_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_16.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
X_0837_ _0177_ vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__inv_2
X_0699_ mem_top_track_2.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__clkbuf_1
X_0768_ net31 vssd1 vssd1 vccd1 vccd1 mux_left_track_37.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_56_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0553_ _0121_ vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__clkbuf_1
X_0484_ mem_top_track_28.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__inv_2
X_0622_ mem_top_track_18.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__inv_2
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1105_ mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_0_out _0245_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1036_ mux_top_track_10.out vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0605_ mem_left_track_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__inv_2
X_0467_ mem_top_track_34.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__inv_2
X_0536_ mem_left_track_17.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__clkbuf_1
X_1019_ mux_left_track_7.out vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__clkbuf_1
XFILLER_26_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0519_ _0110_ vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__clkbuf_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0870_ _0180_ vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__inv_2
XFILLER_9_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0853_ _0179_ vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__inv_2
X_0922_ clknet_3_3__leaf_prog_clk mem_left_track_11.DFFR_0_.Q _0011_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_11.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
X_0784_ net14 vssd1 vssd1 vccd1 vccd1 mux_top_track_32.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_1198_ net128 _0338_ vssd1 vssd1 vccd1 vccd1 mux_top_track_32.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_2
Xinput1 ccff_head vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0_prog_clk prog_clk vssd1 vssd1 vccd1 vccd1 clknet_0_prog_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_59_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1121_ net113 _0261_ vssd1 vssd1 vccd1 vccd1 mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
X_1052_ mux_top_track_2.INVTX1_2_.out _0192_ vssd1 vssd1 vccd1 vccd1 mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_33_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0836_ _0177_ vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__inv_2
X_0905_ clknet_3_3__leaf_prog_clk mem_top_track_12.DFFR_1_.Q _0070_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_14.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
X_0767_ mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_2_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_37.out sky130_fd_sc_hd__inv_2
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0698_ mem_top_track_2.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__inv_2
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0621_ _0144_ vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0552_ mem_left_track_13.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0483_ _0098_ vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1104_ mux_top_track_16.INVTX1_1_.out _0244_ vssd1 vssd1 vccd1 vccd1 mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1035_ mux_top_track_12.out vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__clkbuf_1
XFILLER_61_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0819_ _0176_ vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__inv_2
XFILLER_29_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0604_ mem_left_track_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__inv_2
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0535_ _0115_ vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__clkbuf_1
X_0466_ mem_top_track_34.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__inv_2
XFILLER_41_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1018_ mux_left_track_9.out vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0518_ net61 vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__clkbuf_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0449_ _0086_ vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__clkbuf_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1218__133 vssd1 vssd1 vccd1 vccd1 net133 _1218__133/LO sky130_fd_sc_hd__conb_1
XFILLER_18_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0921_ clknet_3_6__leaf_prog_clk mem_left_track_7.DFFR_1_.Q _0010_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_9.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_18_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0783_ mux_top_track_32.mux_2level_tapbuf_basis_input2_mem1_1_out vssd1 vssd1 vccd1
+ vccd1 mux_top_track_32.out sky130_fd_sc_hd__inv_2
X_1121__113 vssd1 vssd1 vccd1 vccd1 net113 _1121__113/LO sky130_fd_sc_hd__conb_1
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0852_ _0179_ vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__inv_2
XFILLER_5_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput2 chanx_left_in[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1197_ mux_top_track_10.INVTX1_1_.out _0337_ vssd1 vssd1 vccd1 vccd1 mux_top_track_30.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_3_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1120_ mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_1_out _0260_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1051_ mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_0_out _0191_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
XFILLER_18_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0904_ clknet_3_2__leaf_prog_clk mem_top_track_14.DFFR_0_.Q _0069_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_14.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
X_0766_ net22 vssd1 vssd1 vccd1 vccd1 mux_left_track_19.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0697_ _0169_ vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__clkbuf_1
X_0835_ _0177_ vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__inv_2
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0551_ mem_left_track_13.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__inv_2
X_0620_ mem_top_track_36.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0482_ mem_top_track_30.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1103_ net110 _0243_ vssd1 vssd1 vccd1 vccd1 mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_21_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1034_ mux_top_track_14.out vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__clkbuf_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0749_ net28 vssd1 vssd1 vccd1 vccd1 mux_left_track_7.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0818_ _0174_ vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__buf_4
Xinput60 top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0603_ _0138_ vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__clkbuf_1
X_0534_ mem_left_track_17.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0465_ _0092_ vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1017_ mux_left_track_11.out vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0517_ _0109_ vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__clkbuf_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0448_ mem_left_track_25.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__clkbuf_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0920_ clknet_3_3__leaf_prog_clk mem_left_track_9.DFFR_0_.Q _0009_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_11.DFFR_0_.D sky130_fd_sc_hd__dfrtp_1
X_0782_ net15 vssd1 vssd1 vccd1 vccd1 mux_top_track_30.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_0851_ net50 vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__buf_4
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput3 chanx_left_in[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1196_ mux_top_track_30.mux_2level_tapbuf_basis_input2_mem1_0_out _0336_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_30.mux_2level_tapbuf_basis_input2_mem1_1_out sky130_fd_sc_hd__ebufn_2
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1151__118 vssd1 vssd1 vccd1 vccd1 net118 _1151__118/LO sky130_fd_sc_hd__conb_1
X_1050_ mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_1_out _0190_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
XFILLER_18_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0903_ clknet_3_1__leaf_prog_clk mem_top_track_10.DFFR_1_.Q _0068_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_12.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_14_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0834_ _0177_ vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__inv_2
X_0696_ mem_top_track_2.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__clkbuf_1
X_0765_ mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_2_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_19.out sky130_fd_sc_hd__inv_2
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1179_ mux_top_track_22.INVTX1_1_.out _0319_ vssd1 vssd1 vccd1 vccd1 mux_top_track_22.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_24_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0550_ mem_left_track_13.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__inv_2
XFILLER_7_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1102_ mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_1_out _0242_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
X_0481_ _0097_ vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__clkbuf_1
XFILLER_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1033_ mux_top_track_16.out vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__clkbuf_1
Xinput50 pReset vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_2
X_0817_ _0175_ vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__inv_2
X_0748_ mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_2_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_7.out sky130_fd_sc_hd__inv_2
X_0679_ _0163_ vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0533_ mem_left_track_17.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__inv_2
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0464_ mem_left_track_21.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__clkbuf_1
X_0602_ mem_left_track_3.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__clkbuf_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1016_ mux_left_track_13.out vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__clkbuf_1
XFILLER_34_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0447_ mem_left_track_25.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__inv_2
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0516_ mem_left_track_37.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__clkbuf_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0850_ _0178_ vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__inv_2
X_0781_ mux_top_track_30.mux_2level_tapbuf_basis_input2_mem1_1_out vssd1 vssd1 vccd1
+ vccd1 mux_top_track_30.out sky130_fd_sc_hd__inv_2
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput4 chanx_left_in[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1195_ mux_top_track_30.INVTX1_1_.out _0335_ vssd1 vssd1 vccd1 vccd1 mux_top_track_30.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0833_ _0177_ vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__inv_2
X_0902_ clknet_3_0__leaf_prog_clk mem_top_track_12.DFFR_0_.Q _0067_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_12.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_14_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0764_ net47 vssd1 vssd1 vccd1 vccd1 mux_left_track_17.INVTX1_2_.out sky130_fd_sc_hd__inv_2
X_0695_ mem_top_track_2.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__inv_2
X_1178_ net123 _0318_ vssd1 vssd1 vccd1 vccd1 mux_top_track_22.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_2_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0480_ mem_top_track_30.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__clkbuf_1
X_1032_ mux_top_track_18.out vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__clkbuf_1
XFILLER_38_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1101_ mux_top_track_0.INVTX1_0_.out _0241_ vssd1 vssd1 vccd1 vccd1 mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_0747_ net29 vssd1 vssd1 vccd1 vccd1 mux_left_track_5.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0816_ _0175_ vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__inv_2
Xinput40 left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_1
Xinput51 top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_ vssd1 vssd1 vccd1
+ vccd1 net51 sky130_fd_sc_hd__clkbuf_1
X_0678_ mem_top_track_6.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0601_ mem_left_track_3.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__inv_2
XFILLER_7_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0463_ _0091_ vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__clkbuf_1
X_0532_ mem_left_track_17.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__inv_2
X_1015_ mux_left_track_15.out vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__clkbuf_1
XFILLER_19_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0515_ mem_left_track_37.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__inv_2
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0446_ mem_left_track_25.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__inv_2
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1043__100 vssd1 vssd1 vccd1 vccd1 net100 _1043__100/LO sky130_fd_sc_hd__conb_1
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1202__129 vssd1 vssd1 vccd1 vccd1 net129 _1202__129/LO sky130_fd_sc_hd__conb_1
XFILLER_5_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0429_ mem_left_track_31.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__inv_2
XFILLER_54_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0780_ net16 vssd1 vssd1 vccd1 vccd1 mux_top_track_28.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XFILLER_41_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput5 chanx_left_in[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
X_1194_ net127 _0334_ vssd1 vssd1 vccd1 vccd1 mux_top_track_30.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0763_ net23 vssd1 vssd1 vccd1 vccd1 mux_left_track_17.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0901_ clknet_3_4__leaf_prog_clk mem_top_track_10.DFFR_0_.D _0066_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_10.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_14_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0832_ _0177_ vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__inv_2
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0694_ mem_top_track_2.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__inv_2
XFILLER_64_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1177_ mux_top_track_0.INVTX1_1_.out _0317_ vssd1 vssd1 vccd1 vccd1 mux_top_track_20.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1100_ mux_top_track_18.INVTX1_2_.out _0240_ vssd1 vssd1 vccd1 vccd1 mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
X_1031_ mux_top_track_20.out vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__clkbuf_1
Xinput41 left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_1
X_0746_ mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_2_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_5.out sky130_fd_sc_hd__inv_2
Xinput30 chany_top_in[18] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
Xinput52 top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_ vssd1 vssd1 vccd1
+ vccd1 net52 sky130_fd_sc_hd__clkbuf_1
X_0815_ _0175_ vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__inv_2
X_0677_ mem_top_track_6.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__inv_2
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1229_ mux_left_track_31.INVTX1_0_.out _0369_ vssd1 vssd1 vccd1 vccd1 mux_left_track_31.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_25_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0531_ _0114_ vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__clkbuf_1
X_0600_ _0137_ vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__clkbuf_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0462_ mem_left_track_21.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1014_ mux_left_track_17.out vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__clkbuf_1
X_0729_ net6 vssd1 vssd1 vccd1 vccd1 mux_top_track_12.INVTX1_2_.out sky130_fd_sc_hd__inv_2
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0514_ net61 vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__inv_2
XFILLER_58_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0445_ _0085_ vssd1 vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__clkbuf_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0428_ mem_left_track_31.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__inv_2
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1073__105 vssd1 vssd1 vccd1 vccd1 net105 _1073__105/LO sky130_fd_sc_hd__conb_1
XFILLER_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput6 chanx_left_in[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
X_1193_ mux_top_track_10.INVTX1_0_.out _0333_ vssd1 vssd1 vccd1 vccd1 mux_top_track_28.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1190__126 vssd1 vssd1 vccd1 vccd1 net126 _1190__126/LO sky130_fd_sc_hd__conb_1
XFILLER_18_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0900_ clknet_3_1__leaf_prog_clk mem_top_track_10.DFFR_0_.Q _0065_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_10.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_2
XFILLER_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0693_ _0168_ vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__clkbuf_1
X_0762_ mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_2_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_17.out sky130_fd_sc_hd__inv_2
X_0831_ _0177_ vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__inv_2
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1176_ mux_top_track_20.mux_2level_tapbuf_basis_input2_mem1_0_out _0316_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_20.mux_2level_tapbuf_basis_input2_mem1_1_out sky130_fd_sc_hd__ebufn_2
XFILLER_32_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1030_ mux_top_track_22.out vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__clkbuf_1
Xinput20 chanx_left_in[9] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
Xinput31 chany_top_in[1] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
X_0814_ _0175_ vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__inv_2
Xinput53 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_1
X_0745_ net30 vssd1 vssd1 vccd1 vccd1 mux_left_track_3.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0676_ mem_top_track_6.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__inv_2
Xinput42 left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net42 sky130_fd_sc_hd__dlymetal6s2s_1
X_1228_ mux_left_track_31.mux_2level_tapbuf_basis_input2_mem1_0_out _0368_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_31.mux_2level_tapbuf_basis_input2_mem1_1_out sky130_fd_sc_hd__ebufn_2
XFILLER_52_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1159_ mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_0_out _0299_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_1
XFILLER_20_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0530_ mem_left_track_19.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__clkbuf_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0461_ mem_left_track_21.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__inv_2
XFILLER_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1013_ mux_left_track_19.out vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__clkbuf_1
XFILLER_8_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0728_ net58 vssd1 vssd1 vccd1 vccd1 mux_top_track_12.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_0659_ mem_top_track_10.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__inv_2
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1163__120 vssd1 vssd1 vccd1 vccd1 net120 _1163__120/LO sky130_fd_sc_hd__conb_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0513_ _0108_ vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__clkbuf_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0444_ mem_left_track_27.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__clkbuf_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0427_ _0079_ vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput7 chanx_left_in[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
X_1192_ mux_top_track_28.mux_2level_tapbuf_basis_input2_mem1_0_out _0332_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_28.mux_2level_tapbuf_basis_input2_mem1_1_out sky130_fd_sc_hd__ebufn_2
XFILLER_51_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0830_ _0177_ vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__inv_2
X_0692_ mem_top_track_4.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__clkbuf_1
X_0761_ net46 vssd1 vssd1 vccd1 vccd1 mux_left_track_15.INVTX1_2_.out sky130_fd_sc_hd__inv_2
XFILLER_49_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1175_ mux_top_track_20.INVTX1_1_.out _0315_ vssd1 vssd1 vccd1 vccd1 mux_top_track_20.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_32_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0959_ clknet_3_3__leaf_prog_clk mem_left_track_27.DFFR_1_.Q _0048_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_29.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_15_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput10 chanx_left_in[17] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
Xinput21 chany_top_in[0] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
Xinput32 chany_top_in[2] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
Xinput43 left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net43 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput54 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0813_ _0175_ vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__inv_2
X_0675_ _0162_ vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__clkbuf_1
X_0744_ mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_2_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_3.out sky130_fd_sc_hd__inv_2
XFILLER_37_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1227_ mux_left_track_11.INVTX1_2_.out _0367_ vssd1 vssd1 vccd1 vccd1 mux_left_track_31.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1158_ mux_left_track_15.INVTX1_2_.out _0298_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_52_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1089_ mux_top_track_12.INVTX1_1_.out _0229_ vssd1 vssd1 vccd1 vccd1 mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_57_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0460_ mem_left_track_21.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__inv_2
X_1012_ mux_left_track_21.out vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__clkbuf_1
X_0727_ mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_2_out vssd1 vssd1 vccd1
+ vccd1 mux_top_track_12.out sky130_fd_sc_hd__inv_2
X_0589_ _0133_ vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__clkbuf_1
X_0658_ mem_top_track_10.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__inv_2
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0443_ _0084_ vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0512_ mem_top_track_20.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__clkbuf_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0426_ mem_left_track_33.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1191_ mux_top_track_28.INVTX1_1_.out _0331_ vssd1 vssd1 vccd1 vccd1 mux_top_track_28.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
Xinput8 chanx_left_in[15] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0760_ net24 vssd1 vssd1 vccd1 vccd1 mux_left_track_15.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0691_ mem_top_track_4.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__inv_2
XFILLER_56_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1174_ net122 _0314_ vssd1 vssd1 vccd1 vccd1 mux_top_track_20.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0958_ clknet_3_4__leaf_prog_clk mem_left_track_29.DFFR_0_.Q _0047_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_29.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
X_0889_ _0174_ vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__inv_2
XFILLER_28_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1127__114 vssd1 vssd1 vccd1 vccd1 net114 _1127__114/LO sky130_fd_sc_hd__conb_1
Xinput44 left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_1
Xinput55 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
X_0743_ net49 vssd1 vssd1 vccd1 vccd1 mux_left_track_1.INVTX1_2_.out sky130_fd_sc_hd__inv_2
Xinput22 chany_top_in[10] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
X_0812_ _0175_ vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__inv_2
Xinput33 chany_top_in[3] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
Xinput11 chanx_left_in[18] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
X_0674_ mem_top_track_8.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__clkbuf_1
X_1226_ net135 _0366_ vssd1 vssd1 vccd1 vccd1 mux_left_track_31.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_37_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1157_ net119 _0297_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1088_ mux_top_track_14.INVTX1_2_.out _0228_ vssd1 vssd1 vccd1 vccd1 mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_20_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1011_ mux_left_track_23.out vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__clkbuf_1
XFILLER_8_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0726_ net7 vssd1 vssd1 vccd1 vccd1 mux_top_track_10.INVTX1_2_.out sky130_fd_sc_hd__inv_2
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0657_ _0156_ vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__clkbuf_1
X_0588_ mem_left_track_5.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1209_ mux_left_track_21.INVTX1_0_.out _0349_ vssd1 vssd1 vccd1 vccd1 mux_left_track_21.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0511_ _0107_ vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0442_ mem_left_track_27.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__clkbuf_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0709_ _0173_ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0425_ _0078_ vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1190_ net126 _0330_ vssd1 vssd1 vccd1 vccd1 mux_top_track_28.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_36_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput9 chanx_left_in[16] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0690_ _0167_ vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__clkbuf_1
XFILLER_25_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1173_ mux_left_track_37.INVTX1_0_.out _0313_ vssd1 vssd1 vccd1 vccd1 mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0888_ _0174_ vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__inv_2
X_0957_ clknet_3_4__leaf_prog_clk mem_left_track_25.DFFR_1_.Q _0046_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_27.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput56 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net56 sky130_fd_sc_hd__clkbuf_1
Xinput45 left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_1
Xinput34 chany_top_in[4] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_1
Xinput12 chanx_left_in[1] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0742_ net21 vssd1 vssd1 vccd1 vccd1 mux_left_track_1.INVTX1_0_.out sky130_fd_sc_hd__inv_2
Xinput23 chany_top_in[11] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
X_0811_ _0175_ vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__inv_2
X_0673_ mem_top_track_8.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__inv_2
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1214__132 vssd1 vssd1 vccd1 vccd1 net132 _1214__132/LO sky130_fd_sc_hd__conb_1
XFILLER_52_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1225_ mux_left_track_29.INVTX1_0_.out _0365_ vssd1 vssd1 vccd1 vccd1 mux_left_track_29.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_25_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1087_ mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_0_out _0227_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_1
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1156_ mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_1_out _0296_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_1
XFILLER_20_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1157__119 vssd1 vssd1 vccd1 vccd1 net119 _1157__119/LO sky130_fd_sc_hd__conb_1
XFILLER_21_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1010_ mux_left_track_25.out vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_1
XFILLER_19_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0725_ net56 vssd1 vssd1 vccd1 vccd1 mux_top_track_10.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0656_ mem_top_track_12.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0587_ mem_left_track_5.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__inv_2
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1208_ mux_left_track_21.mux_2level_tapbuf_basis_input2_mem1_0_out _0348_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_21.mux_2level_tapbuf_basis_input2_mem1_1_out sky130_fd_sc_hd__ebufn_2
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1139_ net116 _0279_ vssd1 vssd1 vccd1 vccd1 mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0510_ mem_top_track_20.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0441_ mem_left_track_27.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__inv_2
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0708_ mem_top_track_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__clkbuf_1
X_0639_ _0150_ vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0424_ mem_left_track_33.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1172_ mux_left_track_17.INVTX1_2_.out _0312_ vssd1 vssd1 vccd1 vccd1 mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_2_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0956_ clknet_3_5__leaf_prog_clk mem_left_track_27.DFFR_0_.Q _0045_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_27.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
X_0887_ _0174_ vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__inv_2
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0810_ _0175_ vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__inv_2
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput13 chanx_left_in[2] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
Xinput24 chany_top_in[12] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
Xinput57 top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_1
Xinput35 chany_top_in[5] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_1
Xinput46 left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_1
X_0741_ net48 vssd1 vssd1 vccd1 vccd1 mux_left_track_1.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_0672_ _0161_ vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1224_ mux_left_track_29.mux_2level_tapbuf_basis_input2_mem1_0_out _0364_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_29.mux_2level_tapbuf_basis_input2_mem1_1_out sky130_fd_sc_hd__ebufn_2
X_1155_ mux_left_track_15.INVTX1_0_.out _0295_ vssd1 vssd1 vccd1 vccd1 mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_37_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1086_ mux_top_track_14.INVTX1_1_.out _0226_ vssd1 vssd1 vccd1 vccd1 mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0939_ clknet_3_7__leaf_prog_clk mem_top_track_22.DFFR_1_.Q _0028_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_24.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0724_ net57 vssd1 vssd1 vccd1 vccd1 mux_top_track_10.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_0586_ mem_left_track_5.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__inv_2
X_0655_ mem_top_track_12.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__inv_2
XFILLER_57_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1207_ mux_left_track_1.INVTX1_2_.out _0347_ vssd1 vssd1 vccd1 vccd1 mux_left_track_21.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1069_ mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_0_out _0209_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
XFILLER_25_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1138_ mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_1_out _0278_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
XFILLER_31_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0440_ mem_left_track_27.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__inv_2
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0707_ _0172_ vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0569_ mem_left_track_9.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__inv_2
X_0638_ mem_top_track_16.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0423_ mem_left_track_33.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__inv_2
XFILLER_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1049__101 vssd1 vssd1 vccd1 vccd1 net101 _1049__101/LO sky130_fd_sc_hd__conb_1
XFILLER_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1171_ mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_0_out _0311_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
XFILLER_64_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0886_ _0174_ vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__inv_2
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0955_ clknet_3_6__leaf_prog_clk mem_left_track_23.DFFR_1_.Q _0044_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_25.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_55_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput25 chany_top_in[13] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
X_0740_ mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_2_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_1.out sky130_fd_sc_hd__inv_2
Xinput14 chanx_left_in[3] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
Xinput36 chany_top_in[6] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput58 top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_1
Xinput47 left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_1
X_0671_ mem_top_track_10.DFFR_0_.D vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__clkbuf_1
X_1154_ mux_left_track_15.INVTX1_2_.out _0294_ vssd1 vssd1 vccd1 vccd1 mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1223_ mux_left_track_11.INVTX1_1_.out _0363_ vssd1 vssd1 vccd1 vccd1 mux_left_track_29.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_37_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1085_ net107 _0225_ vssd1 vssd1 vccd1 vccd1 mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_20_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0869_ _0180_ vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__inv_2
X_0938_ clknet_3_7__leaf_prog_clk mem_top_track_24.DFFR_0_.Q _0027_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_24.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_43_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0723_ mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_2_out vssd1 vssd1 vccd1
+ vccd1 mux_top_track_10.out sky130_fd_sc_hd__inv_2
X_0585_ _0132_ vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__clkbuf_1
X_0654_ _0155_ vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1137_ mux_left_track_9.INVTX1_0_.out _0277_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1206_ net130 _0346_ vssd1 vssd1 vccd1 vccd1 mux_left_track_21.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1068_ mux_top_track_10.INVTX1_0_.out _0208_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0706_ mem_top_track_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0637_ mem_top_track_16.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__inv_2
X_0499_ _0103_ vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__clkbuf_1
X_0568_ mem_left_track_11.DFFR_0_.D vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__inv_2
XFILLER_13_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1186__125 vssd1 vssd1 vccd1 vccd1 net125 _1186__125/LO sky130_fd_sc_hd__conb_1
XFILLER_5_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1234__137 vssd1 vssd1 vccd1 vccd1 net137 _1234__137/LO sky130_fd_sc_hd__conb_1
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0422_ mem_left_track_33.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__inv_2
XFILLER_5_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1170_ mux_left_track_1.INVTX1_1_.out _0310_ vssd1 vssd1 vccd1 vccd1 mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_1_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0885_ _0174_ vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__inv_2
X_0954_ clknet_3_5__leaf_prog_clk mem_left_track_25.DFFR_0_.Q _0043_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_25.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1079__106 vssd1 vssd1 vccd1 vccd1 net106 _1079__106/LO sky130_fd_sc_hd__conb_1
XFILLER_11_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput37 chany_top_in[7] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_1
Xinput15 chanx_left_in[4] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
X_0670_ _0160_ vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__clkbuf_1
Xinput48 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_ vssd1 vssd1 vccd1
+ vccd1 net48 sky130_fd_sc_hd__clkbuf_1
Xinput26 chany_top_in[14] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
Xinput59 top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_1
X_1153_ mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_0_out _0293_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
X_1222_ net134 _0362_ vssd1 vssd1 vccd1 vccd1 mux_left_track_29.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1084_ mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_1_out _0224_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_1
XFILLER_20_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0799_ net35 vssd1 vssd1 vccd1 vccd1 mux_left_track_29.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0868_ _0180_ vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__inv_2
XFILLER_9_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0937_ clknet_3_7__leaf_prog_clk mem_top_track_20.DFFR_1_.Q _0026_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_22.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_43_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0653_ mem_top_track_12.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_7__f_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_3_7__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
X_0722_ net8 vssd1 vssd1 vccd1 vccd1 mux_top_track_8.INVTX1_2_.out sky130_fd_sc_hd__inv_2
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0584_ mem_left_track_7.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1067_ net104 _0207_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
X_1205_ mux_top_track_14.INVTX1_1_.out _0345_ vssd1 vssd1 vccd1 vccd1 mux_top_track_34.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1136_ mux_left_track_11.INVTX1_1_.out _0276_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_40_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0636_ _0149_ vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__clkbuf_1
X_0705_ mem_top_track_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__inv_2
XFILLER_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0567_ _0126_ vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__clkbuf_1
X_0498_ mem_top_track_24.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__clkbuf_1
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1119_ mux_left_track_3.INVTX1_0_.out _0259_ vssd1 vssd1 vccd1 vccd1 mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_44_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0421_ _0077_ vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0619_ mem_top_track_36.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__inv_2
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1169__121 vssd1 vssd1 vccd1 vccd1 net121 _1169__121/LO sky130_fd_sc_hd__conb_1
XFILLER_50_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0884_ _0174_ vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__inv_2
XFILLER_9_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0953_ clknet_3_2__leaf_prog_clk mem_left_track_21.DFFR_1_.Q _0042_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_23.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput49 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_ vssd1 vssd1 vccd1
+ vccd1 net49 sky130_fd_sc_hd__clkbuf_1
Xinput27 chany_top_in[15] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
Xinput16 chanx_left_in[5] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_6__f_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_3_6__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xinput38 chany_top_in[8] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_1
X_1221_ mux_left_track_27.INVTX1_0_.out _0361_ vssd1 vssd1 vccd1 vccd1 mux_left_track_27.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1152_ mux_left_track_13.INVTX1_2_.out _0292_ vssd1 vssd1 vccd1 vccd1 mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1083_ mux_top_track_10.INVTX1_1_.out _0223_ vssd1 vssd1 vccd1 vccd1 mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_0936_ clknet_3_5__leaf_prog_clk mem_top_track_22.DFFR_0_.Q _0025_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_22.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
X_0798_ mux_left_track_29.mux_2level_tapbuf_basis_input2_mem1_1_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_29.out sky130_fd_sc_hd__inv_2
X_0867_ _0180_ vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__inv_2
XFILLER_51_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0652_ _0154_ vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__clkbuf_1
X_0721_ mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_2_out vssd1 vssd1 vccd1
+ vccd1 mux_top_track_8.out sky130_fd_sc_hd__inv_2
X_0583_ mem_left_track_7.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__inv_2
XFILLER_10_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1204_ mux_top_track_34.mux_2level_tapbuf_basis_input2_mem1_0_out _0344_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_34.mux_2level_tapbuf_basis_input2_mem1_1_out sky130_fd_sc_hd__ebufn_2
X_1066_ mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_1_out _0206_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
X_1135_ mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_0_out _0275_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_1
X_0919_ clknet_3_1__leaf_prog_clk mem_left_track_5.DFFR_1_.Q _0008_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_7.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0566_ mem_left_track_11.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__clkbuf_1
X_0635_ mem_top_track_16.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__clkbuf_1
X_0704_ mem_top_track_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__inv_2
X_0497_ mem_top_track_24.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__inv_2
X_1118_ mux_left_track_23.INVTX1_1_.out _0258_ vssd1 vssd1 vccd1 vccd1 mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_21_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1049_ net101 _0189_ vssd1 vssd1 vccd1 vccd1 mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0420_ mem_left_track_35.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0549_ _0120_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__clkbuf_1
X_0618_ _0143_ vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__clkbuf_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_5__f_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_3_5__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0952_ clknet_3_2__leaf_prog_clk mem_left_track_23.DFFR_0_.Q _0041_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_23.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0883_ _0181_ vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__inv_2
XFILLER_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput28 chany_top_in[16] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
Xinput17 chanx_left_in[6] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput39 chany_top_in[9] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
XFILLER_42_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1151_ net118 _0291_ vssd1 vssd1 vccd1 vccd1 mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
X_1220_ mux_left_track_27.mux_2level_tapbuf_basis_input2_mem1_0_out _0360_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_27.mux_2level_tapbuf_basis_input2_mem1_1_out sky130_fd_sc_hd__ebufn_2
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1082_ mux_top_track_12.INVTX1_2_.out _0222_ vssd1 vssd1 vccd1 vccd1 mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0866_ _0180_ vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__inv_2
X_0935_ clknet_3_1__leaf_prog_clk mem_top_track_18.DFFR_1_.Q _0024_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_20.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0797_ net42 vssd1 vssd1 vccd1 vccd1 mux_left_track_27.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XFILLER_28_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0720_ net9 vssd1 vssd1 vccd1 vccd1 mux_top_track_6.INVTX1_2_.out sky130_fd_sc_hd__inv_2
X_0582_ _0131_ vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__clkbuf_1
X_0651_ mem_top_track_12.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1134_ mux_left_track_27.INVTX1_1_.out _0274_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1203_ mux_top_track_34.INVTX1_1_.out _0343_ vssd1 vssd1 vccd1 vccd1 mux_top_track_34.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1065_ mux_top_track_24.INVTX1_0_.out _0205_ vssd1 vssd1 vccd1 vccd1 mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_18_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0849_ _0178_ vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__inv_2
X_0918_ clknet_3_5__leaf_prog_clk mem_left_track_7.DFFR_0_.Q _0007_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_7.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0703_ mem_top_track_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__inv_2
X_0565_ mem_left_track_11.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__inv_2
X_0496_ mem_top_track_24.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__inv_2
X_0634_ _0148_ vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1117_ mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_0_out _0257_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_1
XFILLER_21_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1048_ mux_top_track_2.INVTX1_1_.out _0188_ vssd1 vssd1 vccd1 vccd1 mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0548_ mem_left_track_15.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__clkbuf_1
X_0617_ mem_left_track_1.DFFR_0_.D vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__clkbuf_1
X_0479_ mem_top_track_30.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__inv_2
XFILLER_41_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_4__f_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_3_4__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0882_ _0181_ vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__inv_2
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0951_ clknet_3_2__leaf_prog_clk mem_left_track_19.DFFR_1_.Q _0040_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_21.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput18 chanx_left_in[7] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput29 chany_top_in[17] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
X_1103__110 vssd1 vssd1 vccd1 vccd1 net110 _1103__110/LO sky130_fd_sc_hd__conb_1
XFILLER_6_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1150_ mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_1_out _0290_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
X_1081_ mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_0_out _0221_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
X_0865_ _0180_ vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__inv_2
X_0934_ clknet_3_3__leaf_prog_clk mem_top_track_20.DFFR_0_.Q _0023_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_20.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0796_ net36 vssd1 vssd1 vccd1 vccd1 mux_left_track_27.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_28_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0581_ mem_left_track_7.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__clkbuf_1
X_0650_ mem_top_track_12.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__inv_2
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1202_ net129 _0342_ vssd1 vssd1 vccd1 vccd1 mux_top_track_34.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1064_ mux_top_track_6.INVTX1_2_.out _0204_ vssd1 vssd1 vccd1 vccd1 mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
X_1133_ net115 _0273_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_33_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0779_ mux_top_track_28.mux_2level_tapbuf_basis_input2_mem1_1_out vssd1 vssd1 vccd1
+ vccd1 mux_top_track_28.out sky130_fd_sc_hd__inv_2
X_0917_ clknet_3_0__leaf_prog_clk mem_left_track_3.DFFR_1_.Q _0006_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_5.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
X_0848_ _0178_ vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__inv_2
XFILLER_56_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0633_ mem_top_track_16.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__clkbuf_1
X_0702_ _0171_ vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__clkbuf_1
X_0564_ _0125_ vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__clkbuf_1
X_0495_ _0102_ vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1047_ mux_top_track_0.INVTX1_2_.out _0187_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
X_1116_ mux_left_track_1.INVTX1_2_.out _0256_ vssd1 vssd1 vccd1 vccd1 mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_3__f_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_3_3__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_56_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0616_ _0142_ vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0547_ mem_left_track_15.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__inv_2
X_0478_ mem_top_track_30.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__inv_2
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0881_ _0181_ vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__inv_2
XFILLER_13_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0950_ clknet_3_2__leaf_prog_clk mem_left_track_21.DFFR_0_.Q _0039_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_21.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput19 chanx_left_in[8] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1080_ mux_top_track_12.INVTX1_1_.out _0220_ vssd1 vssd1 vccd1 vccd1 mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0795_ mux_left_track_27.mux_2level_tapbuf_basis_input2_mem1_1_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_27.out sky130_fd_sc_hd__inv_2
X_0864_ _0180_ vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__inv_2
X_0933_ clknet_3_7__leaf_prog_clk mem_left_track_35.DFFR_1_.Q _0022_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_37.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_13_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1133__115 vssd1 vssd1 vccd1 vccd1 net115 _1133__115/LO sky130_fd_sc_hd__conb_1
XFILLER_63_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0580_ _0130_ vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__clkbuf_1
X_1201_ mux_top_track_12.INVTX1_1_.out _0341_ vssd1 vssd1 vccd1 vccd1 mux_top_track_32.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_6_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1063_ mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_0_out _0203_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
X_1132_ mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_1_out _0272_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_1
XFILLER_18_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0916_ clknet_3_1__leaf_prog_clk mem_left_track_5.DFFR_0_.Q _0005_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_5.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_2
Xclkbuf_3_2__f_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_3_2__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
X_0778_ net17 vssd1 vssd1 vccd1 vccd1 mux_top_track_26.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_0847_ _0178_ vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__inv_2
XFILLER_56_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0563_ mem_left_track_11.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__clkbuf_1
X_0701_ mem_top_track_2.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__clkbuf_1
X_0632_ mem_top_track_16.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__inv_2
XFILLER_38_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0494_ mem_top_track_26.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1115_ net112 _0255_ vssd1 vssd1 vccd1 vccd1 mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1046_ mux_top_track_0.INVTX1_0_.out _0186_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1210__131 vssd1 vssd1 vccd1 vccd1 net131 _1210__131/LO sky130_fd_sc_hd__conb_1
XFILLER_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0546_ _0119_ vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__clkbuf_1
X_0615_ mem_top_track_36.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0477_ _0096_ vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1029_ mux_top_track_24.out vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__clkbuf_1
XFILLER_30_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0529_ mem_left_track_19.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__inv_2
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0880_ _0181_ vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__inv_2
XFILLER_13_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_1__f_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_3_1__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
X_0932_ clknet_3_6__leaf_prog_clk mem_left_track_37.DFFR_0_.Q _0021_ vssd1 vssd1 vccd1
+ vccd1 net61 sky130_fd_sc_hd__dfrtp_4
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0794_ net41 vssd1 vssd1 vccd1 vccd1 mux_left_track_25.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_0863_ _0180_ vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__inv_2
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1200_ mux_top_track_32.mux_2level_tapbuf_basis_input2_mem1_0_out _0340_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_32.mux_2level_tapbuf_basis_input2_mem1_1_out sky130_fd_sc_hd__ebufn_2
XFILLER_2_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1131_ mux_left_track_7.INVTX1_0_.out _0271_ vssd1 vssd1 vccd1 vccd1 mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1062_ mux_top_track_26.INVTX1_0_.out _0202_ vssd1 vssd1 vccd1 vccd1 mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0915_ clknet_3_0__leaf_prog_clk mem_left_track_1.DFFR_1_.Q _0004_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_3.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
X_0777_ net55 vssd1 vssd1 vccd1 vccd1 mux_top_track_26.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0846_ _0178_ vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__inv_2
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0700_ _0170_ vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__clkbuf_1
X_0562_ _0124_ vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__clkbuf_1
X_0631_ mem_top_track_16.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__inv_2
XFILLER_53_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0493_ _0101_ vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__clkbuf_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1114_ mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_1_out _0254_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_1
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1045_ mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_0_out _0185_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_1
X_0829_ _0174_ vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__buf_4
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0545_ mem_left_track_15.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__clkbuf_1
X_0476_ mem_top_track_32.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__clkbuf_1
X_0614_ mem_top_track_36.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__inv_2
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1028_ mux_top_track_26.out vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0528_ _0113_ vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__clkbuf_1
X_0459_ _0090_ vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_0__f_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_3_0__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 chany_top_out[18] sky130_fd_sc_hd__buf_2
XFILLER_55_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0862_ net50 vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__buf_4
X_0931_ clknet_3_7__leaf_prog_clk mem_left_track_17.DFFR_1_.Q _0020_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_19.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0793_ net37 vssd1 vssd1 vccd1 vccd1 mux_left_track_25.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1130_ mux_left_track_27.INVTX1_1_.out _0270_ vssd1 vssd1 vccd1 vccd1 mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_2_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1061_ net103 _0201_ vssd1 vssd1 vccd1 vccd1 mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_18_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0845_ _0178_ vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__inv_2
X_0914_ clknet_3_2__leaf_prog_clk mem_left_track_3.DFFR_0_.Q _0003_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_3.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
X_0776_ mux_top_track_26.mux_2level_tapbuf_basis_input2_mem1_1_out vssd1 vssd1 vccd1
+ vccd1 mux_top_track_26.out sky130_fd_sc_hd__inv_2
XFILLER_56_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0630_ _0147_ vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__clkbuf_1
X_0492_ mem_top_track_26.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__clkbuf_1
X_0561_ mem_left_track_11.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1113_ mux_left_track_1.INVTX1_0_.out _0253_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1044_ mux_top_track_0.INVTX1_1_.out _0184_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0759_ mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_2_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_15.out sky130_fd_sc_hd__inv_2
X_0828_ _0176_ vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__inv_2
XFILLER_28_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0613_ mem_left_track_1.DFFR_0_.D vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__inv_2
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0544_ _0118_ vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__clkbuf_1
X_0475_ _0095_ vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1027_ mux_top_track_28.out vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__clkbuf_1
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0527_ mem_left_track_19.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__clkbuf_1
X_0458_ mem_left_track_23.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__clkbuf_1
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1182__124 vssd1 vssd1 vccd1 vccd1 net124 _1182__124/LO sky130_fd_sc_hd__conb_1
XFILLER_63_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 chany_top_out[1] sky130_fd_sc_hd__buf_2
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 chanx_left_out[9] sky130_fd_sc_hd__buf_2
X_1230__136 vssd1 vssd1 vccd1 vccd1 net136 _1230__136/LO sky130_fd_sc_hd__conb_1
XFILLER_31_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1055__102 vssd1 vssd1 vccd1 vccd1 net102 _1055__102/LO sky130_fd_sc_hd__conb_1
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0792_ mux_left_track_25.mux_2level_tapbuf_basis_input2_mem1_1_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_25.out sky130_fd_sc_hd__inv_2
X_0861_ _0179_ vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__inv_2
XFILLER_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0930_ clknet_3_7__leaf_prog_clk mem_left_track_19.DFFR_0_.Q _0019_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_19.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1060_ mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_1_out _0200_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
XFILLER_18_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0775_ net18 vssd1 vssd1 vccd1 vccd1 mux_top_track_24.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_0844_ _0178_ vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__inv_2
X_0913_ clknet_3_1__leaf_prog_clk mem_left_track_1.DFFR_0_.D _0002_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_1.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_64_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1189_ mux_top_track_26.INVTX1_0_.out _0329_ vssd1 vssd1 vccd1 vccd1 mux_top_track_26.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0491_ mem_top_track_26.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__inv_2
X_0560_ mem_left_track_11.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__inv_2
XFILLER_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1112_ mux_left_track_1.INVTX1_2_.out _0252_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
X_1043_ net100 _0183_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0758_ net45 vssd1 vssd1 vccd1 vccd1 mux_left_track_13.INVTX1_2_.out sky130_fd_sc_hd__inv_2
X_0827_ _0176_ vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__inv_2
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0689_ mem_top_track_4.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0612_ _0141_ vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0543_ mem_left_track_15.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__clkbuf_1
X_0474_ mem_top_track_32.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1026_ mux_top_track_30.out vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__clkbuf_1
XFILLER_61_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0526_ _0112_ vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__clkbuf_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0457_ _0089_ vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__clkbuf_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1009_ mux_left_track_27.out vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_1
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 chanx_left_out[17] sky130_fd_sc_hd__buf_2
XFILLER_31_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 chany_top_out[2] sky130_fd_sc_hd__buf_2
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 chany_top_out[0] sky130_fd_sc_hd__buf_2
XFILLER_51_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0509_ mem_top_track_20.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__inv_2
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0860_ _0179_ vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__inv_2
XFILLER_9_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0791_ net40 vssd1 vssd1 vccd1 vccd1 mux_left_track_23.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XFILLER_3_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1085__107 vssd1 vssd1 vccd1 vccd1 net107 _1085__107/LO sky130_fd_sc_hd__conb_1
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0912_ clknet_3_0__leaf_prog_clk mem_left_track_1.DFFR_0_.Q _0001_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_1.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_2
X_0774_ net54 vssd1 vssd1 vccd1 vccd1 mux_top_track_24.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_5_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0843_ _0178_ vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__inv_2
XFILLER_56_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1188_ mux_top_track_26.mux_2level_tapbuf_basis_input2_mem1_0_out _0328_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_26.mux_2level_tapbuf_basis_input2_mem1_1_out sky130_fd_sc_hd__ebufn_2
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0490_ mem_top_track_26.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__inv_2
X_1111_ mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_0_out _0251_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
X_1042_ mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_1_out _0182_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_1
XFILLER_61_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0757_ net25 vssd1 vssd1 vccd1 vccd1 mux_left_track_13.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0688_ _0166_ vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__clkbuf_1
X_0826_ _0176_ vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__inv_2
XFILLER_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0542_ mem_left_track_15.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__inv_2
X_0611_ mem_left_track_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0473_ mem_top_track_32.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__inv_2
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1025_ mux_top_track_32.out vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__clkbuf_1
XFILLER_53_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0809_ _0175_ vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__inv_2
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_1 _0034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0525_ mem_left_track_19.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__clkbuf_1
X_0456_ mem_top_track_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__clkbuf_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1008_ mux_left_track_29.out vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__clkbuf_1
XFILLER_22_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 chany_top_out[3] sky130_fd_sc_hd__buf_2
XFILLER_49_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 chany_top_out[10] sky130_fd_sc_hd__buf_2
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 chanx_left_out[18] sky130_fd_sc_hd__buf_2
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0439_ _0083_ vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__clkbuf_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0508_ mem_top_track_20.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__inv_2
XFILLER_54_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0790_ net38 vssd1 vssd1 vccd1 vccd1 mux_left_track_23.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0842_ _0178_ vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__inv_2
X_0911_ clknet_3_6__leaf_prog_clk mem_top_track_34.DFFR_1_.Q _0000_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_36.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0773_ mux_top_track_24.mux_2level_tapbuf_basis_input2_mem1_1_out vssd1 vssd1 vccd1
+ vccd1 mux_top_track_24.out sky130_fd_sc_hd__inv_2
XFILLER_56_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1187_ mux_top_track_26.INVTX1_1_.out _0327_ vssd1 vssd1 vccd1 vccd1 mux_top_track_26.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1109__111 vssd1 vssd1 vccd1 vccd1 net111 _1109__111/LO sky130_fd_sc_hd__conb_1
XFILLER_31_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1110_ mux_left_track_1.INVTX1_1_.out _0250_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_64_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1041_ mux_top_track_0.out vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__clkbuf_1
X_0825_ _0176_ vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__inv_2
X_0756_ mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_2_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_13.out sky130_fd_sc_hd__inv_2
X_0687_ mem_top_track_4.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0541_ mem_left_track_15.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__inv_2
X_0472_ mem_top_track_32.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__inv_2
X_0610_ mem_left_track_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__inv_2
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1024_ mux_top_track_34.out vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__clkbuf_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0808_ _0175_ vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__inv_2
X_0739_ net12 vssd1 vssd1 vccd1 vccd1 mux_top_track_36.INVTX1_2_.out sky130_fd_sc_hd__inv_2
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_2 _0040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0524_ mem_left_track_19.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__inv_2
X_0455_ _0088_ vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__clkbuf_1
X_1007_ mux_left_track_31.out vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__clkbuf_1
XFILLER_26_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 ccff_tail sky130_fd_sc_hd__buf_2
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 chany_top_out[4] sky130_fd_sc_hd__buf_2
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 chany_top_out[11] sky130_fd_sc_hd__buf_2
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 chanx_left_out[1] sky130_fd_sc_hd__buf_2
XFILLER_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0507_ _0106_ vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__clkbuf_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0438_ mem_left_track_29.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_54_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1206__130 vssd1 vssd1 vccd1 vccd1 net130 _1206__130/LO sky130_fd_sc_hd__conb_1
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0772_ net19 vssd1 vssd1 vccd1 vccd1 mux_top_track_22.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_0841_ _0178_ vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__inv_2
X_0910_ clknet_3_1__leaf_prog_clk mem_top_track_36.DFFR_0_.Q _0075_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_1.DFFR_0_.D sky130_fd_sc_hd__dfrtp_1
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1186_ net125 _0326_ vssd1 vssd1 vccd1 vccd1 mux_top_track_26.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1040_ mux_top_track_2.out vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0755_ net44 vssd1 vssd1 vccd1 vccd1 mux_left_track_11.INVTX1_2_.out sky130_fd_sc_hd__inv_2
X_0824_ _0176_ vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__inv_2
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0686_ mem_top_track_4.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__inv_2
XFILLER_52_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1169_ net121 _0309_ vssd1 vssd1 vccd1 vccd1 mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1139__116 vssd1 vssd1 vccd1 vccd1 net116 _1139__116/LO sky130_fd_sc_hd__conb_1
XFILLER_34_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0540_ _0117_ vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__clkbuf_1
X_0471_ _0094_ vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__clkbuf_1
X_1023_ mux_top_track_36.out vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__clkbuf_1
XFILLER_34_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0738_ mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_2_out vssd1 vssd1 vccd1
+ vccd1 mux_top_track_36.out sky130_fd_sc_hd__inv_2
X_0807_ _0174_ vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__buf_4
X_0669_ mem_top_track_8.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_3 mux_left_track_37.out vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0523_ mem_left_track_19.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__inv_2
X_0454_ mem_left_track_23.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__clkbuf_1
X_1006_ mux_left_track_33.out vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 chanx_left_out[2] sky130_fd_sc_hd__buf_2
XFILLER_48_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 chanx_left_out[0] sky130_fd_sc_hd__buf_2
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 chany_top_out[5] sky130_fd_sc_hd__buf_2
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 chany_top_out[12] sky130_fd_sc_hd__buf_2
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0506_ mem_top_track_22.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0437_ _0082_ vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0771_ mux_top_track_22.mux_2level_tapbuf_basis_input2_mem1_1_out vssd1 vssd1 vccd1
+ vccd1 mux_top_track_22.out sky130_fd_sc_hd__inv_2
X_0840_ _0174_ vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__buf_4
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1185_ mux_top_track_24.INVTX1_0_.out _0325_ vssd1 vssd1 vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0685_ mem_top_track_4.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__inv_2
X_0754_ net26 vssd1 vssd1 vccd1 vccd1 mux_left_track_11.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0823_ _0176_ vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__inv_2
XFILLER_52_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1099_ mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_0_out _0239_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
X_1237_ mux_left_track_35.INVTX1_0_.out _0377_ vssd1 vssd1 vccd1 vccd1 mux_left_track_35.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1168_ mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_1_out _0308_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_2_out sky130_fd_sc_hd__ebufn_2
XFILLER_47_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0470_ mem_top_track_34.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__clkbuf_1
X_1022_ mux_left_track_1.out vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_1
XFILLER_38_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0737_ net3 vssd1 vssd1 vccd1 vccd1 mux_top_track_18.INVTX1_2_.out sky130_fd_sc_hd__inv_2
X_0668_ mem_top_track_8.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__inv_2
X_0806_ net50 vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__clkbuf_4
X_0599_ mem_left_track_3.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0522_ _0111_ vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__clkbuf_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_4 mux_top_track_10.out vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0453_ mem_left_track_23.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__inv_2
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1005_ mux_left_track_35.out vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__clkbuf_1
XFILLER_34_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 chanx_left_out[3] sky130_fd_sc_hd__buf_2
XFILLER_48_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 chanx_left_out[10] sky130_fd_sc_hd__buf_2
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 chany_top_out[6] sky130_fd_sc_hd__buf_2
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 chany_top_out[13] sky130_fd_sc_hd__buf_2
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0505_ _0105_ vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__clkbuf_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0436_ mem_left_track_29.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__clkbuf_1
.ends

