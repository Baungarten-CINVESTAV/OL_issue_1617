* NGSPICE file created from sb_1__1_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_4 abstract view
.subckt sky130_fd_sc_hd__ebufn_4 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

.subckt sb_1__1_ bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_ bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
+ bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_ bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
+ ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11] chanx_left_in[12]
+ chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16] chanx_left_in[17]
+ chanx_left_in[18] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4]
+ chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_in[9]
+ chanx_left_out[0] chanx_left_out[10] chanx_left_out[11] chanx_left_out[12] chanx_left_out[13]
+ chanx_left_out[14] chanx_left_out[15] chanx_left_out[16] chanx_left_out[17] chanx_left_out[18]
+ chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chanx_right_in[0]
+ chanx_right_in[10] chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14]
+ chanx_right_in[15] chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10]
+ chanx_right_out[11] chanx_right_out[12] chanx_right_out[13] chanx_right_out[14]
+ chanx_right_out[15] chanx_right_out[16] chanx_right_out[17] chanx_right_out[18]
+ chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4] chanx_right_out[5]
+ chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chanx_right_out[9] chany_bottom_in[0]
+ chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13]
+ chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17]
+ chany_bottom_in[18] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4]
+ chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_in[9]
+ chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11] chany_bottom_out[12]
+ chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15] chany_bottom_out[16]
+ chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[1] chany_bottom_out[2]
+ chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6]
+ chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9] chany_top_in[0] chany_top_in[10]
+ chany_top_in[11] chany_top_in[12] chany_top_in[13] chany_top_in[14] chany_top_in[15]
+ chany_top_in[16] chany_top_in[17] chany_top_in[18] chany_top_in[1] chany_top_in[2]
+ chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7]
+ chany_top_in[8] chany_top_in[9] chany_top_out[0] chany_top_out[10] chany_top_out[11]
+ chany_top_out[12] chany_top_out[13] chany_top_out[14] chany_top_out[15] chany_top_out[16]
+ chany_top_out[17] chany_top_out[18] chany_top_out[1] chany_top_out[2] chany_top_out[3]
+ chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8]
+ chany_top_out[9] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_ left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
+ left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_ left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
+ pReset prog_clk right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
+ right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_ right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
+ top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_ top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
+ vccd1 vssd1 vssd1_uq0 vccd1_uq0
XFILLER_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1270_ net13 vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0985_ _0160_ vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__inv_2
XFILLER_8_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1606_ mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out _0449_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out
+ sky130_fd_sc_hd__ebufn_2
X_1537_ mux_left_track_9.INVTX1_9_.out _0380_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1468_ mux_bottom_track_1.INVTX1_4_.out _0311_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1399_ mux_bottom_track_1.INVTX1_1_.out _0242_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_63_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0770_ mem_top_track_16.DFFR_0_.D vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__inv_2
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1322_ net55 vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__clkbuf_1
X_1253_ net30 vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1184_ clknet_4_8_0_prog_clk mem_left_track_9.DFFR_4_.Q _0106_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_9.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
X_0968_ _0159_ vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__inv_2
XFILLER_20_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0899_ net28 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.INVTX1_3_.out sky130_fd_sc_hd__inv_2
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0822_ net67 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.INVTX1_2_.out sky130_fd_sc_hd__inv_2
XFILLER_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0684_ mem_right_track_24.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__inv_2
X_0753_ mem_top_track_16.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__inv_2
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1305_ net63 vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1167_ clknet_4_1_0_prog_clk mem_bottom_track_25.DFFR_5_.Q _0089_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_25.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
X_1098_ clknet_4_3_0_prog_clk mem_top_track_16.DFFR_2_.Q _0020_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_16.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1021_ _0152_ vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__buf_4
X_0805_ mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1 vccd1
+ vccd1 mux_right_track_0.out sky130_fd_sc_hd__inv_2
X_0667_ mem_bottom_track_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__inv_2
X_0736_ mem_top_track_24.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__inv_2
X_0598_ mem_left_track_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__inv_2
XFILLER_55_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1219_ clknet_4_4_0_prog_clk mem_bottom_track_33.DFFR_3_.Q _0141_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_33.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1570_ mux_left_track_25.INVTX1_10_.out _0413_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_0521_ mem_bottom_track_1.DFFR_0_.D vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__inv_2
XANTENNA_5 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1004_ _0162_ vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__inv_2
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0719_ mem_right_track_0.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__inv_2
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 chanx_left_out[10] sky130_fd_sc_hd__buf_2
XFILLER_16_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1622_ mux_bottom_track_33.INVTX1_3_.out _0465_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1484_ mux_bottom_track_9.INVTX1_4_.out _0327_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1553_ mux_left_track_17.INVTX1_9_.out _0396_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0504_ mem_left_track_33.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__inv_2
XFILLER_52_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0984_ _0160_ vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__inv_2
X_1536_ net185 _0379_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
X_1605_ mux_bottom_track_33.INVTX1_0_.out _0448_ vssd1 vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1467_ mux_bottom_track_1.INVTX1_8_.out _0310_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1398_ mux_left_track_1.INVTX1_9_.out _0241_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_6_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_6_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_49_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1321_ mux_top_track_8.out vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__clkbuf_1
X_1252_ mux_left_track_33.out vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1183_ clknet_4_8_0_prog_clk mem_left_track_9.DFFR_5_.Q _0105_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_9.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0967_ _0159_ vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__inv_2
XFILLER_32_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0898_ net34 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.INVTX1_4_.out sky130_fd_sc_hd__inv_2
X_1519_ mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out _0362_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_23_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0821_ net25 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.INVTX1_3_.out sky130_fd_sc_hd__inv_2
XFILLER_9_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0752_ mem_top_track_16.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__inv_2
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0683_ mem_right_track_24.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__inv_2
X_1166_ clknet_4_0_0_prog_clk mem_bottom_track_25.DFFR_6_.Q _0088_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_25.DFFR_7_.Q sky130_fd_sc_hd__dfrtp_1
X_1304_ net73 vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__clkbuf_2
XFILLER_52_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1097_ clknet_4_1_0_prog_clk mem_top_track_16.DFFR_3_.Q _0019_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_16.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1020_ _0163_ vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__inv_2
XFILLER_61_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0735_ mem_top_track_24.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__inv_2
X_0804_ net94 vssd1 vssd1 vccd1 vccd1 mux_top_track_24.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_1504__183 vssd1 vssd1 vccd1 vccd1 net183 _1504__183/LO sky130_fd_sc_hd__conb_1
XFILLER_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0666_ mem_bottom_track_1.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__inv_2
X_0597_ mem_left_track_1.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__inv_2
XFILLER_52_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1149_ clknet_4_15_0_prog_clk mem_bottom_track_1.DFFR_0_.D _0071_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_1.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_1_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1218_ clknet_4_1_0_prog_clk mem_bottom_track_33.DFFR_4_.Q _0140_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_33.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_52_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_6 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_ vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0520_ mem_right_track_32.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__inv_2
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1003_ _0162_ vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__inv_2
XFILLER_22_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0718_ mem_right_track_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__inv_2
XFILLER_57_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0649_ mem_bottom_track_9.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__inv_2
XFILLER_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 chanx_left_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1552_ net186 _0395_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
X_1621_ net191 _0464_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1483_ mux_bottom_track_9.INVTX1_8_.out _0326_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_39_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0503_ mem_left_track_33.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__inv_2
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0983_ _0160_ vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__inv_2
X_1535_ mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out _0378_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1604_ mux_left_track_33.INVTX1_5_.out _0447_ vssd1 vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1466_ mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out _0309_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
X_1397_ mux_left_track_1.INVTX1_8_.out _0240_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_50_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1320_ net57 vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1251_ net32 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1182_ clknet_4_2_0_prog_clk mem_left_track_9.DFFR_6_.Q _0104_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_17.DFFR_0_.D sky130_fd_sc_hd__dfrtp_1
XFILLER_64_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0897_ net18 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.INVTX1_5_.out sky130_fd_sc_hd__inv_2
X_0966_ _0153_ vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__buf_4
XFILLER_59_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1449_ mux_bottom_track_25.INVTX1_2_.out _0292_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1518_ mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out _0361_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_4_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0820_ net40 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.INVTX1_4_.out sky130_fd_sc_hd__inv_2
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0751_ mem_top_track_16.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__inv_2
X_1303_ net74 vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0682_ mem_right_track_24.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__inv_2
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1165_ clknet_4_9_0_prog_clk mem_bottom_track_17.DFFR_0_.D _0087_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_17.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
X_1096_ clknet_4_0_0_prog_clk mem_top_track_16.DFFR_4_.Q _0018_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_16.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0949_ _0157_ vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__inv_2
XFILLER_18_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0803_ mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1 vccd1
+ vccd1 mux_top_track_24.out sky130_fd_sc_hd__clkinv_2
X_0665_ mem_bottom_track_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__inv_2
X_0734_ mem_top_track_24.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__inv_2
X_0596_ mem_left_track_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__inv_2
XFILLER_52_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1079_ clknet_4_0_0_prog_clk mem_top_track_0.DFFR_5_.Q _0001_ vssd1 vssd1 vccd1 vccd1
+ mem_top_track_0.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
X_1148_ clknet_4_7_0_prog_clk mem_bottom_track_1.DFFR_0_.Q _0070_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_1.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
X_1217_ clknet_4_7_0_prog_clk mem_right_track_24.DFFR_7_.Q _0139_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_32.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_7 chany_bottom_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1002_ _0162_ vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__inv_2
XFILLER_34_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0648_ mem_bottom_track_9.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__inv_2
X_0717_ mem_right_track_0.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__inv_2
XFILLER_57_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0579_ mem_left_track_9.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__inv_2
XFILLER_40_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 chanx_left_out[12] sky130_fd_sc_hd__buf_2
XFILLER_48_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1482_ mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out _0325_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
X_1551_ mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out _0394_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
X_0502_ mem_left_track_33.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__inv_2
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1620_ mux_left_track_33.INVTX1_7_.out _0463_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_39_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0982_ _0160_ vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__inv_2
X_1534_ mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out _0377_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
X_1603_ mux_bottom_track_33.INVTX1_6_.out _0446_ vssd1 vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1465_ mux_bottom_track_1.INVTX1_3_.out _0308_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1396_ mux_left_track_1.INVTX1_7_.out _0239_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1250_ net33 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__clkbuf_2
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1181_ clknet_4_4_0_prog_clk mem_bottom_track_33.DFFR_5_.Q _0103_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_1.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0965_ _0158_ vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__inv_2
X_0896_ net20 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.INVTX1_6_.out sky130_fd_sc_hd__inv_2
XFILLER_55_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1448_ mux_left_track_25.INVTX1_2_.out _0291_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1517_ mux_bottom_track_25.INVTX1_0_.out _0360_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1379_ mux_bottom_track_25.INVTX1_10_.out _0222_ vssd1 vssd1 vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_23_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0681_ mem_right_track_24.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__inv_2
X_0750_ mem_top_track_16.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__inv_2
X_1302_ mux_bottom_track_9.out vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__clkbuf_1
XFILLER_56_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1392__176 vssd1 vssd1 vccd1 vccd1 net176 _1392__176/LO sky130_fd_sc_hd__conb_1
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1164_ clknet_4_14_0_prog_clk mem_bottom_track_17.DFFR_0_.Q _0086_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_17.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
X_1095_ clknet_4_1_0_prog_clk mem_top_track_16.DFFR_5_.Q _0017_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_16.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
X_0948_ _0157_ vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__inv_2
X_0879_ mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_17.out sky130_fd_sc_hd__inv_2
XFILLER_28_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0802_ net93 vssd1 vssd1 vccd1 vccd1 mux_top_track_16.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0664_ mem_bottom_track_1.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__inv_2
X_0733_ mem_top_track_24.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__inv_2
XFILLER_29_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1216_ clknet_4_6_0_prog_clk mem_right_track_32.DFFR_0_.Q _0138_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_32.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
X_0595_ mem_left_track_1.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__inv_2
XFILLER_52_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1147_ clknet_4_5_0_prog_clk mem_bottom_track_1.DFFR_1_.Q _0069_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_1.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
X_1078_ clknet_4_2_0_prog_clk mem_top_track_0.DFFR_6_.Q _0000_ vssd1 vssd1 vccd1 vccd1
+ mem_top_track_0.DFFR_7_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_8 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_ vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1001_ _0162_ vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__inv_2
XFILLER_34_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0578_ mem_left_track_17.DFFR_0_.D vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__inv_2
X_0647_ mem_bottom_track_9.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__inv_2
X_0716_ mem_right_track_8.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__inv_2
XFILLER_57_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1481_ mux_bottom_track_9.INVTX1_3_.out _0324_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1550_ mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out _0393_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0501_ mem_left_track_33.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__inv_2
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0981_ _0160_ vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__inv_2
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1602_ mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out _0445_ vssd1
+ vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1533_ mux_bottom_track_1.INVTX1_0_.out _0376_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1395_ mux_bottom_track_1.INVTX1_11_.out _0238_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1464_ mux_bottom_track_1.INVTX1_2_.out _0307_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_23_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1180_ clknet_4_6_0_prog_clk mem_left_track_1.DFFR_0_.Q _0102_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_1.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
X_0964_ _0158_ vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__inv_2
XFILLER_32_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1516_ mux_bottom_track_25.INVTX1_4_.out _0359_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_0895_ mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out vssd1 vssd1
+ vccd1 vccd1 mux_bottom_track_33.out sky130_fd_sc_hd__inv_2
XFILLER_55_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1447_ mux_bottom_track_25.INVTX1_1_.out _0290_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1378_ mux_bottom_track_9.INVTX1_10_.out _0221_ vssd1 vssd1 vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0680_ mem_right_track_24.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__inv_2
XFILLER_64_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1301_ net76 vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__clkbuf_2
X_1163_ clknet_4_9_0_prog_clk mem_bottom_track_17.DFFR_1_.Q _0085_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_17.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
X_1094_ clknet_4_1_0_prog_clk mem_top_track_16.DFFR_6_.Q _0016_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_16.DFFR_7_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0947_ _0157_ vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__inv_2
X_0878_ net85 vssd1 vssd1 vccd1 vccd1 mux_left_track_9.INVTX1_11_.out sky130_fd_sc_hd__inv_2
XFILLER_43_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_5_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_5_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0801_ mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1 vccd1
+ vccd1 mux_top_track_16.out sky130_fd_sc_hd__inv_2
X_0594_ mem_left_track_1.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__inv_2
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0663_ mem_bottom_track_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__inv_2
X_0732_ mem_right_track_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__inv_2
XFILLER_37_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1146_ clknet_4_1_0_prog_clk mem_bottom_track_1.DFFR_2_.Q _0068_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_1.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
X_1215_ clknet_4_5_0_prog_clk mem_right_track_32.DFFR_1_.Q _0137_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_32.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_52_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1077_ _0153_ vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__inv_2
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_9 top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_ vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_1000_ _0162_ vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__inv_2
XFILLER_19_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0715_ mem_right_track_8.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__inv_2
XFILLER_57_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0646_ mem_bottom_track_9.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__inv_2
X_0577_ mem_left_track_9.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__inv_2
X_1129_ clknet_4_11_0_prog_clk mem_right_track_16.DFFR_3_.Q _0051_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_16.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1480_ mux_bottom_track_9.INVTX1_2_.out _0323_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0500_ mem_left_track_33.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__inv_2
XFILLER_22_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0629_ mem_bottom_track_17.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__inv_2
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0980_ _0160_ vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__inv_2
X_1601_ mux_left_track_17.INVTX1_2_.out _0444_ vssd1 vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1532_ mux_bottom_track_1.INVTX1_3_.out _0375_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1394_ mux_bottom_track_1.INVTX1_9_.out _0237_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1463_ mux_bottom_track_1.INVTX1_1_.out _0306_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_35_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0894_ mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out vssd1 vssd1 vccd1
+ vccd1 mux_right_track_32.out sky130_fd_sc_hd__inv_2
XFILLER_32_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0963_ _0158_ vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__inv_2
XFILLER_59_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1515_ mux_bottom_track_25.INVTX1_8_.out _0358_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_55_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1377_ mux_bottom_track_25.INVTX1_9_.out _0220_ vssd1 vssd1 vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1446_ mux_left_track_25.INVTX1_8_.out _0289_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_4_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1162_ clknet_4_8_0_prog_clk mem_bottom_track_17.DFFR_2_.Q _0084_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_17.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
X_1300_ net77 vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1093_ clknet_4_10_0_prog_clk mem_top_track_0.DFFR_7_.Q _0015_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_8.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1440__179 vssd1 vssd1 vccd1 vccd1 net179 _1440__179/LO sky130_fd_sc_hd__conb_1
XFILLER_20_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0946_ _0157_ vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__inv_2
X_0877_ net72 vssd1 vssd1 vccd1 vccd1 mux_left_track_9.INVTX1_3_.out sky130_fd_sc_hd__inv_2
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1429_ mux_left_track_17.INVTX1_8_.out _0272_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0800_ net92 vssd1 vssd1 vccd1 vccd1 mux_top_track_8.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0731_ mem_right_track_0.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__inv_2
X_0662_ mem_bottom_track_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__inv_2
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0593_ mem_left_track_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__inv_2
XFILLER_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1145_ clknet_4_0_0_prog_clk mem_bottom_track_1.DFFR_3_.Q _0067_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_1.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_2
X_1214_ clknet_4_6_0_prog_clk mem_right_track_32.DFFR_2_.Q _0136_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_32.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1076_ _0153_ vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__inv_2
X_0929_ _0155_ vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__inv_2
XFILLER_20_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0714_ mem_right_track_8.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__inv_2
X_0645_ mem_bottom_track_9.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__inv_2
XFILLER_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0576_ mem_left_track_9.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__inv_2
X_1128_ clknet_4_11_0_prog_clk mem_right_track_16.DFFR_4_.Q _0050_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_16.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1059_ _0167_ vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__inv_2
XFILLER_0_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0628_ mem_bottom_track_17.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__inv_2
XFILLER_7_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0559_ mem_left_track_17.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__inv_2
XFILLER_21_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1600_ mux_bottom_track_33.INVTX1_1_.out _0443_ vssd1 vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1531_ mux_left_track_1.INVTX1_8_.out _0374_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1462_ mux_bottom_track_1.INVTX1_7_.out _0305_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1393_ mux_bottom_track_1.INVTX1_8_.out _0236_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_50_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0962_ _0158_ vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__inv_2
X_0893_ mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out vssd1 vssd1 vccd1
+ vccd1 mux_top_track_32.out sky130_fd_sc_hd__inv_2
X_1445_ mux_left_track_25.INVTX1_7_.out _0288_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1514_ mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out _0357_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1376_ net175 _0219_ vssd1 vssd1 vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_23_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1472__181 vssd1 vssd1 vccd1 vccd1 net181 _1472__181/LO sky130_fd_sc_hd__conb_1
XFILLER_50_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1161_ clknet_4_11_0_prog_clk mem_bottom_track_17.DFFR_3_.Q _0083_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_17.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
X_1092_ clknet_4_10_0_prog_clk mem_top_track_8.DFFR_0_.Q _0014_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_8.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
X_0876_ net54 vssd1 vssd1 vccd1 vccd1 mux_left_track_9.INVTX1_7_.out sky130_fd_sc_hd__inv_2
X_0945_ _0157_ vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__inv_2
XFILLER_9_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1428_ mux_left_track_17.INVTX1_7_.out _0271_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_18_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1359_ mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out _0202_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_51_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0661_ mem_bottom_track_1.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__inv_2
XFILLER_6_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0730_ mem_right_track_0.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__inv_2
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0592_ mem_left_track_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__inv_2
X_1213_ clknet_4_3_0_prog_clk mem_right_track_32.DFFR_3_.Q _0135_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_32.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
X_1075_ _0168_ vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__inv_2
X_1144_ clknet_4_0_0_prog_clk mem_bottom_track_1.DFFR_4_.Q _0066_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_1.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0928_ _0155_ vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__inv_2
X_0859_ net38 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.INVTX1_4_.out sky130_fd_sc_hd__inv_2
XFILLER_28_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0713_ mem_right_track_8.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__inv_2
X_0644_ mem_bottom_track_9.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__inv_2
X_0575_ mem_left_track_9.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__inv_2
X_1127_ clknet_4_14_0_prog_clk mem_right_track_16.DFFR_5_.Q _0049_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_16.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1058_ _0167_ vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__inv_2
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0558_ mem_left_track_17.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__inv_2
X_0627_ mem_bottom_track_17.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__inv_2
XFILLER_53_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1530_ mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out _0373_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
X_1461_ mux_bottom_track_1.INVTX1_6_.out _0304_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1392_ net176 _0235_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_4_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0961_ _0158_ vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__inv_2
XFILLER_27_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0892_ net83 vssd1 vssd1 vccd1 vccd1 mux_left_track_25.INVTX1_11_.out sky130_fd_sc_hd__inv_2
XFILLER_40_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1513_ mux_bottom_track_25.INVTX1_3_.out _0356_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1375_ mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out _0218_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
X_1444_ mux_left_track_9.INVTX1_8_.out _0287_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_4_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1160_ clknet_4_10_0_prog_clk mem_bottom_track_17.DFFR_4_.Q _0082_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_17.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_37_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1091_ clknet_4_9_0_prog_clk mem_top_track_8.DFFR_1_.Q _0013_ vssd1 vssd1 vccd1 vccd1
+ mem_top_track_8.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0944_ _0153_ vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__buf_4
X_0875_ net56 vssd1 vssd1 vccd1 vccd1 mux_left_track_9.INVTX1_8_.out sky130_fd_sc_hd__inv_2
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1427_ mux_bottom_track_17.INVTX1_11_.out _0270_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_28_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1358_ mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out _0201_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_63_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1289_ net70 vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0660_ mem_bottom_track_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__inv_2
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0591_ mem_left_track_1.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__inv_2
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1212_ clknet_4_13_0_prog_clk mem_right_track_32.DFFR_4_.Q _0134_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_1.DFFR_0_.D sky130_fd_sc_hd__dfrtp_1
XFILLER_52_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1074_ _0168_ vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__inv_2
X_1143_ clknet_4_0_0_prog_clk mem_bottom_track_1.DFFR_5_.Q _0065_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_1.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0927_ _0155_ vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__inv_2
XFILLER_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0789_ mem_top_track_0.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__inv_2
X_0858_ net26 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.INVTX1_5_.out sky130_fd_sc_hd__inv_2
XFILLER_45_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0712_ mem_right_track_8.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__inv_2
X_0643_ mem_bottom_track_9.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__inv_2
Xclkbuf_4_4_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_4_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
X_0574_ mem_left_track_9.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__inv_2
X_1126_ clknet_4_11_0_prog_clk mem_right_track_16.DFFR_6_.Q _0048_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_16.DFFR_7_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1057_ _0167_ vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__inv_2
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0626_ mem_bottom_track_17.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__inv_2
X_0557_ mem_left_track_17.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0405_ sky130_fd_sc_hd__inv_2
X_1109_ clknet_4_5_0_prog_clk mem_top_track_16.DFFR_7_.Q _0031_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_24.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1460_ mux_bottom_track_1.INVTX1_5_.out _0303_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1391_ mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out _0234_ vssd1 vssd1
+ vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_50_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0609_ mem_bottom_track_25.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__inv_2
X_1589_ mux_bottom_track_33.INVTX1_3_.out _0432_ vssd1 vssd1 vccd1 vccd1 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_53_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0960_ _0158_ vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__inv_2
XFILLER_32_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0891_ net65 vssd1 vssd1 vccd1 vccd1 mux_left_track_25.INVTX1_2_.out sky130_fd_sc_hd__inv_2
X_1512_ mux_bottom_track_25.INVTX1_2_.out _0355_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1443_ mux_bottom_track_25.INVTX1_10_.out _0286_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1374_ mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out _0217_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1090_ clknet_4_12_0_prog_clk mem_top_track_8.DFFR_2_.Q _0012_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_8.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
X_1520__184 vssd1 vssd1 vccd1 vccd1 net184 _1520__184/LO sky130_fd_sc_hd__conb_1
X_0874_ net61 vssd1 vssd1 vccd1 vccd1 mux_left_track_9.INVTX1_9_.out sky130_fd_sc_hd__inv_2
X_0943_ _0156_ vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__inv_2
XFILLER_9_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1357_ mux_top_track_8.INVTX1_0_.out _0200_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1288_ net71 vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__clkbuf_2
X_1426_ mux_bottom_track_17.INVTX1_9_.out _0269_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0590_ mem_left_track_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__inv_2
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1211_ clknet_4_12_0_prog_clk mem_top_track_24.DFFR_7_.Q _0133_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_32.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
X_1142_ clknet_4_2_0_prog_clk mem_bottom_track_1.DFFR_6_.Q _0064_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_1.DFFR_7_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1073_ _0168_ vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__inv_2
XFILLER_18_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0926_ _0155_ vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__inv_2
X_0857_ net33 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.INVTX1_6_.out sky130_fd_sc_hd__inv_2
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0788_ mem_top_track_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__inv_2
X_1409_ mux_bottom_track_9.INVTX1_8_.out _0252_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_56_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0711_ mem_right_track_8.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__inv_2
XFILLER_42_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0642_ mem_bottom_track_17.DFFR_0_.D vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__inv_2
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0573_ mem_left_track_9.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__inv_2
XFILLER_38_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1125_ clknet_4_7_0_prog_clk mem_right_track_0.DFFR_7_.Q _0047_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_8.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1056_ _0167_ vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__inv_2
XFILLER_15_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0909_ net86 vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0625_ mem_bottom_track_17.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__inv_2
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0556_ mem_left_track_25.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__inv_2
XFILLER_53_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1039_ _0165_ vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__inv_2
X_1108_ clknet_4_5_0_prog_clk mem_top_track_24.DFFR_0_.Q _0030_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_24.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1390_ mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out _0233_ vssd1 vssd1
+ vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_35_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0608_ mem_bottom_track_25.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__inv_2
X_1588_ mux_bottom_track_33.INVTX1_2_.out _0431_ vssd1 vssd1 vccd1 vccd1 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0539_ mem_top_track_32.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__inv_2
XFILLER_53_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0890_ net57 vssd1 vssd1 vccd1 vccd1 mux_left_track_25.INVTX1_7_.out sky130_fd_sc_hd__inv_2
X_1511_ mux_bottom_track_25.INVTX1_1_.out _0354_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1442_ mux_bottom_track_25.INVTX1_9_.out _0285_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_4_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1373_ mux_top_track_16.INVTX1_0_.out _0216_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_63_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0873_ net49 vssd1 vssd1 vccd1 vccd1 mux_left_track_9.INVTX1_10_.out sky130_fd_sc_hd__inv_2
XFILLER_20_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0942_ _0156_ vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__inv_2
XFILLER_9_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1425_ mux_bottom_track_17.INVTX1_8_.out _0268_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_55_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1356_ mux_bottom_track_9.INVTX1_6_.out _0199_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1287_ mux_right_track_0.out vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__clkbuf_1
XFILLER_11_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1141_ clknet_4_9_0_prog_clk mem_right_track_16.DFFR_7_.Q _0063_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_24.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
X_1210_ clknet_4_3_0_prog_clk mem_top_track_32.DFFR_0_.Q _0132_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_32.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
X_1072_ _0168_ vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__inv_2
XFILLER_18_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0787_ mem_top_track_0.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__inv_2
X_0925_ _0155_ vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__inv_2
X_0856_ net2 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.INVTX1_7_.out sky130_fd_sc_hd__inv_2
X_1408_ net177 _0251_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
X_1339_ mux_bottom_track_1.INVTX1_8_.out _0182_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_28_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0710_ mem_right_track_8.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__inv_2
X_0641_ mem_bottom_track_9.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__inv_2
X_0572_ mem_left_track_17.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__inv_2
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1124_ clknet_4_15_0_prog_clk mem_right_track_8.DFFR_0_.Q _0046_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_8.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
X_1055_ _0167_ vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__inv_2
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0839_ mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1
+ vccd1 vccd1 mux_bottom_track_17.out sky130_fd_sc_hd__inv_2
X_0908_ net50 vssd1 vssd1 vccd1 vccd1 mux_left_track_33.INVTX1_7_.out sky130_fd_sc_hd__inv_2
XFILLER_56_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0624_ mem_bottom_track_17.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__inv_2
X_0555_ mem_left_track_25.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__inv_2
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1038_ _0165_ vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__inv_2
X_1107_ clknet_4_7_0_prog_clk mem_top_track_24.DFFR_1_.Q _0029_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_24.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0607_ mem_bottom_track_25.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__inv_2
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0538_ mem_top_track_32.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__inv_2
X_1587_ mux_bottom_track_33.INVTX1_6_.out _0430_ vssd1 vssd1 vccd1 vccd1 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1441_ mux_bottom_track_25.INVTX1_8_.out _0284_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1510_ mux_bottom_track_25.INVTX1_7_.out _0353_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_4_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1372_ mux_bottom_track_17.INVTX1_6_.out _0215_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_4_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0941_ _0156_ vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__inv_2
X_0872_ mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_9.out sky130_fd_sc_hd__clkinv_2
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1355_ mux_bottom_track_9.INVTX1_8_.out _0198_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1424_ net178 _0267_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_55_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1286_ net6 vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__clkbuf_2
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1071_ _0168_ vssd1 vssd1 vccd1 vccd1 _0145_ sky130_fd_sc_hd__inv_2
X_1140_ clknet_4_3_0_prog_clk mem_right_track_24.DFFR_0_.Q _0062_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_24.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0924_ _0155_ vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__inv_2
XFILLER_33_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0786_ mem_top_track_0.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__inv_2
X_0855_ net19 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.INVTX1_8_.out sky130_fd_sc_hd__inv_2
X_1407_ mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out _0250_ vssd1 vssd1
+ vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
X_1338_ mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out _0181_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_51_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1269_ net14 vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0571_ mem_left_track_17.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__inv_2
X_0640_ mem_bottom_track_9.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__inv_2
XFILLER_2_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1123_ clknet_4_8_0_prog_clk mem_right_track_8.DFFR_1_.Q _0045_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_8.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
X_1054_ _0152_ vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__buf_4
X_0907_ net79 vssd1 vssd1 vccd1 vccd1 mux_left_track_33.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_0769_ mem_top_track_8.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__inv_2
X_0838_ net11 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.INVTX1_11_.out sky130_fd_sc_hd__inv_2
XFILLER_56_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0623_ mem_bottom_track_17.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__inv_2
X_0554_ mem_left_track_25.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__inv_2
X_1106_ clknet_4_7_0_prog_clk mem_top_track_24.DFFR_2_.Q _0028_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_24.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1037_ _0165_ vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__inv_2
Xinput90 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_ vssd1 vssd1 vccd1
+ vccd1 net90 sky130_fd_sc_hd__clkbuf_1
XFILLER_21_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_3_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_3_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_8_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0606_ mem_bottom_track_25.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__inv_2
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1586_ mux_left_track_33.INVTX1_6_.out _0429_ vssd1 vssd1 vccd1 vccd1 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
X_0537_ mem_top_track_32.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__inv_2
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1371_ mux_bottom_track_17.INVTX1_8_.out _0214_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1440_ net179 _0283_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_4_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1569_ mux_left_track_25.INVTX1_9_.out _0412_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0940_ _0156_ vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__inv_2
XFILLER_13_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0871_ net84 vssd1 vssd1 vccd1 vccd1 mux_left_track_1.INVTX1_11_.out sky130_fd_sc_hd__inv_2
XFILLER_9_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1423_ mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out _0266_ vssd1
+ vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_2
X_1354_ mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out _0197_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
X_1285_ net16 vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__clkbuf_2
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1488__182 vssd1 vssd1 vccd1 vccd1 net182 _1488__182/LO sky130_fd_sc_hd__conb_1
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1070_ _0168_ vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__inv_2
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0854_ net7 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.INVTX1_9_.out sky130_fd_sc_hd__inv_2
X_0923_ _0155_ vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__inv_2
X_0785_ mem_top_track_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__inv_2
X_1268_ mux_left_track_1.out vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__clkbuf_1
X_1337_ mux_bottom_track_17.INVTX1_4_.out _0180_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1406_ mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out _0249_ vssd1 vssd1
+ vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_61_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1199_ clknet_4_11_0_prog_clk mem_left_track_25.DFFR_5_.Q _0121_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_25.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_36_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0570_ mem_left_track_17.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__inv_2
X_1122_ clknet_4_9_0_prog_clk mem_right_track_8.DFFR_2_.Q _0044_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_8.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1053_ _0166_ vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__inv_2
XFILLER_18_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0837_ net73 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0906_ net58 vssd1 vssd1 vccd1 vccd1 mux_left_track_33.INVTX1_5_.out sky130_fd_sc_hd__inv_2
X_0768_ mem_top_track_8.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__inv_2
X_0699_ mem_right_track_16.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__inv_2
XFILLER_56_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0553_ mem_left_track_25.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__inv_2
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0622_ mem_bottom_track_17.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__inv_2
XFILLER_53_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1105_ clknet_4_9_0_prog_clk mem_top_track_24.DFFR_3_.Q _0027_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_24.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1036_ _0165_ vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__inv_2
XFILLER_21_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput91 top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_ vssd1 vssd1 vccd1
+ vccd1 net91 sky130_fd_sc_hd__clkbuf_1
Xinput80 chany_top_in[8] vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__clkbuf_1
XFILLER_44_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1585_ net188 _0428_ vssd1 vssd1 vccd1 vccd1 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
X_0536_ mem_top_track_32.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__inv_2
X_0605_ mem_bottom_track_25.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__inv_2
XFILLER_53_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1019_ _0163_ vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__inv_2
XFILLER_57_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1370_ mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out _0213_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_48_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1568_ net187 _0411_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1499_ mux_bottom_track_17.INVTX1_8_.out _0342_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_39_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0519_ mem_right_track_32.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__inv_2
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0870_ net75 vssd1 vssd1 vccd1 vccd1 mux_left_track_1.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XFILLER_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1422_ mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out _0265_ vssd1
+ vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_2
X_1353_ mux_bottom_track_9.INVTX1_5_.out _0196_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1284_ net17 vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0999_ _0152_ vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__buf_4
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0853_ net14 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.INVTX1_10_.out sky130_fd_sc_hd__inv_2
X_0922_ _0153_ vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__buf_4
X_0784_ mem_top_track_0.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__inv_2
X_1405_ mux_bottom_track_1.INVTX1_0_.out _0248_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
Xinput1 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_ vssd1 vssd1 vccd1
+ vccd1 net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_45_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1198_ clknet_4_14_0_prog_clk mem_left_track_25.DFFR_6_.Q _0120_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_25.DFFR_7_.Q sky130_fd_sc_hd__dfrtp_1
X_1336_ mux_bottom_track_1.INVTX1_4_.out _0179_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_36_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1267_ net25 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_2
XFILLER_51_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0_prog_clk prog_clk vssd1 vssd1 vccd1 vccd1 clknet_0_prog_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_59_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1121_ clknet_4_10_0_prog_clk mem_right_track_8.DFFR_3_.Q _0043_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_8.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1052_ _0166_ vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__inv_2
XFILLER_21_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0767_ mem_top_track_8.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__inv_2
X_0905_ net47 vssd1 vssd1 vccd1 vccd1 mux_left_track_33.INVTX1_6_.out sky130_fd_sc_hd__inv_2
X_0836_ net80 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0698_ mem_right_track_16.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__inv_2
XFILLER_29_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1319_ net58 vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__clkbuf_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0621_ mem_bottom_track_17.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__inv_2
XFILLER_7_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0552_ mem_left_track_25.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__inv_2
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1035_ _0165_ vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__inv_2
X_1104_ clknet_4_13_0_prog_clk mem_top_track_24.DFFR_4_.Q _0026_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_24.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_61_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput92 top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_ vssd1 vssd1 vccd1
+ vccd1 net92 sky130_fd_sc_hd__clkbuf_1
Xinput81 chany_top_in[9] vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__clkbuf_1
Xinput70 chany_top_in[16] vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__clkbuf_2
X_0819_ net29 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.INVTX1_5_.out sky130_fd_sc_hd__inv_2
XFILLER_37_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1584_ mux_bottom_track_33.INVTX1_7_.out _0427_ vssd1 vssd1 vccd1 vccd1 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
X_0604_ mem_left_track_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__inv_2
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0535_ mem_top_track_32.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__inv_2
XFILLER_34_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1018_ _0163_ vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__inv_2
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1567_ mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out _0410_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
X_0518_ mem_right_track_32.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__inv_2
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1498_ mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out _0341_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1421_ mux_bottom_track_9.INVTX1_0_.out _0264_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1352_ mux_bottom_track_9.INVTX1_4_.out _0195_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1283_ mux_right_track_8.out vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0998_ _0161_ vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__inv_2
X_1536__185 vssd1 vssd1 vccd1 vccd1 net185 _1536__185/LO sky130_fd_sc_hd__conb_1
X_1619_ mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out _0462_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0921_ _0154_ vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__inv_2
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0783_ mem_top_track_0.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__inv_2
X_0852_ mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1
+ vccd1 vccd1 mux_bottom_track_25.out sky130_fd_sc_hd__inv_2
X_1404_ mux_right_track_0.INVTX1_4_.out _0247_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1335_ mux_bottom_track_1.INVTX1_3_.out _0178_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1266_ net35 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1197_ clknet_4_8_0_prog_clk mem_left_track_17.DFFR_0_.D _0119_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_17.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_2
Xinput2 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_ vssd1 vssd1 vccd1
+ vccd1 net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1328__172 vssd1 vssd1 vccd1 vccd1 net172 _1328__172/LO sky130_fd_sc_hd__conb_1
XFILLER_27_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1051_ _0166_ vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__inv_2
X_1120_ clknet_4_10_0_prog_clk mem_right_track_8.DFFR_4_.Q _0042_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_8.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0904_ mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_33.out sky130_fd_sc_hd__inv_2
X_0766_ mem_top_track_8.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__inv_2
X_0697_ mem_right_track_16.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__inv_2
X_0835_ net68 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.INVTX1_2_.out sky130_fd_sc_hd__inv_2
X_1318_ net59 vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_1
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0551_ mem_left_track_25.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0412_ sky130_fd_sc_hd__inv_2
X_0620_ mem_bottom_track_25.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__inv_2
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1103_ clknet_4_12_0_prog_clk mem_top_track_24.DFFR_5_.Q _0025_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_24.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
X_1034_ _0165_ vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__inv_2
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput71 chany_top_in[17] vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__clkbuf_2
X_0818_ net31 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.INVTX1_6_.out sky130_fd_sc_hd__inv_2
X_0749_ mem_top_track_16.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__inv_2
Xinput93 top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_ vssd1 vssd1 vccd1
+ vccd1 net93 sky130_fd_sc_hd__clkbuf_1
Xinput60 chany_bottom_in[7] vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_1
Xinput82 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_ vssd1 vssd1 vccd1
+ vccd1 net82 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0534_ mem_top_track_32.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__inv_2
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1583_ mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out _0426_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_4
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0603_ mem_left_track_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__inv_2
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1017_ _0163_ vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__inv_2
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_2_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_2_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
X_0517_ mem_right_track_32.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__inv_2
X_1566_ mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out _0409_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1497_ mux_bottom_track_17.INVTX1_3_.out _0340_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1420_ mux_right_track_8.INVTX1_4_.out _0263_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1351_ mux_bottom_track_9.INVTX1_3_.out _0194_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1282_ net19 vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__clkbuf_1
XFILLER_63_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0997_ _0161_ vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__inv_2
X_1618_ mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out _0461_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
X_1549_ mux_bottom_track_9.INVTX1_0_.out _0392_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0920_ _0154_ vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__inv_2
X_0851_ net13 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.INVTX1_11_.out sky130_fd_sc_hd__inv_2
X_0782_ mem_top_track_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__inv_2
X_1265_ net36 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__clkbuf_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1334_ mux_left_track_1.INVTX1_9_.out _0177_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1403_ mux_left_track_33.INVTX1_7_.out _0246_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_51_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput3 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_ vssd1 vssd1 vccd1
+ vccd1 net3 sky130_fd_sc_hd__clkbuf_1
X_1196_ clknet_4_2_0_prog_clk mem_left_track_17.DFFR_0_.Q _0118_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_17.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1050_ _0166_ vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__inv_2
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0834_ net35 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.INVTX1_3_.out sky130_fd_sc_hd__inv_2
X_0903_ net9 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.INVTX1_7_.out sky130_fd_sc_hd__inv_2
X_0696_ mem_right_track_16.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__inv_2
X_0765_ mem_top_track_8.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__inv_2
X_1317_ mux_top_track_16.out vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1179_ clknet_4_2_0_prog_clk mem_left_track_1.DFFR_1_.Q _0101_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_1.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_15_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_15_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xoutput170 net170 vssd1 vssd1 vccd1 vccd1 chany_top_out[8] sky130_fd_sc_hd__buf_2
XFILLER_62_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0550_ mem_left_track_25.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__inv_2
XFILLER_7_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1102_ clknet_4_15_0_prog_clk mem_top_track_24.DFFR_6_.Q _0024_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_24.DFFR_7_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1033_ _0165_ vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__inv_2
Xinput50 chany_bottom_in[15] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_1
Xinput72 chany_top_in[18] vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__clkbuf_1
X_0817_ net3 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.INVTX1_7_.out sky130_fd_sc_hd__inv_2
Xinput61 chany_bottom_in[8] vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_2
Xinput83 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_ vssd1 vssd1 vccd1
+ vccd1 net83 sky130_fd_sc_hd__clkbuf_1
X_0679_ mem_right_track_24.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__inv_2
X_0748_ mem_top_track_24.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__inv_2
Xinput94 top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_ vssd1 vssd1 vccd1
+ vccd1 net94 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0533_ mem_right_track_0.DFFR_0_.D vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__inv_2
X_1582_ mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out _0425_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_4
X_0602_ mem_left_track_1.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__inv_2
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1016_ _0163_ vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__inv_2
XFILLER_57_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0516_ mem_bottom_track_33.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__inv_2
X_1565_ mux_bottom_track_17.INVTX1_0_.out _0408_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1496_ mux_bottom_track_17.INVTX1_2_.out _0339_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1350_ mux_left_track_9.INVTX1_10_.out _0193_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1281_ net20 vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__clkbuf_1
XFILLER_63_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0996_ _0161_ vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__inv_2
X_1617_ mux_bottom_track_33.INVTX1_0_.out _0460_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_59_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1548_ mux_bottom_track_9.INVTX1_3_.out _0391_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_39_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1479_ mux_bottom_track_9.INVTX1_1_.out _0322_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_54_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0850_ net74 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0781_ mem_top_track_0.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__inv_2
X_1402_ mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out _0245_ vssd1 vssd1
+ vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
X_1264_ mux_left_track_9.out vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__clkbuf_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1333_ mux_left_track_1.INVTX1_8_.out _0176_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
Xinput4 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_ vssd1 vssd1 vccd1
+ vccd1 net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1195_ clknet_4_3_0_prog_clk mem_left_track_17.DFFR_1_.Q _0117_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_17.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_3_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0979_ _0160_ vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__inv_2
XFILLER_10_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0833_ net42 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.INVTX1_4_.out sky130_fd_sc_hd__inv_2
X_0902_ net77 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0695_ mem_right_track_16.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__inv_2
X_0764_ mem_top_track_16.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__inv_2
X_1316_ net61 vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__clkbuf_2
X_1178_ clknet_4_6_0_prog_clk mem_left_track_1.DFFR_2_.Q _0100_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_1.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_20 mem_bottom_track_25.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput171 net171 vssd1 vssd1 vccd1 vccd1 chany_top_out[9] sky130_fd_sc_hd__buf_2
Xoutput160 net160 vssd1 vssd1 vccd1 vccd1 chany_top_out[16] sky130_fd_sc_hd__buf_2
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1032_ _0152_ vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__buf_4
X_1101_ clknet_4_0_0_prog_clk mem_top_track_16.DFFR_0_.D _0023_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_16.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput40 chanx_right_in[6] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput62 chany_bottom_in[9] vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput51 chany_bottom_in[16] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__dlymetal6s2s_1
X_0816_ net6 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.INVTX1_8_.out sky130_fd_sc_hd__inv_2
X_0747_ mem_top_track_24.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__inv_2
Xinput73 chany_top_in[1] vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__clkbuf_2
Xinput84 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_ vssd1 vssd1 vccd1
+ vccd1 net84 sky130_fd_sc_hd__clkbuf_1
X_0678_ mem_right_track_24.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__inv_2
XFILLER_29_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1581_ mux_bottom_track_25.INVTX1_0_.out _0424_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
X_0601_ mem_left_track_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__inv_2
XFILLER_7_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0532_ mem_top_track_32.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0431_ sky130_fd_sc_hd__inv_2
XFILLER_26_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1015_ _0163_ vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__inv_2
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1564_ mux_bottom_track_17.INVTX1_3_.out _0407_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_58_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0515_ mem_bottom_track_33.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__inv_2
X_1495_ mux_bottom_track_17.INVTX1_1_.out _0338_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1280_ net21 vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__clkbuf_2
XFILLER_63_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0995_ _0161_ vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__inv_2
X_1547_ mux_left_track_9.INVTX1_8_.out _0390_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1616_ mux_bottom_track_33.INVTX1_3_.out _0459_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1478_ mux_bottom_track_9.INVTX1_7_.out _0321_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_54_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0780_ mem_top_track_8.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__inv_2
X_1401_ mux_left_track_9.INVTX1_3_.out _0244_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_36_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1263_ net38 vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__clkbuf_1
Xinput5 ccff_head vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__dlymetal6s2s_1
X_1332_ mux_left_track_1.INVTX1_7_.out _0175_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1194_ clknet_4_2_0_prog_clk mem_left_track_17.DFFR_2_.Q _0116_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_17.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0978_ _0160_ vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__inv_2
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0832_ net27 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.INVTX1_5_.out sky130_fd_sc_hd__inv_2
X_0901_ net66 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_0763_ mem_top_track_16.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__inv_2
X_1315_ net62 vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0694_ mem_right_track_16.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__inv_2
X_1177_ clknet_4_1_0_prog_clk mem_left_track_1.DFFR_3_.Q _0099_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_1.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_21 mem_left_track_25.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_10 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput150 net150 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[7] sky130_fd_sc_hd__buf_2
Xoutput161 net161 vssd1 vssd1 vccd1 vccd1 chany_top_out[17] sky130_fd_sc_hd__buf_2
XFILLER_46_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1031_ _0164_ vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__inv_2
X_1100_ clknet_4_0_0_prog_clk mem_top_track_16.DFFR_0_.Q _0022_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_16.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
Xinput63 chany_top_in[0] vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__clkbuf_2
Xinput41 chanx_right_in[7] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_1
Xinput30 chanx_right_in[14] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput52 chany_bottom_in[17] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__dlymetal6s2s_1
X_0815_ net21 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.INVTX1_9_.out sky130_fd_sc_hd__inv_2
X_0746_ mem_top_track_24.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__inv_2
Xinput85 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_ vssd1 vssd1 vccd1
+ vccd1 net85 sky130_fd_sc_hd__clkbuf_1
Xinput74 chany_top_in[2] vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__clkbuf_2
X_0677_ mem_right_track_24.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__inv_2
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1229_ clknet_4_9_0_prog_clk mem_left_track_25.DFFR_7_.Q _0151_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_33.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_12_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1580_ mux_bottom_track_25.INVTX1_4_.out _0423_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
X_0531_ mem_top_track_32.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__inv_2
X_0600_ mem_left_track_1.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__inv_2
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1014_ _0163_ vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__inv_2
XFILLER_8_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0729_ mem_right_track_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__inv_2
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1494_ mux_bottom_track_17.INVTX1_7_.out _0337_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1563_ mux_left_track_17.INVTX1_8_.out _0406_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0514_ mem_bottom_track_33.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__inv_2
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0994_ _0161_ vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__inv_2
X_1477_ mux_bottom_track_9.INVTX1_6_.out _0320_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1546_ mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out _0389_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1615_ mux_bottom_track_33.INVTX1_6_.out _0458_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_1_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_1_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_41_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1331_ mux_bottom_track_1.INVTX1_11_.out _0174_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1400_ mux_bottom_track_1.INVTX1_2_.out _0243_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
Xinput6 chanx_left_in[0] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_2
X_1262_ net39 vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1193_ clknet_4_3_0_prog_clk mem_left_track_17.DFFR_3_.Q _0115_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_17.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_51_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0977_ _0153_ vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__buf_4
XFILLER_59_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1529_ mux_bottom_track_1.INVTX1_2_.out _0372_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_42_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0900_ net39 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.INVTX1_2_.out sky130_fd_sc_hd__inv_2
X_0693_ mem_right_track_16.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__inv_2
X_0831_ net30 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.INVTX1_6_.out sky130_fd_sc_hd__inv_2
X_0762_ mem_top_track_16.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__inv_2
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1314_ net45 vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1176_ clknet_4_0_0_prog_clk mem_left_track_1.DFFR_4_.Q _0098_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_1.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_11 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 mem_top_track_32.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput140 net140 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[15] sky130_fd_sc_hd__buf_2
Xoutput151 net151 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[8] sky130_fd_sc_hd__buf_2
Xoutput162 net162 vssd1 vssd1 vccd1 vccd1 chany_top_out[18] sky130_fd_sc_hd__buf_2
XFILLER_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1030_ _0164_ vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__inv_2
X_0814_ net22 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.INVTX1_10_.out sky130_fd_sc_hd__inv_2
Xinput31 chanx_right_in[15] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
Xinput20 chanx_left_in[5] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_2
Xinput42 chanx_right_in[8] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__dlymetal6s2s_1
X_0676_ mem_right_track_24.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__inv_2
X_0745_ mem_top_track_24.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__inv_2
Xinput53 chany_bottom_in[18] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_1
Xinput86 pReset vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__clkbuf_1
Xinput64 chany_top_in[10] vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__clkbuf_2
Xinput75 chany_top_in[3] vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__clkbuf_1
X_1228_ clknet_4_2_0_prog_clk mem_left_track_33.DFFR_0_.Q _0150_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_33.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_52_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1159_ clknet_4_10_0_prog_clk mem_bottom_track_17.DFFR_5_.Q _0081_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_17.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_16_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0530_ mem_top_track_32.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__inv_2
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1013_ _0163_ vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__inv_2
Xclkbuf_4_14_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_14_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
X_0659_ mem_bottom_track_1.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__inv_2
X_0728_ mem_right_track_0.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__inv_2
XFILLER_27_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1493_ mux_bottom_track_17.INVTX1_6_.out _0336_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1562_ mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out _0405_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
X_0513_ mem_bottom_track_33.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__inv_2
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0993_ _0161_ vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__inv_2
X_1614_ mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out _0457_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_8_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1476_ mux_bottom_track_9.INVTX1_5_.out _0319_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1545_ mux_left_track_9.INVTX1_3_.out _0388_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_39_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1261_ net40 vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__clkbuf_1
X_1330_ mux_bottom_track_1.INVTX1_9_.out _0173_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_30_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput7 chanx_left_in[10] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_2
X_1192_ clknet_4_9_0_prog_clk mem_left_track_17.DFFR_4_.Q _0114_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_17.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_17_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0976_ _0159_ vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__inv_2
XFILLER_32_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1459_ mux_bottom_track_1.INVTX1_11_.out _0302_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1528_ mux_bottom_track_1.INVTX1_1_.out _0371_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_42_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0830_ net4 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.INVTX1_7_.out sky130_fd_sc_hd__inv_2
XFILLER_14_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0692_ mem_right_track_16.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__inv_2
X_0761_ mem_top_track_16.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__inv_2
X_1313_ mux_top_track_24.out vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1175_ clknet_4_0_0_prog_clk mem_left_track_1.DFFR_5_.Q _0097_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_1.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_23 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0959_ _0158_ vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__inv_2
XFILLER_32_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_12 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput152 net152 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[9] sky130_fd_sc_hd__buf_2
Xoutput141 net141 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[16] sky130_fd_sc_hd__buf_2
Xoutput163 net163 vssd1 vssd1 vccd1 vccd1 chany_top_out[1] sky130_fd_sc_hd__buf_2
Xoutput130 net130 vssd1 vssd1 vccd1 vccd1 chanx_right_out[6] sky130_fd_sc_hd__buf_2
XFILLER_62_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput32 chanx_right_in[16] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_2
Xinput21 chanx_left_in[6] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__dlymetal6s2s_1
X_0813_ mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1 vccd1
+ vccd1 mux_bottom_track_1.out sky130_fd_sc_hd__clkinv_2
Xinput10 chanx_left_in[13] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_2
Xinput43 chanx_right_in[9] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput54 chany_bottom_in[1] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_2
Xinput76 chany_top_in[4] vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput65 chany_top_in[11] vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_1
Xinput87 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_ vssd1 vssd1 vccd1
+ vccd1 net87 sky130_fd_sc_hd__clkbuf_1
X_0675_ mem_right_track_24.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__inv_2
X_0744_ mem_top_track_24.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__inv_2
X_1158_ clknet_4_11_0_prog_clk mem_bottom_track_17.DFFR_6_.Q _0080_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_17.DFFR_7_.Q sky130_fd_sc_hd__dfrtp_1
X_1227_ clknet_4_1_0_prog_clk mem_left_track_33.DFFR_1_.Q _0149_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_33.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_52_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1089_ clknet_4_8_0_prog_clk mem_top_track_8.DFFR_3_.Q _0011_ vssd1 vssd1 vccd1 vccd1
+ mem_top_track_8.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1012_ _0163_ vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__inv_2
XFILLER_34_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0727_ mem_right_track_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__inv_2
X_0658_ mem_bottom_track_1.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__inv_2
X_0589_ mem_left_track_1.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__inv_2
XFILLER_25_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1492_ mux_bottom_track_17.INVTX1_5_.out _0335_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_0512_ mem_bottom_track_33.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__inv_2
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1561_ mux_bottom_track_17.INVTX1_2_.out _0404_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_46 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0992_ _0161_ vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__inv_2
XFILLER_12_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1544_ mux_bottom_track_9.INVTX1_2_.out _0387_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1613_ mux_bottom_track_33.INVTX1_2_.out _0456_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_8_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1475_ mux_bottom_track_9.INVTX1_11_.out _0318_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1260_ mux_left_track_17.out vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__clkbuf_1
XFILLER_39_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1191_ clknet_4_11_0_prog_clk mem_left_track_17.DFFR_5_.Q _0113_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_17.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
Xinput8 chanx_left_in[11] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0975_ _0159_ vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__inv_2
XFILLER_59_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1527_ mux_left_track_1.INVTX1_1_.out _0370_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1458_ mux_bottom_track_1.INVTX1_10_.out _0301_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1389_ mux_top_track_24.INVTX1_0_.out _0232_ vssd1 vssd1 vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0760_ mem_top_track_16.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__inv_2
X_0691_ mem_right_track_16.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__inv_2
XFILLER_56_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1312_ net47 vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1174_ clknet_4_1_0_prog_clk mem_left_track_1.DFFR_6_.Q _0096_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_1.DFFR_7_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_13 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0958_ _0158_ vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__inv_2
XFILLER_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0889_ net45 vssd1 vssd1 vccd1 vccd1 mux_left_track_25.INVTX1_8_.out sky130_fd_sc_hd__inv_2
XFILLER_20_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_24 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput164 net164 vssd1 vssd1 vccd1 vccd1 chany_top_out[2] sky130_fd_sc_hd__buf_2
Xoutput153 net153 vssd1 vssd1 vccd1 vccd1 chany_top_out[0] sky130_fd_sc_hd__buf_2
Xoutput131 net131 vssd1 vssd1 vccd1 vccd1 chanx_right_out[7] sky130_fd_sc_hd__buf_2
Xoutput120 net120 vssd1 vssd1 vccd1 vccd1 chanx_right_out[14] sky130_fd_sc_hd__buf_2
Xoutput142 net142 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[17] sky130_fd_sc_hd__buf_2
XFILLER_55_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput66 chany_top_in[12] vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput33 chanx_right_in[17] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_2
Xinput22 chanx_left_in[7] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
Xinput55 chany_bottom_in[2] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
XFILLER_52_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput77 chany_top_in[5] vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput11 chanx_left_in[14] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__dlymetal6s2s_1
X_0743_ mem_top_track_24.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__inv_2
Xinput44 chany_bottom_in[0] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_2
Xinput88 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_ vssd1 vssd1 vccd1
+ vccd1 net88 sky130_fd_sc_hd__clkbuf_1
X_0812_ net88 vssd1 vssd1 vccd1 vccd1 mux_right_track_24.INVTX1_4_.out sky130_fd_sc_hd__inv_2
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0674_ mem_right_track_24.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__inv_2
XFILLER_29_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1157_ clknet_4_8_0_prog_clk mem_bottom_track_1.DFFR_7_.Q _0079_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_9.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
X_1226_ clknet_4_0_0_prog_clk mem_left_track_33.DFFR_2_.Q _0148_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_33.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_52_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1088_ clknet_4_8_0_prog_clk mem_top_track_8.DFFR_4_.Q _0010_ vssd1 vssd1 vccd1 vccd1
+ mem_top_track_8.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1011_ _0163_ vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__inv_2
XFILLER_34_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0726_ mem_right_track_0.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__inv_2
XFILLER_8_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0588_ mem_left_track_9.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__inv_2
X_0657_ mem_bottom_track_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__inv_2
X_1209_ clknet_4_6_0_prog_clk mem_top_track_32.DFFR_1_.Q _0131_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_32.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0511_ mem_bottom_track_33.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__inv_2
X_1560_ mux_left_track_17.INVTX1_2_.out _0403_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1491_ mux_bottom_track_17.INVTX1_11_.out _0334_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1552__186 vssd1 vssd1 vccd1 vccd1 net186 _1552__186/LO sky130_fd_sc_hd__conb_1
X_0709_ mem_right_track_8.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__inv_2
XFILLER_1_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1609__190 vssd1 vssd1 vccd1 vccd1 net190 _1609__190/LO sky130_fd_sc_hd__conb_1
X_0991_ _0161_ vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__inv_2
XFILLER_8_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1474_ mux_bottom_track_9.INVTX1_10_.out _0317_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1612_ mux_bottom_track_33.INVTX1_1_.out _0455_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1543_ mux_bottom_track_9.INVTX1_1_.out _0386_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_5_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1344__173 vssd1 vssd1 vccd1 vccd1 net173 _1344__173/LO sky130_fd_sc_hd__conb_1
XFILLER_14_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput9 chanx_left_in[12] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_2
X_1190_ clknet_4_14_0_prog_clk mem_left_track_17.DFFR_6_.Q _0112_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_17.DFFR_7_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_51_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0974_ _0159_ vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__inv_2
X_1457_ mux_bottom_track_1.INVTX1_9_.out _0300_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1526_ mux_left_track_1.INVTX1_7_.out _0369_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1388_ mux_bottom_track_33.INVTX1_4_.out _0231_ vssd1 vssd1 vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_27_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0690_ mem_right_track_16.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__inv_2
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1311_ net48 vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__clkbuf_1
XFILLER_52_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1173_ clknet_4_14_0_prog_clk mem_bottom_track_17.DFFR_7_.Q _0095_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_25.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_64_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_25 mem_left_track_25.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_14 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput132 net132 vssd1 vssd1 vccd1 vccd1 chanx_right_out[8] sky130_fd_sc_hd__buf_2
X_0888_ net46 vssd1 vssd1 vccd1 vccd1 mux_left_track_25.INVTX1_9_.out sky130_fd_sc_hd__inv_2
X_0957_ _0158_ vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__inv_2
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 chanx_left_out[5] sky130_fd_sc_hd__buf_2
Xoutput121 net121 vssd1 vssd1 vccd1 vccd1 chanx_right_out[15] sky130_fd_sc_hd__buf_2
Xoutput143 net143 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[18] sky130_fd_sc_hd__buf_2
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_0_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_0_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xoutput154 net154 vssd1 vssd1 vccd1 vccd1 chany_top_out[10] sky130_fd_sc_hd__buf_2
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput165 net165 vssd1 vssd1 vccd1 vccd1 chany_top_out[3] sky130_fd_sc_hd__buf_2
X_1509_ mux_bottom_track_25.INVTX1_6_.out _0352_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_46_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput89 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_ vssd1 vssd1 vccd1
+ vccd1 net89 sky130_fd_sc_hd__clkbuf_1
Xinput23 chanx_left_in[8] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__dlymetal6s2s_1
X_0811_ mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1 vccd1
+ vccd1 mux_right_track_24.out sky130_fd_sc_hd__inv_2
X_0673_ mem_right_track_24.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__inv_2
Xinput34 chanx_right_in[18] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_1
Xinput56 chany_bottom_in[3] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__clkbuf_1
X_0742_ mem_top_track_24.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__inv_2
Xinput78 chany_top_in[6] vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__clkbuf_2
Xinput67 chany_top_in[13] vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput12 chanx_left_in[15] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
Xinput45 chany_bottom_in[10] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1156_ clknet_4_14_0_prog_clk mem_bottom_track_9.DFFR_0_.Q _0078_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_9.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_25_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1225_ clknet_4_5_0_prog_clk mem_left_track_33.DFFR_3_.Q _0147_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_33.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1087_ clknet_4_2_0_prog_clk mem_top_track_8.DFFR_5_.Q _0009_ vssd1 vssd1 vccd1 vccd1
+ mem_top_track_8.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1010_ _0152_ vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__buf_4
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0656_ mem_bottom_track_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__inv_2
X_0725_ mem_right_track_0.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__inv_2
XFILLER_57_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0587_ mem_left_track_9.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__inv_2
X_1208_ clknet_4_0_0_prog_clk mem_top_track_32.DFFR_2_.Q _0130_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_32.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_1
X_1585__188 vssd1 vssd1 vccd1 vccd1 net188 _1585__188/LO sky130_fd_sc_hd__conb_1
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1139_ clknet_4_6_0_prog_clk mem_right_track_24.DFFR_1_.Q _0061_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_24.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_4_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1490_ mux_bottom_track_17.INVTX1_10_.out _0333_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0510_ mem_bottom_track_33.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__inv_2
XFILLER_39_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0708_ mem_right_track_8.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__inv_2
X_0639_ mem_bottom_track_9.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__inv_2
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_13_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_13_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1611_ mux_bottom_track_33.INVTX1_5_.out _0454_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
X_0990_ _0161_ vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__inv_2
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1473_ mux_bottom_track_9.INVTX1_9_.out _0316_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1542_ mux_left_track_9.INVTX1_7_.out _0385_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_5_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0973_ _0159_ vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__inv_2
X_1387_ mux_bottom_track_25.INVTX1_8_.out _0230_ vssd1 vssd1 vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1456_ net180 _0299_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
X_1525_ mux_bottom_track_1.INVTX1_5_.out _0368_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_23_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1310_ net49 vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__clkbuf_2
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1172_ clknet_4_13_0_prog_clk mem_bottom_track_25.DFFR_0_.Q _0094_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_25.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
X_0956_ _0158_ vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__inv_2
XFILLER_32_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_15 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 chanx_left_out[6] sky130_fd_sc_hd__buf_2
Xoutput122 net122 vssd1 vssd1 vccd1 vccd1 chanx_right_out[16] sky130_fd_sc_hd__buf_2
X_0887_ net52 vssd1 vssd1 vccd1 vccd1 mux_left_track_25.INVTX1_10_.out sky130_fd_sc_hd__inv_2
Xoutput133 net133 vssd1 vssd1 vccd1 vccd1 chanx_right_out[9] sky130_fd_sc_hd__buf_2
Xoutput155 net155 vssd1 vssd1 vccd1 vccd1 chany_top_out[11] sky130_fd_sc_hd__buf_2
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 chanx_left_out[13] sky130_fd_sc_hd__buf_2
Xoutput166 net166 vssd1 vssd1 vccd1 vccd1 chany_top_out[4] sky130_fd_sc_hd__buf_2
Xoutput144 net144 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[1] sky130_fd_sc_hd__buf_2
X_1439_ mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out _0282_ vssd1
+ vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_2
X_1508_ mux_bottom_track_25.INVTX1_5_.out _0351_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_23_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput13 chanx_left_in[16] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_2
X_0810_ net87 vssd1 vssd1 vccd1 vccd1 mux_right_track_16.INVTX1_4_.out sky130_fd_sc_hd__inv_2
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput35 chanx_right_in[1] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput79 chany_top_in[7] vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__clkbuf_1
Xinput46 chany_bottom_in[11] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_1
X_0672_ mem_right_track_24.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__inv_2
X_0741_ mem_top_track_24.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__inv_2
Xinput24 chanx_left_in[9] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_2
Xinput57 chany_bottom_in[4] vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput68 chany_top_in[14] vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1224_ clknet_4_7_0_prog_clk mem_left_track_33.DFFR_4_.Q _0146_ vssd1 vssd1 vccd1
+ vccd1 net95 sky130_fd_sc_hd__dfrtp_2
XFILLER_52_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1155_ clknet_4_12_0_prog_clk mem_bottom_track_9.DFFR_1_.Q _0077_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_9.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
X_1086_ clknet_4_0_0_prog_clk mem_top_track_8.DFFR_6_.Q _0008_ vssd1 vssd1 vccd1 vccd1
+ mem_top_track_16.DFFR_0_.D sky130_fd_sc_hd__dfrtp_1
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0939_ _0156_ vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__inv_2
XFILLER_20_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0586_ mem_left_track_9.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__inv_2
X_0724_ mem_right_track_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__inv_2
X_0655_ mem_bottom_track_1.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__inv_2
XFILLER_57_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1207_ clknet_4_0_0_prog_clk mem_top_track_32.DFFR_3_.Q _0129_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_32.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_40_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1138_ clknet_4_13_0_prog_clk mem_right_track_24.DFFR_2_.Q _0060_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_24.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
X_1069_ _0168_ vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__inv_2
XFILLER_0_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0707_ mem_right_track_8.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__inv_2
XFILLER_57_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0569_ mem_left_track_17.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__inv_2
X_0638_ mem_bottom_track_9.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__inv_2
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1610_ mux_bottom_track_33.INVTX1_4_.out _0453_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1472_ net181 _0315_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
X_1541_ mux_bottom_track_9.INVTX1_6_.out _0384_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_5_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0972_ _0159_ vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__inv_2
XFILLER_44_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1524_ mux_bottom_track_1.INVTX1_4_.out _0367_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1455_ mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out _0298_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
X_1386_ mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out _0229_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1171_ clknet_4_12_0_prog_clk mem_bottom_track_25.DFFR_1_.Q _0093_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_25.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0886_ mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_25.out sky130_fd_sc_hd__inv_2
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0955_ _0153_ vssd1 vssd1 vccd1 vccd1 _0158_ sky130_fd_sc_hd__buf_4
XFILLER_20_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_16 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput145 net145 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[2] sky130_fd_sc_hd__buf_2
Xoutput156 net156 vssd1 vssd1 vccd1 vccd1 chany_top_out[12] sky130_fd_sc_hd__buf_2
Xoutput123 net123 vssd1 vssd1 vccd1 vccd1 chanx_right_out[17] sky130_fd_sc_hd__buf_2
X_1507_ mux_bottom_track_25.INVTX1_11_.out _0350_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 chanx_left_out[7] sky130_fd_sc_hd__buf_2
Xoutput134 net134 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[0] sky130_fd_sc_hd__buf_2
Xoutput167 net167 vssd1 vssd1 vccd1 vccd1 chany_top_out[5] sky130_fd_sc_hd__buf_2
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 chanx_left_out[14] sky130_fd_sc_hd__buf_2
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1438_ mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out _0281_ vssd1
+ vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_2
X_1369_ mux_bottom_track_1.INVTX1_6_.out _0212_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_62_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0740_ mem_top_track_24.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__inv_2
Xinput25 chanx_right_in[0] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput36 chanx_right_in[2] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_2
Xinput14 chanx_left_in[17] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput47 chany_bottom_in[12] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_2
X_0671_ mem_right_track_24.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__inv_2
Xinput69 chany_top_in[15] vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_1
Xinput58 chany_bottom_in[5] vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1154_ clknet_4_13_0_prog_clk mem_bottom_track_9.DFFR_2_.Q _0076_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_9.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
X_1223_ clknet_4_1_0_prog_clk mem_bottom_track_25.DFFR_7_.Q _0145_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_33.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_37_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1085_ clknet_4_12_0_prog_clk net5 _0007_ vssd1 vssd1 vccd1 vccd1 mem_top_track_0.DFFR_0_.Q
+ sky130_fd_sc_hd__dfrtp_4
X_0869_ net44 vssd1 vssd1 vccd1 vccd1 mux_left_track_1.INVTX1_7_.out sky130_fd_sc_hd__inv_2
X_0938_ _0156_ vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__inv_2
XFILLER_20_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0723_ mem_right_track_0.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__inv_2
X_0585_ mem_left_track_9.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__inv_2
X_0654_ mem_bottom_track_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__inv_2
XFILLER_6_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1137_ clknet_4_15_0_prog_clk mem_right_track_24.DFFR_3_.Q _0059_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_24.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
X_1206_ clknet_4_0_0_prog_clk mem_top_track_32.DFFR_4_.Q _0128_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_0.DFFR_0_.D sky130_fd_sc_hd__dfrtp_1
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1068_ _0168_ vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__inv_2
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0706_ mem_right_track_16.DFFR_0_.D vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__inv_2
XFILLER_30_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0568_ mem_left_track_17.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__inv_2
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0637_ mem_bottom_track_9.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__inv_2
X_0499_ mem_left_track_33.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__inv_2
XFILLER_38_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1540_ mux_bottom_track_9.INVTX1_4_.out _0383_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_8_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1471_ mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out _0314_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_5_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0971_ _0159_ vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__inv_2
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1454_ mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out _0297_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
X_1523_ mux_left_track_1.INVTX1_11_.out _0366_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1385_ mux_bottom_track_25.INVTX1_6_.out _0228_ vssd1 vssd1 vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_27_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1170_ clknet_4_7_0_prog_clk mem_bottom_track_25.DFFR_2_.Q _0092_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_25.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_64_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0885_ net82 vssd1 vssd1 vccd1 vccd1 mux_left_track_17.INVTX1_11_.out sky130_fd_sc_hd__inv_2
XFILLER_20_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0954_ _0157_ vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__inv_2
XFILLER_9_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_17 _0002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 chanx_left_out[8] sky130_fd_sc_hd__buf_2
Xoutput146 net146 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[3] sky130_fd_sc_hd__buf_2
Xoutput124 net124 vssd1 vssd1 vccd1 vccd1 chanx_right_out[18] sky130_fd_sc_hd__buf_2
Xoutput135 net135 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[10] sky130_fd_sc_hd__buf_2
Xoutput157 net157 vssd1 vssd1 vccd1 vccd1 chany_top_out[13] sky130_fd_sc_hd__buf_2
X_1506_ mux_bottom_track_25.INVTX1_10_.out _0349_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1437_ mux_bottom_track_17.INVTX1_0_.out _0280_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 chanx_left_out[15] sky130_fd_sc_hd__buf_2
Xoutput168 net168 vssd1 vssd1 vccd1 vccd1 chany_top_out[6] sky130_fd_sc_hd__buf_2
XFILLER_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1299_ net78 vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__clkbuf_1
X_1368_ mux_bottom_track_17.INVTX1_5_.out _0211_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_23_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput15 chanx_left_in[18] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
Xinput37 chanx_right_in[3] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_1
XFILLER_52_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0670_ mem_right_track_24.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__inv_2
Xinput59 chany_bottom_in[6] vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_2
Xinput48 chany_bottom_in[13] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_2
Xinput26 chanx_right_in[10] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_2
XFILLER_52_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1084_ clknet_4_14_0_prog_clk mem_top_track_0.DFFR_0_.Q _0006_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_0.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
X_1153_ clknet_4_13_0_prog_clk mem_bottom_track_9.DFFR_3_.Q _0075_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_9.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
X_1222_ clknet_4_6_0_prog_clk mem_bottom_track_33.DFFR_0_.Q _0144_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_33.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
X_0868_ net59 vssd1 vssd1 vccd1 vccd1 mux_left_track_1.INVTX1_8_.out sky130_fd_sc_hd__inv_2
X_0799_ mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1 vccd1
+ vccd1 mux_top_track_8.out sky130_fd_sc_hd__inv_2
X_0937_ _0156_ vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__inv_2
XFILLER_57_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0653_ mem_bottom_track_1.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__inv_2
XFILLER_6_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0722_ mem_right_track_0.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__inv_2
X_0584_ mem_left_track_9.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__inv_2
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1205_ clknet_4_15_0_prog_clk mem_left_track_17.DFFR_7_.Q _0127_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_25.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
X_1136_ clknet_4_15_0_prog_clk mem_right_track_24.DFFR_4_.Q _0058_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_24.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
X_1067_ _0168_ vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__inv_2
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0705_ mem_right_track_8.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__inv_2
X_0636_ mem_bottom_track_17.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__inv_2
XFILLER_57_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0567_ mem_left_track_17.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__inv_2
X_0498_ mem_left_track_33.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__inv_2
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1119_ clknet_4_11_0_prog_clk mem_right_track_8.DFFR_5_.Q _0041_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_8.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1470_ mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out _0313_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0619_ mem_bottom_track_25.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__inv_2
X_1599_ mux_left_track_1.INVTX1_10_.out _0442_ vssd1 vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0970_ _0159_ vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__inv_2
X_1453_ mux_bottom_track_25.INVTX1_0_.out _0296_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1522_ mux_left_track_1.INVTX1_10_.out _0365_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1384_ mux_bottom_track_25.INVTX1_5_.out _0227_ vssd1 vssd1 vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_50_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_12_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_12_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_18 _0079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 chanx_left_out[9] sky130_fd_sc_hd__buf_2
Xoutput125 net125 vssd1 vssd1 vccd1 vccd1 chanx_right_out[1] sky130_fd_sc_hd__buf_2
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 chanx_left_out[16] sky130_fd_sc_hd__buf_2
X_0953_ _0157_ vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__inv_2
XFILLER_9_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0884_ net69 vssd1 vssd1 vccd1 vccd1 mux_left_track_17.INVTX1_2_.out sky130_fd_sc_hd__inv_2
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput147 net147 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[4] sky130_fd_sc_hd__buf_2
Xoutput169 net169 vssd1 vssd1 vccd1 vccd1 chany_top_out[7] sky130_fd_sc_hd__buf_2
Xoutput136 net136 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[11] sky130_fd_sc_hd__buf_2
Xoutput158 net158 vssd1 vssd1 vccd1 vccd1 chany_top_out[14] sky130_fd_sc_hd__buf_2
X_1436_ mux_right_track_16.INVTX1_4_.out _0279_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1505_ mux_bottom_track_25.INVTX1_9_.out _0348_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1367_ mux_bottom_track_17.INVTX1_3_.out _0210_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1298_ mux_bottom_track_17.out vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__clkbuf_1
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput27 chanx_right_in[11] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
Xinput49 chany_bottom_in[14] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_2
Xinput16 chanx_left_in[1] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_2
Xinput38 chanx_right_in[4] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1221_ clknet_4_6_0_prog_clk mem_bottom_track_33.DFFR_1_.Q _0143_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_33.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_52_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1152_ clknet_4_15_0_prog_clk mem_bottom_track_9.DFFR_4_.Q _0074_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_9.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
X_1083_ clknet_4_13_0_prog_clk mem_top_track_0.DFFR_1_.Q _0005_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_0.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
X_0936_ _0156_ vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__inv_2
X_0798_ net91 vssd1 vssd1 vccd1 vccd1 mux_top_track_0.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0867_ net48 vssd1 vssd1 vccd1 vccd1 mux_left_track_1.INVTX1_9_.out sky130_fd_sc_hd__inv_2
X_1419_ mux_left_track_9.INVTX1_10_.out _0262_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_28_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0652_ mem_bottom_track_9.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__inv_2
X_0583_ mem_left_track_9.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__inv_2
XFILLER_10_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0721_ mem_right_track_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__inv_2
X_1204_ clknet_4_15_0_prog_clk mem_left_track_25.DFFR_0_.Q _0126_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_25.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1135_ clknet_4_14_0_prog_clk mem_right_track_24.DFFR_5_.Q _0057_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_24.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1066_ _0168_ vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__inv_2
XFILLER_33_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0919_ _0154_ vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__inv_2
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0566_ mem_left_track_17.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__inv_2
X_0635_ mem_bottom_track_17.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__inv_2
X_0704_ mem_right_track_8.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__inv_2
X_0497_ net95 vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__inv_2
X_1049_ _0166_ vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__inv_2
X_1118_ clknet_4_10_0_prog_clk mem_right_track_8.DFFR_6_.Q _0040_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_16.DFFR_0_.D sky130_fd_sc_hd__dfrtp_1
XFILLER_21_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1568__187 vssd1 vssd1 vccd1 vccd1 net187 _1568__187/LO sky130_fd_sc_hd__conb_1
XFILLER_44_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0549_ mem_left_track_25.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__inv_2
X_1598_ mux_left_track_33.INVTX1_6_.out _0441_ vssd1 vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
X_0618_ mem_bottom_track_25.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__inv_2
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1383_ mux_bottom_track_25.INVTX1_4_.out _0226_ vssd1 vssd1 vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1521_ mux_left_track_1.INVTX1_9_.out _0364_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1452_ mux_right_track_24.INVTX1_4_.out _0295_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_35_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0952_ _0157_ vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__inv_2
XANTENNA_19 chany_top_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0883_ net55 vssd1 vssd1 vccd1 vccd1 mux_left_track_17.INVTX1_7_.out sky130_fd_sc_hd__inv_2
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 chanx_left_out[17] sky130_fd_sc_hd__buf_2
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 chanx_right_out[0] sky130_fd_sc_hd__buf_2
Xoutput137 net137 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[12] sky130_fd_sc_hd__buf_2
Xoutput159 net159 vssd1 vssd1 vccd1 vccd1 chany_top_out[15] sky130_fd_sc_hd__buf_2
Xoutput148 net148 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[5] sky130_fd_sc_hd__buf_2
Xoutput126 net126 vssd1 vssd1 vccd1 vccd1 chanx_right_out[2] sky130_fd_sc_hd__buf_2
X_1504_ net183 _0347_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1435_ mux_left_track_17.INVTX1_10_.out _0278_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1366_ mux_left_track_17.INVTX1_10_.out _0209_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1297_ net80 vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__clkbuf_1
XFILLER_23_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput17 chanx_left_in[2] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_2
Xinput39 chanx_right_in[5] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_2
Xinput28 chanx_right_in[12] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1151_ clknet_4_12_0_prog_clk mem_bottom_track_9.DFFR_5_.Q _0073_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_9.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
X_1220_ clknet_4_5_0_prog_clk mem_bottom_track_33.DFFR_2_.Q _0142_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_33.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1082_ clknet_4_15_0_prog_clk mem_top_track_0.DFFR_2_.Q _0004_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_0.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_37_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0866_ net53 vssd1 vssd1 vccd1 vccd1 mux_left_track_1.INVTX1_10_.out sky130_fd_sc_hd__inv_2
X_0935_ _0156_ vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__inv_2
X_0797_ mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1 vccd1
+ vccd1 mux_top_track_0.out sky130_fd_sc_hd__inv_2
X_1349_ mux_left_track_9.INVTX1_9_.out _0192_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1418_ mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out _0261_ vssd1 vssd1
+ vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_43_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0720_ mem_right_track_0.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__inv_2
X_0582_ mem_left_track_9.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__inv_2
X_0651_ mem_bottom_track_9.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__inv_2
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1134_ clknet_4_15_0_prog_clk mem_right_track_24.DFFR_6_.Q _0056_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_24.DFFR_7_.Q sky130_fd_sc_hd__dfrtp_1
X_1203_ clknet_4_15_0_prog_clk mem_left_track_25.DFFR_1_.Q _0125_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_25.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1065_ _0152_ vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__buf_4
XFILLER_18_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0849_ net81 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_0918_ _0154_ vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__inv_2
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0703_ mem_right_track_8.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__inv_2
X_0634_ mem_bottom_track_17.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__inv_2
X_0496_ mem_left_track_33.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__inv_2
X_0565_ mem_left_track_17.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__inv_2
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1117_ clknet_4_3_0_prog_clk mem_right_track_0.DFFR_0_.D _0039_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_0.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1048_ _0166_ vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__inv_2
XFILLER_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0548_ mem_left_track_25.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__inv_2
X_0617_ mem_bottom_track_25.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__inv_2
X_1597_ net189 _0440_ vssd1 vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_41_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1520_ net184 _0363_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
X_1451_ mux_left_track_25.INVTX1_10_.out _0294_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1382_ mux_left_track_25.INVTX1_10_.out _0225_ vssd1 vssd1 vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_50_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0882_ net60 vssd1 vssd1 vccd1 vccd1 mux_left_track_17.INVTX1_8_.out sky130_fd_sc_hd__inv_2
XFILLER_40_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0951_ _0157_ vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__inv_2
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput138 net138 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[13] sky130_fd_sc_hd__buf_2
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1503_ mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out _0346_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
Xoutput127 net127 vssd1 vssd1 vccd1 vccd1 chanx_right_out[3] sky130_fd_sc_hd__buf_2
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 chanx_right_out[10] sky130_fd_sc_hd__buf_2
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 chanx_left_out[18] sky130_fd_sc_hd__buf_2
Xoutput149 net149 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[6] sky130_fd_sc_hd__buf_2
X_1296_ net81 vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__clkbuf_1
XFILLER_55_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1365_ mux_left_track_17.INVTX1_9_.out _0208_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1434_ mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out _0277_ vssd1
+ vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 chanx_left_in[3] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput29 chanx_right_in[13] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1150_ clknet_4_13_0_prog_clk mem_bottom_track_9.DFFR_6_.Q _0072_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_17.DFFR_0_.D sky130_fd_sc_hd__dfrtp_1
XFILLER_45_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1081_ clknet_4_10_0_prog_clk mem_top_track_0.DFFR_3_.Q _0003_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_0.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
X_0865_ mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_1.out sky130_fd_sc_hd__inv_2
X_0934_ _0156_ vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__inv_2
XFILLER_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1417_ mux_bottom_track_9.INVTX1_2_.out _0260_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_0796_ mem_top_track_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__inv_2
X_1279_ mux_right_track_16.out vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__clkbuf_1
X_1348_ mux_left_track_9.INVTX1_7_.out _0191_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_11_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0581_ mem_left_track_9.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__inv_2
X_0650_ mem_bottom_track_9.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__inv_2
X_1202_ clknet_4_15_0_prog_clk mem_left_track_25.DFFR_2_.Q _0124_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_25.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
X_1133_ clknet_4_10_0_prog_clk mem_right_track_16.DFFR_0_.D _0055_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_16.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
X_1064_ _0167_ vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__inv_2
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0779_ mem_top_track_8.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__inv_2
X_0917_ _0154_ vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__inv_2
X_0848_ net70 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.INVTX1_2_.out sky130_fd_sc_hd__inv_2
XFILLER_0_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0633_ mem_bottom_track_17.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__inv_2
X_0702_ mem_right_track_8.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__inv_2
X_0564_ mem_left_track_17.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__inv_2
X_0495_ mem_left_track_33.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__inv_2
X_1047_ _0166_ vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__inv_2
XFILLER_38_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_9_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_9_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1116_ clknet_4_3_0_prog_clk mem_right_track_0.DFFR_0_.Q _0038_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_0.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1360__174 vssd1 vssd1 vccd1 vccd1 net174 _1360__174/LO sky130_fd_sc_hd__conb_1
XFILLER_8_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1596_ mux_bottom_track_33.INVTX1_7_.out _0439_ vssd1 vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0616_ mem_bottom_track_25.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__inv_2
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0547_ mem_left_track_25.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__inv_2
XFILLER_38_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1450_ mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out _0293_ vssd1
+ vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_2
X_1381_ mux_left_track_25.INVTX1_8_.out _0224_ vssd1 vssd1 vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1408__177 vssd1 vssd1 vccd1 vccd1 net177 _1408__177/LO sky130_fd_sc_hd__conb_1
XFILLER_50_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1579_ mux_left_track_25.INVTX1_8_.out _0422_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0881_ net62 vssd1 vssd1 vccd1 vccd1 mux_left_track_17.INVTX1_9_.out sky130_fd_sc_hd__inv_2
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0950_ _0157_ vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__inv_2
XFILLER_13_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 chanx_right_out[11] sky130_fd_sc_hd__buf_2
Xoutput128 net128 vssd1 vssd1 vccd1 vccd1 chanx_right_out[4] sky130_fd_sc_hd__buf_2
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1433_ mux_bottom_track_17.INVTX1_2_.out _0276_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
Xoutput139 net139 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[14] sky130_fd_sc_hd__buf_2
X_1502_ mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out _0345_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 chanx_left_out[1] sky130_fd_sc_hd__buf_2
XFILLER_55_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1295_ net64 vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__clkbuf_1
X_1364_ mux_left_track_17.INVTX1_7_.out _0207_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_63_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput19 chanx_left_in[4] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_11_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_11_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1080_ clknet_4_2_0_prog_clk mem_top_track_0.DFFR_4_.Q _0002_ vssd1 vssd1 vccd1 vccd1
+ mem_top_track_0.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0864_ net15 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.INVTX1_11_.out sky130_fd_sc_hd__inv_2
X_0795_ mem_top_track_0.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__inv_2
X_0933_ _0153_ vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__buf_4
XFILLER_9_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1347_ mux_bottom_track_25.INVTX1_11_.out _0190_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1416_ mux_bottom_track_9.INVTX1_1_.out _0259_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1278_ net23 vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__clkbuf_2
XFILLER_36_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1201_ clknet_4_14_0_prog_clk mem_left_track_25.DFFR_3_.Q _0123_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_25.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
X_0580_ mem_left_track_9.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__inv_2
XFILLER_6_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1132_ clknet_4_10_0_prog_clk mem_right_track_16.DFFR_0_.Q _0054_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_16.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_2
X_1063_ _0167_ vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__inv_2
X_0916_ _0154_ vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__inv_2
XFILLER_33_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0847_ net36 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.INVTX1_3_.out sky130_fd_sc_hd__inv_2
X_0778_ mem_top_track_8.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__inv_2
XFILLER_56_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0632_ mem_bottom_track_17.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__inv_2
X_0701_ mem_right_track_8.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__inv_2
X_0563_ mem_left_track_17.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__inv_2
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0494_ mem_left_track_33.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__inv_2
XFILLER_2_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1046_ _0166_ vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__inv_2
XFILLER_21_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1115_ clknet_4_5_0_prog_clk mem_right_track_0.DFFR_1_.Q _0037_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_0.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0546_ mem_left_track_25.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__inv_2
X_0615_ mem_bottom_track_25.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__inv_2
X_1595_ mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out _0438_ vssd1
+ vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_7_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1029_ _0164_ vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__inv_2
XFILLER_39_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1380_ mux_left_track_25.INVTX1_7_.out _0223_ vssd1 vssd1 vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_4_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1578_ mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out _0421_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0529_ mem_top_track_32.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__inv_2
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0880_ net51 vssd1 vssd1 vccd1 vccd1 mux_left_track_17.INVTX1_10_.out sky130_fd_sc_hd__inv_2
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 chanx_left_out[2] sky130_fd_sc_hd__buf_2
XFILLER_13_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput129 net129 vssd1 vssd1 vccd1 vccd1 chanx_right_out[5] sky130_fd_sc_hd__buf_2
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 chanx_right_out[12] sky130_fd_sc_hd__buf_2
X_1363_ mux_bottom_track_17.INVTX1_11_.out _0206_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1501_ mux_bottom_track_17.INVTX1_0_.out _0344_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1432_ mux_bottom_track_17.INVTX1_1_.out _0275_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1294_ mux_bottom_track_25.out vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__clkbuf_1
XFILLER_23_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0932_ _0155_ vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__inv_2
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0863_ net76 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0794_ mem_top_track_0.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__inv_2
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1346_ mux_bottom_track_9.INVTX1_11_.out _0189_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_28_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1415_ mux_left_track_1.INVTX1_1_.out _0258_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_36_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1277_ net24 vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__clkbuf_2
XFILLER_22_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1200_ clknet_4_14_0_prog_clk mem_left_track_25.DFFR_4_.Q _0122_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_25.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1131_ clknet_4_10_0_prog_clk mem_right_track_16.DFFR_1_.Q _0053_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_16.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_2
X_1062_ _0167_ vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__inv_2
XFILLER_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0915_ _0154_ vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__inv_2
X_0846_ net41 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.INVTX1_4_.out sky130_fd_sc_hd__inv_2
X_0777_ mem_top_track_8.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__inv_2
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1329_ mux_bottom_track_33.INVTX1_5_.out _0172_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_17_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0700_ mem_right_track_16.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__inv_2
XFILLER_30_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0562_ mem_left_track_17.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__inv_2
X_0631_ mem_bottom_track_17.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__inv_2
XFILLER_53_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0493_ mem_left_track_33.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__inv_2
X_1114_ clknet_4_4_0_prog_clk mem_right_track_0.DFFR_2_.Q _0036_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_0.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1045_ _0166_ vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__inv_2
X_0829_ net16 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.INVTX1_8_.out sky130_fd_sc_hd__inv_2
XFILLER_21_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0545_ mem_left_track_25.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__inv_2
X_0614_ mem_bottom_track_25.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__inv_2
X_1594_ mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out _0437_ vssd1
+ vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1028_ _0164_ vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__inv_2
XFILLER_14_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1577_ mux_bottom_track_25.INVTX1_2_.out _0420_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0528_ mem_right_track_32.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__inv_2
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 chanx_left_out[3] sky130_fd_sc_hd__buf_2
X_1500_ mux_bottom_track_17.INVTX1_4_.out _0343_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_40_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 chanx_right_out[13] sky130_fd_sc_hd__buf_2
X_1293_ net66 vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__clkbuf_1
X_1431_ mux_left_track_33.INVTX1_1_.out _0274_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1362_ mux_bottom_track_17.INVTX1_10_.out _0205_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_48_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1629_ mux_bottom_track_33.INVTX1_0_.out _0472_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0862_ net64 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_0931_ _0155_ vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__inv_2
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0793_ mem_top_track_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__inv_2
X_1345_ mux_bottom_track_9.INVTX1_9_.out _0188_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1414_ mux_left_track_25.INVTX1_9_.out _0257_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1276_ net7 vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__clkbuf_1
XFILLER_28_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1130_ clknet_4_11_0_prog_clk mem_right_track_16.DFFR_2_.Q _0052_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_16.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_33_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1061_ _0167_ vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__inv_2
XFILLER_18_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0845_ net43 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.INVTX1_5_.out sky130_fd_sc_hd__inv_2
X_0914_ _0154_ vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__inv_2
X_0776_ mem_top_track_8.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__inv_2
X_1259_ net42 vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__clkbuf_1
XFILLER_56_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1328_ net172 _0171_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_64_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0561_ mem_left_track_17.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__inv_2
X_0630_ mem_bottom_track_17.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__inv_2
XFILLER_53_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1044_ _0166_ vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__inv_2
XFILLER_38_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1113_ clknet_4_5_0_prog_clk mem_right_track_0.DFFR_3_.Q _0035_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_0.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0759_ mem_top_track_16.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__inv_2
X_0828_ net23 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.INVTX1_9_.out sky130_fd_sc_hd__inv_2
XFILLER_29_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0613_ mem_bottom_track_25.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__inv_2
XFILLER_7_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0544_ mem_left_track_25.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__inv_2
X_1593_ mux_bottom_track_25.INVTX1_3_.out _0436_ vssd1 vssd1 vccd1 vccd1 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1027_ _0164_ vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__inv_2
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_8_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_8_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1576_ mux_left_track_25.INVTX1_2_.out _0419_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0527_ mem_right_track_32.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0442_ sky130_fd_sc_hd__inv_2
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 chanx_left_out[4] sky130_fd_sc_hd__buf_2
X_1430_ mux_left_track_17.INVTX1_9_.out _0273_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1361_ mux_bottom_track_17.INVTX1_9_.out _0204_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_36_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1292_ net67 vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__clkbuf_1
XFILLER_63_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1559_ mux_bottom_track_17.INVTX1_1_.out _0402_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1628_ mux_bottom_track_33.INVTX1_2_.out _0471_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0861_ net71 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.INVTX1_2_.out sky130_fd_sc_hd__inv_2
X_0930_ _0155_ vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__inv_2
X_0792_ mem_top_track_0.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__inv_2
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1413_ mux_left_track_9.INVTX1_9_.out _0256_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1275_ mux_right_track_24.out vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1344_ net173 _0187_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1060_ _0167_ vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__inv_2
XFILLER_2_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0775_ mem_top_track_8.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__inv_2
X_0844_ net32 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.INVTX1_6_.out sky130_fd_sc_hd__inv_2
X_0913_ _0154_ vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__inv_2
XFILLER_56_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1327_ mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out _0170_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
X_1258_ net43 vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__clkbuf_1
X_1189_ clknet_4_2_0_prog_clk mem_left_track_1.DFFR_7_.Q _0111_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_9.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_4_10_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_10_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_24_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0560_ mem_left_track_17.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__inv_2
XFILLER_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1112_ clknet_4_1_0_prog_clk mem_right_track_0.DFFR_4_.Q _0034_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_0.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
X_1043_ _0152_ vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__buf_4
XFILLER_61_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0758_ mem_top_track_16.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__inv_2
X_0827_ net8 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.INVTX1_10_.out sky130_fd_sc_hd__inv_2
X_0689_ mem_right_track_16.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__inv_2
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0612_ mem_bottom_track_25.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__inv_2
XFILLER_7_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1592_ mux_left_track_33.INVTX1_5_.out _0435_ vssd1 vssd1 vccd1 vccd1 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0543_ mem_left_track_25.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__inv_2
XFILLER_53_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1026_ _0164_ vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__inv_2
XFILLER_61_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1575_ mux_bottom_track_25.INVTX1_1_.out _0418_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0526_ mem_right_track_32.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__inv_2
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1009_ _0162_ vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__inv_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1360_ net174 _0203_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_2
X_1291_ net68 vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__clkbuf_1
XFILLER_63_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1489_ mux_bottom_track_17.INVTX1_9_.out _0332_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1627_ mux_left_track_33.INVTX1_6_.out _0470_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0509_ mem_bottom_track_33.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__inv_2
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1558_ mux_left_track_17.INVTX1_7_.out _0401_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_54_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0860_ net37 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.INVTX1_3_.out sky130_fd_sc_hd__inv_2
XFILLER_42_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0791_ mem_top_track_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__inv_2
XFILLER_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1412_ mux_left_track_9.INVTX1_7_.out _0255_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1343_ mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out _0186_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_3_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1274_ net9 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__clkbuf_1
XFILLER_24_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0989_ _0161_ vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__inv_2
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0912_ _0154_ vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__inv_2
X_0843_ net1 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.INVTX1_7_.out sky130_fd_sc_hd__inv_2
X_0774_ mem_top_track_8.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__inv_2
XFILLER_5_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1326_ mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out _0169_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_64_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1188_ clknet_4_9_0_prog_clk mem_left_track_9.DFFR_0_.Q _0110_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_9.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
X_1257_ net26 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1042_ _0165_ vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__inv_2
X_1111_ clknet_4_4_0_prog_clk mem_right_track_0.DFFR_5_.Q _0033_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_0.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_61_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0826_ mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1 vccd1
+ vccd1 mux_bottom_track_9.out sky130_fd_sc_hd__inv_2
X_0688_ mem_right_track_16.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__inv_2
X_0757_ mem_top_track_16.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__inv_2
XFILLER_29_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1309_ mux_top_track_32.out vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__clkbuf_1
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1376__175 vssd1 vssd1 vccd1 vccd1 net175 _1376__175/LO sky130_fd_sc_hd__conb_1
X_0542_ mem_left_track_25.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__inv_2
X_1591_ mux_bottom_track_1.INVTX1_10_.out _0434_ vssd1 vssd1 vccd1 vccd1 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
X_0611_ mem_bottom_track_25.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__inv_2
XFILLER_7_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1025_ _0164_ vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__inv_2
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0809_ mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1 vccd1
+ vccd1 mux_right_track_16.out sky130_fd_sc_hd__inv_2
XFILLER_55_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_1 _0010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1574_ mux_left_track_25.INVTX1_7_.out _0417_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0525_ mem_right_track_32.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__inv_2
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1008_ _0162_ vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__inv_2
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1290_ mux_bottom_track_33.out vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__clkbuf_1
XFILLER_63_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1626_ mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out _0469_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
X_1488_ net182 _0331_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
X_1557_ mux_bottom_track_17.INVTX1_6_.out _0400_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
X_0508_ mem_bottom_track_33.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__inv_2
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0790_ mem_top_track_0.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__inv_2
XFILLER_5_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1411_ mux_bottom_track_9.INVTX1_11_.out _0254_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1342_ mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out _0185_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_3_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1273_ net10 vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0988_ _0153_ vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__buf_4
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1609_ net190 _0452_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_59_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0842_ net17 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.INVTX1_8_.out sky130_fd_sc_hd__inv_2
XFILLER_33_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0911_ _0153_ vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__buf_4
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0773_ mem_top_track_8.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__inv_2
X_1256_ mux_left_track_25.out vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1325_ mux_top_track_0.out vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__clkbuf_1
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1187_ clknet_4_13_0_prog_clk mem_left_track_9.DFFR_1_.Q _0109_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_9.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_24_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1110_ clknet_4_4_0_prog_clk mem_right_track_0.DFFR_6_.Q _0032_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_0.DFFR_7_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1041_ _0165_ vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__inv_2
X_0825_ net10 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.INVTX1_11_.out sky130_fd_sc_hd__inv_2
XFILLER_14_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0756_ mem_top_track_16.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__inv_2
X_0687_ mem_right_track_16.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__inv_2
X_1308_ net51 vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__clkbuf_2
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0541_ mem_left_track_25.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__inv_2
X_0610_ mem_bottom_track_25.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__inv_2
X_1590_ mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out _0433_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_4
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1024_ _0164_ vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__inv_2
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0808_ net90 vssd1 vssd1 vccd1 vccd1 mux_right_track_8.INVTX1_4_.out sky130_fd_sc_hd__inv_2
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0739_ mem_top_track_24.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__inv_2
XFILLER_37_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_2 _0064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1573_ mux_bottom_track_25.INVTX1_6_.out _0416_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0524_ mem_right_track_32.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__inv_2
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1007_ _0162_ vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__inv_2
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1556_ mux_bottom_track_17.INVTX1_5_.out _0399_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1625_ mux_bottom_track_33.INVTX1_1_.out _0468_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1487_ mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out _0330_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_39_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0507_ mem_bottom_track_33.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__inv_2
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_7_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_7_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1410_ mux_bottom_track_9.INVTX1_9_.out _0253_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1341_ mux_top_track_0.INVTX1_0_.out _0184_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1272_ net11 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0987_ _0160_ vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__inv_2
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1608_ mux_bottom_track_33.INVTX1_7_.out _0451_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1539_ mux_left_track_9.INVTX1_11_.out _0382_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0772_ mem_top_track_8.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__inv_2
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0841_ net24 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.INVTX1_9_.out sky130_fd_sc_hd__inv_2
X_0910_ _0152_ vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__clkbuf_4
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1255_ net28 vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__clkbuf_1
X_1324_ net44 vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__clkbuf_2
X_1186_ clknet_4_7_0_prog_clk mem_left_track_9.DFFR_2_.Q _0108_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_9.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_32_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1040_ _0165_ vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__inv_2
XFILLER_64_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0824_ net63 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0755_ mem_top_track_16.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__inv_2
XFILLER_9_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0686_ mem_right_track_16.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__inv_2
XFILLER_29_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1307_ net52 vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__clkbuf_2
XFILLER_37_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1169_ clknet_4_2_0_prog_clk mem_bottom_track_25.DFFR_3_.Q _0091_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_25.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0540_ mem_top_track_32.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__inv_2
XFILLER_53_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1023_ _0164_ vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__inv_2
X_1424__178 vssd1 vssd1 vccd1 vccd1 net178 _1424__178/LO sky130_fd_sc_hd__conb_1
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0807_ mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1 vccd1
+ vccd1 mux_right_track_8.out sky130_fd_sc_hd__inv_2
X_0738_ mem_top_track_24.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__inv_2
X_0669_ mem_right_track_24.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__inv_2
XFILLER_39_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1572_ mux_bottom_track_25.INVTX1_5_.out _0415_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
XANTENNA_3 _0119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1597__189 vssd1 vssd1 vccd1 vccd1 net189 _1597__189/LO sky130_fd_sc_hd__conb_1
XFILLER_6_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0523_ mem_right_track_32.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__inv_2
XFILLER_54_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1006_ _0162_ vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__inv_2
XFILLER_19_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 ccff_tail sky130_fd_sc_hd__buf_2
XFILLER_48_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1624_ mux_left_track_33.INVTX1_1_.out _0467_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1555_ mux_left_track_17.INVTX1_11_.out _0398_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_0506_ mem_bottom_track_33.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__inv_2
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1486_ mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out _0329_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_39_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1340_ mux_bottom_track_1.INVTX1_5_.out _0183_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1271_ mux_right_track_32.out vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__clkbuf_1
X_0986_ _0160_ vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__inv_2
XFILLER_59_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1538_ mux_left_track_9.INVTX1_10_.out _0381_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1469_ mux_bottom_track_1.INVTX1_0_.out _0312_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1607_ mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out _0450_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_63_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0771_ mem_top_track_8.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__inv_2
X_0840_ net12 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.INVTX1_10_.out sky130_fd_sc_hd__inv_2
X_1323_ net54 vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__clkbuf_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1254_ net29 vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__clkbuf_1
X_1185_ clknet_4_4_0_prog_clk mem_left_track_9.DFFR_3_.Q _0107_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_9.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_24_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0969_ _0159_ vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__inv_2
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0685_ mem_right_track_16.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__inv_2
X_0754_ mem_top_track_16.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__inv_2
X_0823_ net78 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_1306_ mux_bottom_track_1.out vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1168_ clknet_4_1_0_prog_clk mem_bottom_track_25.DFFR_4_.Q _0090_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_25.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
X_1099_ clknet_4_0_0_prog_clk mem_top_track_16.DFFR_1_.Q _0021_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_16.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_47_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1456__180 vssd1 vssd1 vccd1 vccd1 net180 _1456__180/LO sky130_fd_sc_hd__conb_1
XFILLER_61_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1022_ _0164_ vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__inv_2
X_0806_ net89 vssd1 vssd1 vccd1 vccd1 mux_right_track_0.INVTX1_4_.out sky130_fd_sc_hd__inv_2
X_0737_ mem_top_track_24.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__inv_2
X_0668_ mem_bottom_track_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__inv_2
XFILLER_55_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0599_ mem_left_track_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__inv_2
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1571_ mux_left_track_25.INVTX1_11_.out _0414_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0522_ mem_right_track_32.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__inv_2
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_4 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1005_ _0162_ vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__inv_2
XFILLER_41_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1621__191 vssd1 vssd1 vccd1 vccd1 net191 _1621__191/LO sky130_fd_sc_hd__conb_1
XFILLER_40_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 chanx_left_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1554_ mux_left_track_17.INVTX1_10_.out _0397_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1485_ mux_bottom_track_9.INVTX1_0_.out _0328_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1623_ mux_left_track_33.INVTX1_5_.out _0466_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
X_0505_ mem_bottom_track_33.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__inv_2
.ends

