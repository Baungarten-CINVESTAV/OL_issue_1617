* NGSPICE file created from sb_1__4_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_4 abstract view
.subckt sky130_fd_sc_hd__ebufn_4 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

.subckt sb_1__4_ bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_ bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
+ bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_ bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
+ ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11] chanx_left_in[12]
+ chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16] chanx_left_in[17]
+ chanx_left_in[18] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4]
+ chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_in[9]
+ chanx_left_out[0] chanx_left_out[10] chanx_left_out[11] chanx_left_out[12] chanx_left_out[13]
+ chanx_left_out[14] chanx_left_out[15] chanx_left_out[16] chanx_left_out[17] chanx_left_out[18]
+ chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chanx_right_in[0]
+ chanx_right_in[10] chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14]
+ chanx_right_in[15] chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10]
+ chanx_right_out[11] chanx_right_out[12] chanx_right_out[13] chanx_right_out[14]
+ chanx_right_out[15] chanx_right_out[16] chanx_right_out[17] chanx_right_out[18]
+ chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4] chanx_right_out[5]
+ chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chanx_right_out[9] chany_bottom_in[0]
+ chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13]
+ chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17]
+ chany_bottom_in[18] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4]
+ chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_in[9]
+ chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11] chany_bottom_out[12]
+ chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15] chany_bottom_out[16]
+ chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[1] chany_bottom_out[2]
+ chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6]
+ chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
+ left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_ left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_ left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_ left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_
+ left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_ left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_
+ left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_ pReset prog_clk right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_ right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_ right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_ right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_
+ right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_ right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_
+ right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_ vccd1 vssd1 vssd1_uq0
+ vccd1_uq0
XFILLER_54_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1119__148 vssd1 vssd1 vccd1 vccd1 net148 _1119__148/LO sky130_fd_sc_hd__conb_1
XFILLER_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0419_ mem_bottom_track_25.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0770_ _0122_ vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__inv_2
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1184_ net158 _0298_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_20_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0899_ clknet_4_1_0_prog_clk mem_right_track_32.DFFR_4_.Q _0012_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_1.DFFR_0_.D sky130_fd_sc_hd__dfrtp_1
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0822_ _0127_ vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__inv_2
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0684_ net9 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_19.INVTX1_2_.out sky130_fd_sc_hd__inv_2
X_0753_ _0120_ vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__inv_2
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1236_ mux_left_track_33.INVTX1_4_.out _0350_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_64_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1167_ mux_bottom_track_5.INVTX1_0_.out _0281_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_5.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1098_ mux_left_track_9.INVTX1_7_.out _0212_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1021_ mux_right_track_8.out vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__clkbuf_1
XFILLER_34_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0805_ _0125_ vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__inv_2
X_0667_ net21 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_11.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_0598_ mem_right_track_0.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__inv_2
X_0736_ _0158_ vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__inv_2
XFILLER_44_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1219_ mux_bottom_track_27.INVTX1_0_.out _0333_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0521_ mem_right_track_32.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__inv_2
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0452_ mem_bottom_track_21.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__clkbuf_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0383_ mem_right_track_0.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__inv_2
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1209__163 vssd1 vssd1 vccd1 vccd1 net163 _1209__163/LO sky130_fd_sc_hd__conb_1
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1004_ net35 vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__clkbuf_1
XFILLER_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0719_ _0156_ vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__inv_2
XFILLER_1_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 chanx_left_out[3] sky130_fd_sc_hd__buf_2
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 chanx_left_out[10] sky130_fd_sc_hd__buf_2
XFILLER_63_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0435_ mem_bottom_track_19.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__inv_2
X_0504_ mem_bottom_track_7.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__inv_2
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0418_ mem_bottom_track_25.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__inv_2
XFILLER_27_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_6_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_6_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_49_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1183_ mux_bottom_track_15.INVTX1_0_.out _0297_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_17_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0898_ clknet_4_6_0_prog_clk mem_left_track_17.DFFR_7_.Q _0011_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_25.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0821_ net73 vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__buf_4
X_0752_ _0120_ vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__inv_2
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0683_ net28 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_19.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_49_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1166_ mux_bottom_track_5.mux_2level_tapbuf_basis_input3_mem3_0_out _0280_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_5.mux_2level_tapbuf_basis_input3_mem3_1_out sky130_fd_sc_hd__ebufn_2
X_1235_ net166 _0349_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_52_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1097_ mux_left_track_9.INVTX1_6_.out _0211_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_20_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1020_ net19 vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__clkbuf_1
XFILLER_38_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0804_ _0125_ vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__inv_2
X_0735_ _0158_ vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__inv_2
XFILLER_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0666_ net40 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_11.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_29_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0597_ mem_right_track_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__inv_2
X_1149_ mux_bottom_track_7.INVTX1_2_.out _0263_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_7.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1218_ mux_bottom_track_27.INVTX1_2_.out _0332_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_52_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0520_ mem_right_track_32.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__inv_2
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0451_ mem_bottom_track_21.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__inv_2
X_1003_ net36 vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__clkbuf_1
XFILLER_34_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0718_ _0156_ vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__inv_2
X_0649_ mux_bottom_track_7.mux_2level_tapbuf_basis_input3_mem3_1_out vssd1 vssd1 vccd1
+ vccd1 mux_bottom_track_7.out sky130_fd_sc_hd__inv_2
XFILLER_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 chanx_left_out[4] sky130_fd_sc_hd__buf_2
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 chanx_left_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0434_ _0137_ vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__clkbuf_1
X_0503_ mem_bottom_track_7.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__inv_2
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0417_ mem_bottom_track_25.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__inv_2
XFILLER_10_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1188__159 vssd1 vssd1 vccd1 vccd1 net159 _1188__159/LO sky130_fd_sc_hd__conb_1
XFILLER_18_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1182_ mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_0_out _0296_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_64_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0897_ clknet_4_12_0_prog_clk mem_left_track_25.DFFR_0_.Q _0010_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_25.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_2
XFILLER_59_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0751_ _0120_ vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__inv_2
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0820_ _0126_ vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__inv_2
X_0682_ mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_2_out vssd1 vssd1
+ vccd1 vccd1 mux_bottom_track_19.out sky130_fd_sc_hd__inv_2
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1165_ mux_bottom_track_5.INVTX1_3_.out _0279_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_5.mux_2level_tapbuf_basis_input2_mem2_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1234_ mux_left_track_33.INVTX1_7_.out _0348_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1096_ mux_left_track_9.INVTX1_5_.out _0210_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_52_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0949_ clknet_4_15_0_prog_clk mem_bottom_track_27.DFFR_0_.Q _0062_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_27.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0665_ mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_1_out vssd1 vssd1
+ vccd1 vccd1 mux_bottom_track_11.out sky130_fd_sc_hd__inv_2
X_0803_ _0125_ vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__inv_2
X_0734_ _0158_ vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__inv_2
X_0596_ mem_right_track_8.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__inv_2
XFILLER_52_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1079_ mux_left_track_17.INVTX1_5_.out _0193_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1148_ mux_bottom_track_25.INVTX1_1_.out _0262_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_7.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1217_ mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_0_out _0331_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_20_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0450_ mem_bottom_track_21.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__inv_2
X_1002_ mux_left_track_9.out vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__clkbuf_1
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0648_ net22 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.INVTX1_3_.out sky130_fd_sc_hd__inv_2
X_0717_ _0156_ vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__inv_2
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0579_ mem_right_track_16.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__inv_2
XFILLER_25_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 chanx_left_out[12] sky130_fd_sc_hd__buf_2
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 chanx_left_out[5] sky130_fd_sc_hd__buf_2
XFILLER_0_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0502_ mem_bottom_track_7.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__inv_2
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0433_ mem_bottom_track_23.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__clkbuf_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1197__161 vssd1 vssd1 vccd1 vccd1 net161 _1197__161/LO sky130_fd_sc_hd__conb_1
XFILLER_3_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0416_ _0131_ vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1181_ mux_bottom_track_15.INVTX1_1_.out _0295_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0896_ clknet_4_12_0_prog_clk mem_left_track_25.DFFR_1_.Q _0009_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_25.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0750_ _0120_ vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__inv_2
X_0681_ net18 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_37.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XFILLER_56_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1233_ mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out _0347_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1164_ mux_bottom_track_25.INVTX1_1_.out _0278_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_5.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1095_ net146 _0209_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_0948_ clknet_4_13_0_prog_clk mem_bottom_track_23.DFFR_1_.Q _0061_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_25.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_2
X_0879_ clknet_4_9_0_prog_clk mem_left_track_9.DFFR_2_.Q _0112_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_9.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0802_ _0125_ vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__inv_2
X_0733_ _0155_ vssd1 vssd1 vccd1 vccd1 _0158_ sky130_fd_sc_hd__buf_4
XFILLER_6_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0664_ net20 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_1216_ mux_bottom_track_27.INVTX1_1_.out _0330_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_2
X_0595_ mem_right_track_8.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__inv_2
XFILLER_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1147_ net151 _0261_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_7.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1078_ mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out _0192_ vssd1
+ vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out sky130_fd_sc_hd__ebufn_4
XFILLER_4_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1001_ net38 vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__clkbuf_2
XFILLER_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0647_ net25 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0716_ _0156_ vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__inv_2
X_0578_ mem_right_track_16.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__inv_2
XFILLER_57_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 chanx_left_out[13] sky130_fd_sc_hd__buf_2
XFILLER_56_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0432_ mem_bottom_track_23.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__inv_2
X_0501_ mem_bottom_track_3.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__inv_2
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1141__150 vssd1 vssd1 vccd1 vccd1 net150 _1141__150/LO sky130_fd_sc_hd__conb_1
X_0415_ mem_bottom_track_27.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1180_ net157 _0294_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_32_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0895_ clknet_4_11_0_prog_clk mem_left_track_25.DFFR_2_.Q _0008_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_25.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_2
XFILLER_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0680_ mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_1_out vssd1 vssd1
+ vccd1 vccd1 mux_bottom_track_37.out sky130_fd_sc_hd__inv_2
X_1232_ mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out _0346_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_64_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1163_ mux_bottom_track_23.INVTX1_1_.out _0277_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_5.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1094_ mux_left_track_9.INVTX1_8_.out _0208_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_0947_ clknet_4_15_0_prog_clk mem_bottom_track_25.DFFR_0_.Q _0060_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_25.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0878_ clknet_4_2_0_prog_clk mem_left_track_9.DFFR_3_.Q _0111_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_9.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_55_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_5_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_5_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0801_ _0125_ vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__inv_2
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0594_ mem_right_track_8.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__inv_2
X_0663_ net39 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0732_ _0157_ vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__inv_2
XFILLER_10_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1215_ net164 _0329_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_1_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1146_ mux_bottom_track_7.INVTX1_3_.out _0260_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_7.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_52_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1077_ mux_left_track_17.INVTX1_4_.out _0191_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_45_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1000_ net39 vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__clkbuf_1
XFILLER_13_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0715_ _0156_ vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__inv_2
XFILLER_57_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0646_ net3 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_0577_ mem_right_track_16.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__inv_2
XFILLER_57_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1129_ net149 _0243_ vssd1 vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input2_mem2_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0431_ _0136_ vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__clkbuf_1
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0500_ mem_bottom_track_3.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__inv_2
XFILLER_47_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0629_ net51 vssd1 vssd1 vccd1 vccd1 mux_left_track_17.INVTX1_6_.out sky130_fd_sc_hd__inv_2
XFILLER_26_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0414_ mem_bottom_track_27.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__inv_2
XFILLER_50_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0894_ clknet_4_6_0_prog_clk mem_left_track_25.DFFR_3_.Q _0007_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_25.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_4_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1162_ net153 _0276_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_5.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1231_ mux_bottom_track_1.INVTX1_0_.out _0345_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_64_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1093_ mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out _0207_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out sky130_fd_sc_hd__ebufn_4
XFILLER_20_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0877_ clknet_4_8_0_prog_clk mem_left_track_9.DFFR_4_.Q _0110_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_9.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
X_0946_ clknet_4_3_0_prog_clk mem_bottom_track_21.DFFR_1_.Q _0059_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_23.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0731_ _0157_ vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__inv_2
X_0800_ _0125_ vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__inv_2
X_0662_ mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_1_out vssd1 vssd1 vccd1
+ vccd1 mux_bottom_track_9.out sky130_fd_sc_hd__inv_2
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0593_ mem_right_track_8.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__inv_2
XFILLER_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1145_ mux_bottom_track_1.INVTX1_0_.out _0259_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_25_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1214_ mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_1_out _0328_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1076_ mux_left_track_17.INVTX1_3_.out _0190_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_0929_ clknet_4_5_0_prog_clk mem_bottom_track_9.DFFR_0_.Q _0042_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_11.DFFR_0_.D sky130_fd_sc_hd__dfrtp_1
XFILLER_29_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0645_ net6 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.INVTX1_2_.out sky130_fd_sc_hd__inv_2
X_0714_ _0156_ vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__inv_2
XFILLER_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0576_ mem_right_track_16.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__inv_2
X_1128_ mux_bottom_track_7.INVTX1_0_.out _0242_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_40_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1059_ net143 _0173_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0430_ mem_bottom_track_23.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__clkbuf_1
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0628_ net67 vssd1 vssd1 vccd1 vccd1 mux_left_track_17.INVTX1_7_.out sky130_fd_sc_hd__inv_2
XFILLER_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0559_ mem_left_track_9.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__inv_2
XFILLER_26_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1047__142 vssd1 vssd1 vccd1 vccd1 net142 _1047__142/LO sky130_fd_sc_hd__conb_1
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0413_ _0130_ vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0962_ clknet_4_11_0_prog_clk mem_left_track_25.DFFR_7_.Q _0075_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_33.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
X_0893_ clknet_4_13_0_prog_clk mem_left_track_25.DFFR_4_.Q _0006_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_25.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1161_ mux_bottom_track_5.mux_2level_tapbuf_basis_input2_mem2_0_out _0275_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_5.mux_2level_tapbuf_basis_input3_mem3_1_out sky130_fd_sc_hd__ebufn_2
X_1092_ mux_right_track_24.INVTX1_0_.out _0206_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1230_ mux_left_track_1.INVTX1_3_.out _0344_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_52_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0876_ clknet_4_8_0_prog_clk mem_left_track_9.DFFR_5_.Q _0109_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_9.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
X_0945_ clknet_4_13_0_prog_clk mem_bottom_track_23.DFFR_0_.Q _0058_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_23.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_43_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0661_ net12 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_5.INVTX1_4_.out sky130_fd_sc_hd__inv_2
X_0730_ _0157_ vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__inv_2
XFILLER_6_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1213_ mux_bottom_track_25.INVTX1_0_.out _0327_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0592_ mem_right_track_8.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__inv_2
XFILLER_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1144_ mux_bottom_track_1.mux_2level_tapbuf_basis_input3_mem3_0_out _0258_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input3_mem3_1_out sky130_fd_sc_hd__ebufn_4
X_1075_ mux_right_track_16.INVTX1_1_.out _0189_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_0859_ clknet_4_2_0_prog_clk mem_right_track_16.DFFR_6_.Q _0092_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_16.DFFR_7_.Q sky130_fd_sc_hd__dfrtp_1
X_0928_ clknet_4_9_0_prog_clk mem_bottom_track_3.DFFR_5_.Q _0041_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_5.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0713_ _0156_ vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__inv_2
X_0644_ mux_bottom_track_1.mux_2level_tapbuf_basis_input3_mem3_1_out vssd1 vssd1 vccd1
+ vccd1 mux_bottom_track_1.out sky130_fd_sc_hd__inv_2
X_0575_ mem_right_track_16.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__inv_2
X_1127_ mux_left_track_25.INVTX1_4_.out _0241_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_25_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1058_ mux_bottom_track_23.INVTX1_2_.out _0172_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0627_ mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_17.out sky130_fd_sc_hd__clkinv_2
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0558_ mem_left_track_9.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__inv_2
X_0489_ mem_bottom_track_5.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__inv_2
XFILLER_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0412_ mem_bottom_track_27.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0961_ clknet_4_14_0_prog_clk mem_left_track_33.DFFR_0_.Q _0074_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_33.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_17_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0892_ clknet_4_13_0_prog_clk mem_left_track_25.DFFR_5_.Q _0005_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_25.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_4_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1160_ mux_bottom_track_5.INVTX1_4_.out _0274_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_5.mux_2level_tapbuf_basis_input2_mem2_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1091_ mux_left_track_9.INVTX1_5_.out _0205_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0944_ clknet_4_1_0_prog_clk mem_bottom_track_17.DFFR_1_.Q _0057_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_19.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_9_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0875_ clknet_4_8_0_prog_clk mem_left_track_9.DFFR_6_.Q _0108_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_17.DFFR_0_.D sky130_fd_sc_hd__dfrtp_1
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1154__152 vssd1 vssd1 vccd1 vccd1 net152 _1154__152/LO sky130_fd_sc_hd__conb_1
XFILLER_18_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0660_ net36 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_5.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0591_ mem_right_track_8.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__inv_2
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1212_ mux_bottom_track_25.INVTX1_2_.out _0326_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1143_ mux_bottom_track_1.INVTX1_2_.out _0257_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_18_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1074_ mux_bottom_track_15.INVTX1_1_.out _0188_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_0927_ clknet_4_12_0_prog_clk mem_bottom_track_5.DFFR_0_.Q _0040_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_5.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_2
X_0789_ _0124_ vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__inv_2
X_0858_ clknet_4_0_0_prog_clk mem_right_track_0.DFFR_7_.Q _0091_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_8.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_2
XFILLER_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0643_ net80 vssd1 vssd1 vccd1 vccd1 mux_right_track_32.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0574_ mem_right_track_16.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__inv_2
X_0712_ _0156_ vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__inv_2
Xclkbuf_4_4_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_4_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1126_ mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out _0240_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out sky130_fd_sc_hd__ebufn_4
XFILLER_40_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1057_ mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out _0171_ vssd1 vssd1
+ vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out sky130_fd_sc_hd__ebufn_4
XFILLER_31_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_46 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0557_ mem_left_track_9.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__inv_2
X_0626_ net71 vssd1 vssd1 vccd1 vccd1 mux_left_track_9.INVTX1_8_.out sky130_fd_sc_hd__inv_2
X_1109_ mux_left_track_17.INVTX1_6_.out _0223_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_0488_ mem_bottom_track_5.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__inv_2
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0411_ _0129_ vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0609_ net81 vssd1 vssd1 vccd1 vccd1 mux_right_track_0.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0960_ clknet_4_9_0_prog_clk mem_left_track_33.DFFR_1_.Q _0073_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_33.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
X_0891_ clknet_4_15_0_prog_clk mem_left_track_25.DFFR_6_.Q _0004_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_25.DFFR_7_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1235__166 vssd1 vssd1 vccd1 vccd1 net166 _1235__166/LO sky130_fd_sc_hd__conb_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1090_ mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out _0204_ vssd1
+ vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out sky130_fd_sc_hd__ebufn_4
X_0874_ clknet_4_9_0_prog_clk mem_right_track_16.DFFR_7_.Q _0107_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_24.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_2
X_0943_ clknet_4_6_0_prog_clk mem_bottom_track_19.DFFR_0_.Q _0056_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_19.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0590_ mem_right_track_16.DFFR_0_.D vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__inv_2
XFILLER_10_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1211_ mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_0_out _0325_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_2_out
+ sky130_fd_sc_hd__ebufn_1
X_1142_ mux_bottom_track_1.INVTX1_1_.out _0256_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1073_ mux_bottom_track_5.INVTX1_3_.out _0187_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_0857_ clknet_4_3_0_prog_clk mem_right_track_8.DFFR_0_.Q _0090_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_8.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
X_0926_ clknet_4_5_0_prog_clk mem_bottom_track_5.DFFR_1_.Q _0039_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_5.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0788_ _0155_ vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__buf_4
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0711_ _0155_ vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__buf_4
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0642_ net75 vssd1 vssd1 vccd1 vccd1 mux_right_track_32.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_0573_ mem_right_track_16.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__inv_2
XFILLER_38_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1125_ mux_left_track_25.INVTX1_3_.out _0239_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1056_ mux_right_track_0.INVTX1_0_.out _0170_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_33_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0909_ clknet_4_6_0_prog_clk mem_bottom_track_1.DFFR_0_.Q _0022_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_1.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_48_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1215__164 vssd1 vssd1 vccd1 vccd1 net164 _1215__164/LO sky130_fd_sc_hd__conb_1
XFILLER_62_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0625_ net44 vssd1 vssd1 vccd1 vccd1 mux_left_track_9.INVTX1_3_.out sky130_fd_sc_hd__inv_2
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0487_ mem_bottom_track_5.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__inv_2
X_0556_ mem_left_track_9.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__inv_2
XFILLER_53_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1108_ mux_left_track_17.INVTX1_5_.out _0222_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_26_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1039_ mux_bottom_track_11.out vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__clkbuf_1
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0410_ mem_bottom_track_27.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__clkbuf_1
X_0608_ mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out vssd1 vssd1 vccd1
+ vccd1 mux_right_track_0.out sky130_fd_sc_hd__inv_2
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0539_ mem_left_track_17.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__inv_2
XFILLER_26_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0890_ clknet_4_14_0_prog_clk mem_left_track_17.DFFR_0_.D _0003_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_17.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_2
XFILLER_4_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0873_ clknet_4_14_0_prog_clk mem_right_track_24.DFFR_0_.Q _0106_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_24.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_2
X_0942_ clknet_4_6_0_prog_clk mem_bottom_track_27.DFFR_1_.Q _0055_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_37.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1072_ mux_left_track_17.INVTX1_6_.out _0186_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1210_ mux_bottom_track_25.INVTX1_1_.out _0324_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_1_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1141_ net150 _0255_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1184__158 vssd1 vssd1 vccd1 vccd1 net158 _1184__158/LO sky130_fd_sc_hd__conb_1
X_0925_ clknet_4_1_0_prog_clk mem_bottom_track_5.DFFR_2_.Q _0038_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_5.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_1
X_0856_ clknet_4_11_0_prog_clk mem_right_track_8.DFFR_1_.Q _0089_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_8.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_2
X_0787_ _0123_ vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__inv_2
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0641_ mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out vssd1 vssd1 vccd1
+ vccd1 mux_right_track_32.out sky130_fd_sc_hd__inv_2
XFILLER_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0710_ net73 vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__buf_2
X_0572_ mem_right_track_24.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__inv_2
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1124_ mux_bottom_track_27.INVTX1_0_.out _0238_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1055_ mux_left_track_33.INVTX1_4_.out _0169_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_33_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0908_ clknet_4_0_0_prog_clk mem_bottom_track_1.DFFR_1_.Q _0021_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_1.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_1
X_0839_ _0128_ vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__inv_2
XFILLER_56_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0624_ net58 vssd1 vssd1 vccd1 vccd1 mux_left_track_9.INVTX1_4_.out sky130_fd_sc_hd__inv_2
XFILLER_7_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0486_ mem_bottom_track_5.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__inv_2
X_0555_ mem_left_track_9.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__inv_2
XFILLER_38_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1107_ net147 _0221_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1038_ mux_bottom_track_13.out vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0538_ mem_left_track_17.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__inv_2
X_0607_ mem_right_track_0.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__inv_2
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0469_ mem_bottom_track_13.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__inv_2
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1147__151 vssd1 vssd1 vccd1 vccd1 net151 _1147__151/LO sky130_fd_sc_hd__conb_1
X_0941_ clknet_4_7_0_prog_clk mem_bottom_track_37.DFFR_0_.Q _0054_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_37.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0872_ clknet_4_15_0_prog_clk mem_right_track_24.DFFR_1_.Q _0105_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_24.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1071_ net144 _0185_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1140_ mux_bottom_track_1.INVTX1_3_.out _0254_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0924_ clknet_4_7_0_prog_clk mem_bottom_track_5.DFFR_3_.Q _0037_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_5.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
X_0855_ clknet_4_14_0_prog_clk mem_right_track_8.DFFR_2_.Q _0088_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_8.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_2
X_0786_ _0123_ vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__inv_2
XFILLER_28_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0640_ net63 vssd1 vssd1 vccd1 vccd1 mux_left_track_25.INVTX1_8_.out sky130_fd_sc_hd__inv_2
X_0571_ mem_right_track_24.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__inv_2
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1123_ mux_bottom_track_17.INVTX1_0_.out _0237_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_25_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1054_ mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out _0168_ vssd1 vssd1
+ vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out sky130_fd_sc_hd__ebufn_4
X_0907_ clknet_4_2_0_prog_clk mem_bottom_track_1.DFFR_2_.Q _0020_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_1.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_1
X_0769_ _0122_ vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__inv_2
X_0838_ _0128_ vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__inv_2
XFILLER_0_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0623_ net45 vssd1 vssd1 vccd1 vccd1 mux_left_track_9.INVTX1_5_.out sky130_fd_sc_hd__inv_2
XFILLER_7_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0554_ mem_left_track_17.DFFR_0_.D vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__inv_2
X_1106_ mux_left_track_17.INVTX1_8_.out _0220_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_38_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0485_ _0154_ vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1037_ mux_bottom_track_15.out vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__clkbuf_1
XFILLER_21_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_3_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_3_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0537_ mem_left_track_17.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__inv_2
X_0606_ mem_right_track_0.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__inv_2
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0399_ mem_left_track_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__inv_2
XFILLER_26_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0468_ mem_bottom_track_13.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__inv_2
XFILLER_53_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0940_ clknet_4_14_0_prog_clk mem_bottom_track_19.DFFR_1_.Q _0053_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_21.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_13_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0871_ clknet_4_15_0_prog_clk mem_right_track_24.DFFR_2_.Q _0104_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_24.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1070_ mux_bottom_track_25.INVTX1_2_.out _0184_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0854_ clknet_4_3_0_prog_clk mem_right_track_8.DFFR_3_.Q _0087_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_8.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
X_0923_ clknet_4_13_0_prog_clk mem_bottom_track_5.DFFR_4_.Q _0036_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_5.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
X_0785_ _0123_ vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__inv_2
X_1199_ mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_0_out _0313_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_36_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0570_ mem_right_track_24.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__inv_2
X_1122_ mux_left_track_25.INVTX1_7_.out _0236_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_2_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1053_ mux_left_track_33.INVTX1_3_.out _0167_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_0837_ _0128_ vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__inv_2
X_0906_ clknet_4_10_0_prog_clk mem_bottom_track_1.DFFR_3_.Q _0019_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_1.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
X_0699_ net49 vssd1 vssd1 vccd1 vccd1 mux_left_track_1.INVTX1_5_.out sky130_fd_sc_hd__inv_2
X_0768_ _0122_ vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__inv_2
XFILLER_0_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0622_ net50 vssd1 vssd1 vccd1 vccd1 mux_left_track_9.INVTX1_6_.out sky130_fd_sc_hd__inv_2
X_0484_ mem_bottom_track_11.DFFR_0_.D vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0553_ mem_left_track_9.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__inv_2
XFILLER_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1105_ mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out _0219_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out sky130_fd_sc_hd__ebufn_4
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1036_ mux_bottom_track_17.out vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__clkbuf_1
Xinput80 right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net80 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0536_ mem_left_track_25.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__inv_2
X_0605_ mem_right_track_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__inv_2
X_0467_ _0148_ vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0398_ mem_left_track_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__inv_2
X_1019_ net20 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__clkbuf_1
XFILLER_57_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1083__145 vssd1 vssd1 vccd1 vccd1 net145 _1083__145/LO sky130_fd_sc_hd__conb_1
XFILLER_54_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0519_ mem_right_track_32.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__inv_2
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0870_ clknet_4_2_0_prog_clk mem_right_track_24.DFFR_3_.Q _0103_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_24.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_63_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0999_ net40 vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__clkbuf_2
XFILLER_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0922_ clknet_4_10_0_prog_clk mem_bottom_track_1.DFFR_5_.Q _0035_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_3.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_2
X_0853_ clknet_4_11_0_prog_clk mem_right_track_8.DFFR_4_.Q _0086_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_8.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
X_0784_ _0123_ vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__inv_2
XFILLER_56_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1198_ mux_bottom_track_1.INVTX1_1_.out _0312_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
Xinput1 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_ vssd1 vssd1 vccd1
+ vccd1 net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_28_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0_prog_clk prog_clk vssd1 vssd1 vccd1 vccd1 clknet_0_prog_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_47_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1121_ mux_left_track_25.INVTX1_6_.out _0235_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1052_ mux_left_track_33.INVTX1_2_.out _0166_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_21_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0767_ _0122_ vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__inv_2
X_0905_ clknet_4_10_0_prog_clk mem_bottom_track_1.DFFR_4_.Q _0018_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_1.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
X_0836_ _0128_ vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__inv_2
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0698_ net65 vssd1 vssd1 vccd1 vccd1 mux_left_track_1.INVTX1_6_.out sky130_fd_sc_hd__inv_2
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0621_ net66 vssd1 vssd1 vccd1 vccd1 mux_left_track_9.INVTX1_7_.out sky130_fd_sc_hd__inv_2
X_0483_ _0153_ vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__clkbuf_1
X_0552_ mem_left_track_9.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__inv_2
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1035_ mux_bottom_track_19.out vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__clkbuf_1
XFILLER_53_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1104_ mux_bottom_track_3.INVTX1_0_.out _0218_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_61_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput81 right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net81 sky130_fd_sc_hd__clkbuf_1
Xinput70 left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net70 sky130_fd_sc_hd__clkbuf_1
X_0819_ _0126_ vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__inv_2
XFILLER_29_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0604_ mem_right_track_0.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__inv_2
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0535_ mem_left_track_25.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__inv_2
X_0397_ mem_left_track_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__inv_2
X_0466_ mem_bottom_track_15.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1018_ net21 vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__clkbuf_2
XFILLER_26_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0518_ mem_bottom_track_1.DFFR_0_.D vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__inv_2
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0449_ _0142_ vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__clkbuf_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0998_ mux_left_track_17.out vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__clkbuf_1
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0921_ clknet_4_8_0_prog_clk mem_bottom_track_3.DFFR_0_.Q _0034_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_3.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_18_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0852_ clknet_4_11_0_prog_clk mem_right_track_8.DFFR_5_.Q _0085_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_8.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
X_0783_ _0123_ vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__inv_2
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1197_ net161 _0311_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput2 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_ vssd1 vssd1 vccd1
+ vccd1 net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1120_ mux_left_track_25.INVTX1_5_.out _0234_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1051_ mux_right_track_0.INVTX1_1_.out _0165_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0904_ clknet_4_3_0_prog_clk mem_right_track_24.DFFR_7_.Q _0017_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_32.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
X_0766_ _0155_ vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__buf_4
X_0697_ mux_left_track_1.mux_2level_tapbuf_basis_input3_mem3_3_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_1.out sky130_fd_sc_hd__inv_2
X_0835_ _0128_ vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__inv_2
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0620_ mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_9.out sky130_fd_sc_hd__inv_2
X_0551_ mem_left_track_9.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__inv_2
XFILLER_7_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0482_ mem_bottom_track_9.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1103_ mux_left_track_9.INVTX1_4_.out _0217_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1034_ mux_bottom_track_21.out vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__clkbuf_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput60 chany_bottom_in[7] vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_1
Xinput82 right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net82 sky130_fd_sc_hd__clkbuf_1
X_0749_ _0120_ vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__inv_2
Xinput71 left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net71 sky130_fd_sc_hd__clkbuf_1
X_0818_ _0126_ vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__inv_2
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0534_ mem_left_track_25.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__inv_2
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0603_ mem_right_track_0.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__inv_2
XFILLER_7_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0465_ _0147_ vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__clkbuf_1
X_0396_ mem_left_track_1.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__inv_2
XFILLER_26_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1017_ mux_right_track_16.out vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_2_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_2_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0517_ mem_right_track_32.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__inv_2
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0448_ mem_bottom_track_37.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__clkbuf_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0997_ net42 vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__clkbuf_1
XFILLER_46_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0920_ clknet_4_0_0_prog_clk mem_bottom_track_3.DFFR_1_.Q _0033_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_3.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0851_ clknet_4_11_0_prog_clk mem_right_track_8.DFFR_6_.Q _0084_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_16.DFFR_0_.D sky130_fd_sc_hd__dfrtp_1
X_0782_ _0123_ vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__inv_2
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput3 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_ vssd1 vssd1 vccd1
+ vccd1 net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1196_ mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_1_out _0310_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1050_ mux_bottom_track_11.INVTX1_1_.out _0164_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_18_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0903_ clknet_4_7_0_prog_clk mem_right_track_32.DFFR_0_.Q _0016_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_32.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
X_0834_ _0128_ vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__inv_2
X_0765_ _0121_ vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__inv_2
X_0696_ net14 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_27.INVTX1_2_.out sky130_fd_sc_hd__inv_2
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1179_ mux_bottom_track_13.INVTX1_0_.out _0293_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
Xclkbuf_4_15_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_15_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0550_ mem_left_track_9.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__inv_2
XFILLER_38_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0481_ mem_bottom_track_9.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__inv_2
X_1102_ mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out _0216_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out sky130_fd_sc_hd__ebufn_4
XFILLER_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1033_ mux_bottom_track_23.out vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__clkbuf_1
Xinput72 left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net72 sky130_fd_sc_hd__clkbuf_1
Xinput50 chany_bottom_in[15] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_1
Xinput61 chany_bottom_in[8] vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_1
X_0817_ _0126_ vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__inv_2
X_0748_ _0120_ vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__inv_2
X_0679_ net10 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_21.INVTX1_1_.out sky130_fd_sc_hd__inv_2
Xinput83 right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net83 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0533_ mem_left_track_25.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__inv_2
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0602_ mem_right_track_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__inv_2
X_0464_ mem_bottom_track_15.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0395_ mem_left_track_33.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__inv_2
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1016_ net23 vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0447_ _0141_ vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__clkbuf_1
X_0516_ mem_right_track_32.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__inv_2
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0996_ net43 vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0850_ clknet_4_10_0_prog_clk net5 _0083_ vssd1 vssd1 vccd1 vccd1 mem_right_track_0.DFFR_0_.Q
+ sky130_fd_sc_hd__dfrtp_2
X_0781_ _0123_ vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__inv_2
XFILLER_5_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput4 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_ vssd1 vssd1 vccd1
+ vccd1 net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1195_ mux_bottom_track_1.INVTX1_1_.out _0309_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_10_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0833_ _0128_ vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__inv_2
X_0902_ clknet_4_7_0_prog_clk mem_right_track_32.DFFR_1_.Q _0015_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_32.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_2
X_0695_ net33 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_27.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0764_ _0121_ vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__inv_2
XFILLER_24_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1178_ mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_0_out _0292_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_2
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0480_ mem_bottom_track_11.DFFR_0_.D vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__inv_2
XFILLER_38_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1032_ mux_bottom_track_25.out vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__clkbuf_1
X_1101_ mux_left_track_9.INVTX1_3_.out _0215_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
Xinput40 chanx_right_in[6] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_2
Xinput51 chany_bottom_in[16] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
X_0816_ _0126_ vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__inv_2
X_0747_ _0120_ vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__inv_2
Xinput62 chany_bottom_in[9] vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_1
Xinput73 pReset vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__dlymetal6s2s_1
X_0678_ net29 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_21.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_37_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0601_ mem_right_track_0.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__inv_2
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0394_ mem_left_track_33.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__inv_2
X_0532_ mem_left_track_25.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__inv_2
X_0463_ mem_bottom_track_15.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__inv_2
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1015_ net24 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0515_ mem_right_track_32.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__inv_2
X_0446_ mem_bottom_track_37.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__clkbuf_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0995_ net26 vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__clkbuf_1
XFILLER_5_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0429_ _0135_ vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__clkbuf_1
XFILLER_54_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0780_ _0123_ vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__inv_2
X_1194_ mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_0_out _0308_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_2
Xinput5 ccff_head vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0832_ net73 vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__buf_4
X_0763_ _0121_ vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__inv_2
X_0901_ clknet_4_1_0_prog_clk mem_right_track_32.DFFR_2_.Q _0014_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_32.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_1
X_0694_ net34 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_27.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1177_ mux_bottom_track_13.INVTX1_1_.out _0291_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_2_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1100_ mux_bottom_track_23.INVTX1_0_.out _0214_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1031_ mux_bottom_track_27.out vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__clkbuf_1
Xinput63 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_ vssd1 vssd1 vccd1
+ vccd1 net63 sky130_fd_sc_hd__clkbuf_1
Xinput52 chany_bottom_in[17] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_1
Xinput41 chanx_right_in[7] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput74 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_ vssd1 vssd1 vccd1
+ vccd1 net74 sky130_fd_sc_hd__clkbuf_1
Xinput30 chanx_right_in[14] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__dlymetal6s2s_1
X_0746_ _0120_ vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__inv_2
X_0815_ _0126_ vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__inv_2
XFILLER_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0677_ mux_bottom_track_21.mux_2level_tapbuf_basis_input2_mem1_1_out vssd1 vssd1
+ vccd1 vccd1 mux_bottom_track_21.out sky130_fd_sc_hd__inv_2
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1229_ mux_left_track_1.INVTX1_6_.out _0343_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_25_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1180__157 vssd1 vssd1 vccd1 vccd1 net157 _1180__157/LO sky130_fd_sc_hd__conb_1
XFILLER_4_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0531_ mem_left_track_25.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__inv_2
XFILLER_7_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0600_ mem_right_track_0.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__inv_2
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0462_ mem_bottom_track_15.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__inv_2
X_0393_ mem_left_track_33.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__inv_2
X_1014_ net7 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_1
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0729_ _0157_ vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__inv_2
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0514_ mem_right_track_32.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__inv_2
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0445_ mem_bottom_track_37.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__inv_2
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0994_ mux_left_track_25.out vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__clkbuf_1
XFILLER_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0428_ mem_bottom_track_23.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_1_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_1_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_18_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput6 chanx_left_in[0] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_2
XFILLER_36_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1193_ mux_bottom_track_37.INVTX1_1_.out _0307_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_32_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0900_ clknet_4_2_0_prog_clk mem_right_track_32.DFFR_3_.Q _0013_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_32.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0831_ _0127_ vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__inv_2
X_0693_ mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_2_out vssd1 vssd1
+ vccd1 vccd1 mux_bottom_track_27.out sky130_fd_sc_hd__inv_2
X_0762_ _0121_ vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__inv_2
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1176_ net156 _0290_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_20_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput140 net140 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[8] sky130_fd_sc_hd__buf_2
XFILLER_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1030_ net31 vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__clkbuf_2
XFILLER_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput31 chanx_right_in[15] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
Xinput20 chanx_left_in[5] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
X_0814_ _0126_ vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__inv_2
XFILLER_14_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput42 chanx_right_in[8] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput64 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_ vssd1 vssd1 vccd1
+ vccd1 net64 sky130_fd_sc_hd__clkbuf_1
X_0676_ net7 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.INVTX1_1_.out sky130_fd_sc_hd__inv_2
Xinput53 chany_bottom_in[18] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_1
Xinput75 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_ vssd1 vssd1 vccd1
+ vccd1 net75 sky130_fd_sc_hd__clkbuf_1
X_0745_ _0120_ vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__inv_2
X_1228_ mux_left_track_1.mux_2level_tapbuf_basis_input3_mem3_0_out _0342_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_52_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1159_ mux_bottom_track_3.INVTX1_0_.out _0273_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_3.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_4_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0530_ mem_left_track_25.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__inv_2
XFILLER_7_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0461_ _0146_ vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__clkbuf_1
X_0392_ mem_left_track_33.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__inv_2
XFILLER_34_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1013_ mux_right_track_24.out vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__clkbuf_1
XFILLER_8_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_14_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_14_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
X_0659_ net17 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_5.INVTX1_3_.out sky130_fd_sc_hd__inv_2
X_0728_ _0157_ vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__inv_2
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0444_ mem_bottom_track_37.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__inv_2
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0513_ mem_bottom_track_1.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__inv_2
XFILLER_39_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0993_ net28 vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__clkbuf_1
XFILLER_8_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0427_ mem_bottom_track_23.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__inv_2
XFILLER_39_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1192_ net160 _0306_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_36_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput7 chanx_left_in[10] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0830_ _0127_ vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__inv_2
X_0692_ net13 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.INVTX1_2_.out sky130_fd_sc_hd__inv_2
X_0761_ _0121_ vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__inv_2
XFILLER_49_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1175_ mux_bottom_track_11.INVTX1_0_.out _0289_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_24_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0959_ clknet_4_2_0_prog_clk mem_left_track_33.DFFR_2_.Q _0072_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_33.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput141 net141 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[9] sky130_fd_sc_hd__buf_2
Xoutput130 net130 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[16] sky130_fd_sc_hd__buf_2
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput54 chany_bottom_in[1] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_1
Xinput32 chanx_right_in[16] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_2
Xinput21 chanx_left_in[6] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_2
XFILLER_21_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0813_ _0126_ vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__inv_2
Xinput10 chanx_left_in[13] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput43 chanx_right_in[9] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput76 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net76 sky130_fd_sc_hd__clkbuf_1
X_0675_ net26 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0744_ _0155_ vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__buf_4
Xinput65 left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1227_ mux_bottom_track_21.INVTX1_0_.out _0341_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1158_ mux_bottom_track_3.mux_2level_tapbuf_basis_input3_mem3_0_out _0272_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_3.mux_2level_tapbuf_basis_input3_mem3_1_out sky130_fd_sc_hd__ebufn_2
XFILLER_52_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1089_ mux_left_track_9.INVTX1_4_.out _0203_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_20_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0460_ mem_bottom_track_17.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__clkbuf_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1012_ net9 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__clkbuf_1
X_0391_ mem_left_track_33.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__inv_2
XFILLER_34_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0727_ _0157_ vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__inv_2
X_0658_ mux_bottom_track_5.mux_2level_tapbuf_basis_input3_mem3_1_out vssd1 vssd1 vccd1
+ vccd1 mux_bottom_track_5.out sky130_fd_sc_hd__inv_2
X_0589_ mem_right_track_8.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__inv_2
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0443_ _0140_ vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0512_ mem_bottom_track_1.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__inv_2
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0992_ net29 vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__clkbuf_1
XFILLER_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0426_ mem_bottom_track_23.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__inv_2
X_1059__143 vssd1 vssd1 vccd1 vccd1 net143 _1059__143/LO sky130_fd_sc_hd__conb_1
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput8 chanx_left_in[11] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_46_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1191_ mux_bottom_track_21.INVTX1_0_.out _0305_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_21.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0409_ mem_bottom_track_27.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__inv_2
XFILLER_19_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0760_ _0121_ vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__inv_2
XFILLER_14_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0691_ net32 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_56_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1174_ mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_0_out _0288_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1243_ mux_bottom_track_9.INVTX1_0_.out _0357_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0958_ clknet_4_10_0_prog_clk mem_left_track_33.DFFR_3_.Q _0071_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_33.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
X_0889_ clknet_4_15_0_prog_clk mem_left_track_17.DFFR_0_.Q _0002_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_17.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput131 net131 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[17] sky130_fd_sc_hd__buf_2
Xoutput120 net120 vssd1 vssd1 vccd1 vccd1 chanx_right_out[7] sky130_fd_sc_hd__buf_2
XFILLER_28_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput33 chanx_right_in[17] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_2
Xinput55 chany_bottom_in[2] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
Xinput22 chanx_left_in[7] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
Xinput44 chany_bottom_in[0] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_1
X_0812_ _0126_ vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__inv_2
Xinput11 chanx_left_in[14] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput77 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net77 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput66 left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_1
X_0743_ _0158_ vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__inv_2
X_0674_ mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_1_out vssd1 vssd1
+ vccd1 vccd1 mux_bottom_track_17.out sky130_fd_sc_hd__inv_2
X_1226_ mux_bottom_track_11.INVTX1_0_.out _0340_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1157_ mux_bottom_track_3.INVTX1_3_.out _0271_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_3.mux_2level_tapbuf_basis_input2_mem2_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_52_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1088_ mux_left_track_9.INVTX1_3_.out _0202_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0390_ mem_left_track_33.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__inv_2
XFILLER_3_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1011_ net10 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__clkbuf_1
XFILLER_19_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0726_ _0157_ vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__inv_2
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0657_ net8 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_3.INVTX1_4_.out sky130_fd_sc_hd__inv_2
X_0588_ mem_right_track_8.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__inv_2
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1209_ net163 _0323_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0511_ mem_bottom_track_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__inv_2
X_0442_ mem_bottom_track_19.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0709_ net64 vssd1 vssd1 vccd1 vccd1 mux_left_track_33.INVTX1_7_.out sky130_fd_sc_hd__inv_2
XFILLER_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0991_ net30 vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0425_ _0134_ vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput9 chanx_left_in[12] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1190_ mux_bottom_track_21.mux_2level_tapbuf_basis_input2_mem1_0_out _0304_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_21.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_51_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0408_ mem_bottom_track_27.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__inv_2
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0690_ net2 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XFILLER_64_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1173_ mux_bottom_track_11.INVTX1_1_.out _0287_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1242_ mux_left_track_33.INVTX1_3_.out _0356_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput132 net132 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[18] sky130_fd_sc_hd__buf_2
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 chanx_right_out[15] sky130_fd_sc_hd__buf_2
Xoutput121 net121 vssd1 vssd1 vccd1 vccd1 chanx_right_out[8] sky130_fd_sc_hd__buf_2
X_0957_ clknet_4_10_0_prog_clk mem_left_track_33.DFFR_4_.Q _0070_ vssd1 vssd1 vccd1
+ vccd1 net84 sky130_fd_sc_hd__dfrtp_1
Xclkbuf_4_0_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_0_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0888_ clknet_4_13_0_prog_clk mem_left_track_17.DFFR_1_.Q _0001_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_17.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_2
XFILLER_21_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput78 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net78 sky130_fd_sc_hd__clkbuf_1
Xinput12 chanx_left_in[15] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
Xinput34 chanx_right_in[18] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_1
X_0811_ _0126_ vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__inv_2
Xinput45 chany_bottom_in[10] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_1
Xinput56 chany_bottom_in[3] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__clkbuf_1
X_0673_ net24 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_15.INVTX1_1_.out sky130_fd_sc_hd__inv_2
Xinput23 chanx_left_in[8] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput67 left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net67 sky130_fd_sc_hd__clkbuf_1
X_0742_ _0158_ vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__inv_2
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1225_ mux_left_track_1.INVTX1_5_.out _0339_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_25_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1087_ mux_right_track_24.INVTX1_1_.out _0201_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1156_ mux_bottom_track_23.INVTX1_1_.out _0270_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_3.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_20_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1010_ net11 vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0725_ _0157_ vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__inv_2
X_0656_ net35 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_3.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_57_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1208_ mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_1_out _0322_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_2_out
+ sky130_fd_sc_hd__ebufn_1
X_0587_ mem_right_track_8.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__inv_2
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1139_ mux_right_track_32.INVTX1_0_.out _0253_ vssd1 vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_63_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0510_ mem_bottom_track_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__inv_2
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0441_ mem_bottom_track_19.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__inv_2
XFILLER_39_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0639_ net55 vssd1 vssd1 vccd1 vccd1 mux_left_track_25.INVTX1_3_.out sky130_fd_sc_hd__inv_2
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0708_ net56 vssd1 vssd1 vccd1 vccd1 mux_left_track_33.INVTX1_2_.out sky130_fd_sc_hd__inv_2
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_13_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_13_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0990_ mux_left_track_33.out vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__clkbuf_1
X_0424_ mem_bottom_track_25.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1192__160 vssd1 vssd1 vccd1 vccd1 net160 _1192__160/LO sky130_fd_sc_hd__conb_1
XFILLER_6_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0407_ mem_left_track_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__inv_2
XFILLER_27_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1241_ mux_left_track_33.INVTX1_6_.out _0355_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1172_ net155 _0286_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0956_ clknet_4_12_0_prog_clk mem_bottom_track_37.DFFR_1_.Q _0069_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_1.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_2
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 chanx_right_out[16] sky130_fd_sc_hd__buf_2
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 chanx_left_out[6] sky130_fd_sc_hd__buf_2
Xoutput133 net133 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[1] sky130_fd_sc_hd__buf_2
X_0887_ clknet_4_5_0_prog_clk mem_left_track_17.DFFR_2_.Q _0000_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_17.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_1
Xoutput122 net122 vssd1 vssd1 vccd1 vccd1 chanx_right_out[9] sky130_fd_sc_hd__buf_2
XFILLER_15_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput13 chanx_left_in[16] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__dlymetal6s2s_1
X_0810_ _0155_ vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__clkbuf_8
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput79 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net79 sky130_fd_sc_hd__clkbuf_1
Xinput68 left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net68 sky130_fd_sc_hd__clkbuf_1
Xinput46 chany_bottom_in[11] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_1
Xinput35 chanx_right_in[1] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput57 chany_bottom_in[4] vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_1
X_0741_ _0158_ vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__inv_2
Xinput24 chanx_left_in[9] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
X_0672_ net43 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_15.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1224_ mux_left_track_1.INVTX1_4_.out _0338_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1086_ mux_bottom_track_17.INVTX1_1_.out _0200_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1155_ mux_bottom_track_3.INVTX1_1_.out _0269_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_3.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0939_ clknet_4_11_0_prog_clk mem_bottom_track_21.DFFR_0_.Q _0052_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_21.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0724_ _0157_ vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__inv_2
X_0586_ mem_right_track_8.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__inv_2
X_0655_ net4 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_3.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XFILLER_57_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1207_ mux_bottom_track_23.INVTX1_0_.out _0321_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_27_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1138_ mux_left_track_1.INVTX1_4_.out _0252_ vssd1 vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1069_ mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out _0183_ vssd1
+ vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out sky130_fd_sc_hd__ebufn_4
XFILLER_0_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0440_ _0139_ vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__clkbuf_1
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0707_ net61 vssd1 vssd1 vccd1 vccd1 mux_left_track_33.INVTX1_3_.out sky130_fd_sc_hd__inv_2
XFILLER_57_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0638_ net60 vssd1 vssd1 vccd1 vccd1 mux_left_track_25.INVTX1_4_.out sky130_fd_sc_hd__inv_2
X_0569_ mem_right_track_24.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__inv_2
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0423_ mem_bottom_track_25.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__inv_2
XFILLER_5_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1107__147 vssd1 vssd1 vccd1 vccd1 net147 _1107__147/LO sky130_fd_sc_hd__conb_1
XFILLER_24_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0406_ mem_left_track_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__inv_2
XFILLER_27_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1176__156 vssd1 vssd1 vccd1 vccd1 net156 _1176__156/LO sky130_fd_sc_hd__conb_1
XFILLER_42_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1171_ mux_bottom_track_9.INVTX1_0_.out _0285_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1240_ mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out _0354_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_64_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0886_ clknet_4_6_0_prog_clk mem_left_track_17.DFFR_3_.Q _0119_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_17.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
X_0955_ clknet_4_13_0_prog_clk mem_left_track_1.DFFR_0_.Q _0068_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_1.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
Xoutput134 net134 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[2] sky130_fd_sc_hd__buf_2
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 chanx_right_out[17] sky130_fd_sc_hd__buf_2
Xoutput123 net123 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[0] sky130_fd_sc_hd__buf_2
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 chanx_left_out[7] sky130_fd_sc_hd__buf_2
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput36 chanx_right_in[2] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput25 chanx_right_in[0] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_2
X_0740_ _0158_ vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__inv_2
Xinput14 chanx_left_in[17] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput58 chany_bottom_in[5] vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_1
Xinput69 left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_ vssd1 vssd1
+ vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput47 chany_bottom_in[12] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_1
X_0671_ mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_1_out vssd1 vssd1
+ vccd1 vccd1 mux_bottom_track_15.out sky130_fd_sc_hd__inv_2
X_1223_ net165 _0337_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1154_ net152 _0268_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_3.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1085_ mux_bottom_track_7.INVTX1_2_.out _0199_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_0869_ clknet_4_2_0_prog_clk mem_right_track_24.DFFR_4_.Q _0102_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_24.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
X_0938_ clknet_4_3_0_prog_clk mem_bottom_track_15.DFFR_1_.Q _0051_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_17.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0723_ _0157_ vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__inv_2
X_0585_ mem_right_track_8.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__inv_2
X_0654_ net16 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_3.INVTX1_3_.out sky130_fd_sc_hd__inv_2
XFILLER_6_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1137_ mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out _0251_ vssd1
+ vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out sky130_fd_sc_hd__ebufn_2
X_1206_ mux_bottom_track_23.INVTX1_2_.out _0320_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_25_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1068_ mux_right_track_8.INVTX1_0_.out _0182_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0706_ net48 vssd1 vssd1 vccd1 vccd1 mux_left_track_33.INVTX1_4_.out sky130_fd_sc_hd__inv_2
XFILLER_57_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0499_ mem_bottom_track_3.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__inv_2
X_0637_ net47 vssd1 vssd1 vccd1 vccd1 mux_left_track_25.INVTX1_5_.out sky130_fd_sc_hd__inv_2
X_0568_ mem_right_track_24.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__inv_2
XFILLER_53_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0422_ _0133_ vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0405_ mem_left_track_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__inv_2
XFILLER_50_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1170_ mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_0_out _0284_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_1_out sky130_fd_sc_hd__ebufn_2
XFILLER_2_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0885_ clknet_4_4_0_prog_clk mem_left_track_17.DFFR_4_.Q _0118_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_17.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
X_0954_ clknet_4_15_0_prog_clk mem_left_track_1.DFFR_1_.Q _0067_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_1.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_2
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 chanx_left_out[8] sky130_fd_sc_hd__buf_2
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 chanx_right_out[18] sky130_fd_sc_hd__buf_2
Xoutput124 net124 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[10] sky130_fd_sc_hd__buf_2
Xoutput135 net135 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[3] sky130_fd_sc_hd__buf_2
XFILLER_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput26 chanx_right_in[10] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_2
Xinput37 chanx_right_in[3] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_1
Xinput15 chanx_left_in[18] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
XFILLER_52_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0670_ net23 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_13.INVTX1_1_.out sky130_fd_sc_hd__inv_2
Xinput48 chany_bottom_in[13] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_1
Xinput59 chany_bottom_in[6] vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1222_ mux_left_track_1.INVTX1_7_.out _0336_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1084_ mux_left_track_9.INVTX1_6_.out _0198_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1153_ mux_bottom_track_3.mux_2level_tapbuf_basis_input2_mem2_0_out _0267_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_3.mux_2level_tapbuf_basis_input3_mem3_1_out sky130_fd_sc_hd__ebufn_2
X_0799_ _0155_ vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__buf_4
X_0868_ clknet_4_8_0_prog_clk mem_right_track_24.DFFR_5_.Q _0101_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_24.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0937_ clknet_4_5_0_prog_clk mem_bottom_track_17.DFFR_0_.Q _0050_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_17.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_43_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0722_ _0155_ vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__buf_4
X_0653_ mux_bottom_track_3.mux_2level_tapbuf_basis_input3_mem3_1_out vssd1 vssd1 vccd1
+ vccd1 mux_bottom_track_3.out sky130_fd_sc_hd__inv_2
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0584_ mem_right_track_16.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__inv_2
X_1136_ mux_bottom_track_19.INVTX1_2_.out _0250_ vssd1 vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input2_mem2_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1205_ mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_0_out _0319_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_25_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1067_ mux_left_track_25.INVTX1_5_.out _0181_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0636_ net52 vssd1 vssd1 vccd1 vccd1 mux_left_track_25.INVTX1_6_.out sky130_fd_sc_hd__inv_2
X_0705_ net53 vssd1 vssd1 vccd1 vccd1 mux_left_track_33.INVTX1_5_.out sky130_fd_sc_hd__inv_2
XFILLER_57_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0498_ mem_bottom_track_3.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__inv_2
X_0567_ mem_right_track_24.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__inv_2
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1119_ net148 _0233_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_21_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0421_ mem_bottom_track_25.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0619_ net79 vssd1 vssd1 vccd1 vccd1 mux_right_track_24.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0404_ mem_left_track_1.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__inv_2
XFILLER_50_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_12_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_12_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 chanx_left_out[9] sky130_fd_sc_hd__buf_2
Xoutput125 net125 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[11] sky130_fd_sc_hd__buf_2
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 chanx_right_out[1] sky130_fd_sc_hd__buf_2
X_0953_ clknet_4_11_0_prog_clk mem_left_track_1.DFFR_2_.Q _0066_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_1.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0884_ clknet_4_7_0_prog_clk mem_left_track_17.DFFR_5_.Q _0117_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_17.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
Xoutput136 net136 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[4] sky130_fd_sc_hd__buf_2
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput38 chanx_right_in[4] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput49 chany_bottom_in[14] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_1
Xinput16 chanx_left_in[1] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput27 chanx_right_in[11] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
X_1221_ mux_left_track_1.mux_2level_tapbuf_basis_input3_mem3_2_out _0335_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1152_ mux_bottom_track_3.INVTX1_4_.out _0266_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_3.mux_2level_tapbuf_basis_input2_mem2_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1083_ net145 _0197_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_0936_ clknet_4_0_0_prog_clk mem_bottom_track_13.DFFR_1_.Q _0049_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_15.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
X_0798_ _0124_ vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__inv_2
X_0867_ clknet_4_8_0_prog_clk mem_right_track_24.DFFR_6_.Q _0100_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_24.DFFR_7_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0652_ net15 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_7.INVTX1_3_.out sky130_fd_sc_hd__inv_2
X_0583_ mem_right_track_16.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__inv_2
X_0721_ _0156_ vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__inv_2
XFILLER_6_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1204_ mux_bottom_track_23.INVTX1_1_.out _0318_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_2_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1135_ mux_left_track_1.INVTX1_3_.out _0249_ vssd1 vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_25_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1066_ mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out _0180_ vssd1 vssd1
+ vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out sky130_fd_sc_hd__ebufn_4
X_0919_ clknet_4_2_0_prog_clk mem_bottom_track_3.DFFR_2_.Q _0032_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_3.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0635_ net68 vssd1 vssd1 vccd1 vccd1 mux_left_track_25.INVTX1_7_.out sky130_fd_sc_hd__inv_2
X_0704_ net69 vssd1 vssd1 vccd1 vccd1 mux_left_track_33.INVTX1_6_.out sky130_fd_sc_hd__inv_2
X_0566_ mem_right_track_24.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__inv_2
X_0497_ mem_bottom_track_3.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__inv_2
XFILLER_53_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1118_ mux_left_track_25.INVTX1_8_.out _0232_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1049_ mux_bottom_track_1.INVTX1_2_.out _0163_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_21_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0420_ _0132_ vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0618_ net74 vssd1 vssd1 vccd1 vccd1 mux_right_track_24.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_0549_ mem_left_track_9.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__inv_2
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0403_ mem_left_track_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__inv_2
XFILLER_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1095__146 vssd1 vssd1 vccd1 vccd1 net146 _1095__146/LO sky130_fd_sc_hd__conb_1
XFILLER_64_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0952_ clknet_4_10_0_prog_clk mem_left_track_1.DFFR_3_.Q _0065_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_1.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput126 net126 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[12] sky130_fd_sc_hd__buf_2
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 chanx_right_out[0] sky130_fd_sc_hd__buf_2
Xoutput137 net137 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[5] sky130_fd_sc_hd__buf_2
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 chanx_right_out[2] sky130_fd_sc_hd__buf_2
X_0883_ clknet_4_4_0_prog_clk mem_left_track_17.DFFR_6_.Q _0116_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_17.DFFR_7_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput17 chanx_left_in[2] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput28 chanx_right_in[12] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput39 chanx_right_in[5] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1151_ mux_bottom_track_7.INVTX1_0_.out _0265_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_7.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1220_ mux_left_track_1.mux_2level_tapbuf_basis_input3_mem3_1_out _0334_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1082_ mux_bottom_track_27.INVTX1_2_.out _0196_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0935_ clknet_4_0_0_prog_clk mem_bottom_track_15.DFFR_0_.Q _0048_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_15.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
X_0866_ clknet_4_15_0_prog_clk mem_right_track_16.DFFR_0_.D _0099_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_16.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
X_0797_ _0124_ vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__inv_2
XFILLER_28_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0720_ _0156_ vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__inv_2
X_0651_ net38 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_7.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0582_ mem_right_track_16.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__inv_2
X_1203_ net162 _0317_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
X_1134_ mux_right_track_32.INVTX1_1_.out _0248_ vssd1 vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1065_ mux_left_track_25.INVTX1_4_.out _0179_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_18_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0918_ clknet_4_11_0_prog_clk mem_bottom_track_3.DFFR_3_.Q _0031_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_3.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
X_0849_ clknet_4_15_0_prog_clk mem_right_track_0.DFFR_0_.Q _0082_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_0.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_2
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0703_ mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_33.out sky130_fd_sc_hd__inv_2
X_0634_ mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_25.out sky130_fd_sc_hd__inv_2
X_0496_ mem_bottom_track_3.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__inv_2
X_0565_ mem_right_track_24.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__inv_2
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1117_ mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out _0231_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out sky130_fd_sc_hd__ebufn_4
XFILLER_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1048_ mux_left_track_33.INVTX1_5_.out _0162_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0548_ mem_left_track_17.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__inv_2
X_0479_ _0152_ vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__clkbuf_1
X_0617_ mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out vssd1 vssd1 vccd1
+ vccd1 mux_right_track_24.out sky130_fd_sc_hd__clkinv_2
XFILLER_41_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0402_ mem_left_track_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__inv_2
XFILLER_35_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0882_ clknet_4_10_0_prog_clk mem_left_track_1.DFFR_5_.Q _0115_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_9.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_2
X_0951_ clknet_4_9_0_prog_clk mem_left_track_1.DFFR_4_.Q _0064_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_1.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 chanx_right_out[3] sky130_fd_sc_hd__buf_2
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput127 net127 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[13] sky130_fd_sc_hd__buf_2
Xoutput138 net138 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[6] sky130_fd_sc_hd__buf_2
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 chanx_right_out[10] sky130_fd_sc_hd__buf_2
XFILLER_55_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_10 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput18 chanx_left_in[3] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
Xinput29 chanx_right_in[13] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1150_ mux_bottom_track_7.mux_2level_tapbuf_basis_input3_mem3_0_out _0264_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_7.mux_2level_tapbuf_basis_input3_mem3_1_out sky130_fd_sc_hd__ebufn_2
XFILLER_45_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1081_ mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out _0195_ vssd1
+ vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out sky130_fd_sc_hd__ebufn_4
X_0934_ clknet_4_1_0_prog_clk mem_bottom_track_11.DFFR_1_.Q _0047_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_13.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_1
X_0865_ clknet_4_4_0_prog_clk mem_right_track_16.DFFR_0_.Q _0098_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_16.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0796_ _0124_ vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__inv_2
XFILLER_43_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0650_ net19 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_7.INVTX1_2_.out sky130_fd_sc_hd__inv_2
X_0581_ mem_right_track_16.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__inv_2
XFILLER_2_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1064_ mux_left_track_25.INVTX1_3_.out _0178_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1202_ mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_1_out _0316_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1133_ mux_bottom_track_9.INVTX1_1_.out _0247_ vssd1 vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0779_ _0123_ vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__inv_2
X_0917_ clknet_4_11_0_prog_clk mem_bottom_track_3.DFFR_4_.Q _0030_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_3.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
X_0848_ clknet_4_12_0_prog_clk mem_right_track_0.DFFR_1_.Q _0081_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_0.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0702_ net70 vssd1 vssd1 vccd1 vccd1 mux_left_track_1.INVTX1_7_.out sky130_fd_sc_hd__inv_2
X_0633_ net72 vssd1 vssd1 vccd1 vccd1 mux_left_track_17.INVTX1_8_.out sky130_fd_sc_hd__inv_2
X_0564_ mem_right_track_24.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__inv_2
X_0495_ mem_bottom_track_3.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__inv_2
XFILLER_38_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1116_ mux_bottom_track_5.INVTX1_0_.out _0230_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_4_9_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_9_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1047_ net142 _0161_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0616_ net78 vssd1 vssd1 vccd1 vccd1 mux_right_track_16.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0547_ mem_left_track_17.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__inv_2
X_0478_ mem_bottom_track_11.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0401_ mem_left_track_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__inv_2
XFILLER_4_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0881_ clknet_4_9_0_prog_clk mem_left_track_9.DFFR_0_.Q _0114_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_9.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_2
XFILLER_9_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0950_ clknet_4_15_0_prog_clk mem_bottom_track_25.DFFR_1_.Q _0063_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_27.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 chanx_right_out[4] sky130_fd_sc_hd__buf_2
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 chanx_right_out[11] sky130_fd_sc_hd__buf_2
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput128 net128 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[14] sky130_fd_sc_hd__buf_2
Xoutput139 net139 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[7] sky130_fd_sc_hd__buf_2
XFILLER_55_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput19 chanx_left_in[4] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_11_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_11_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1080_ mux_right_track_16.INVTX1_0_.out _0194_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0933_ clknet_4_0_0_prog_clk mem_bottom_track_13.DFFR_0_.Q _0046_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_13.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
X_0795_ _0124_ vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__inv_2
XFILLER_13_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0864_ clknet_4_5_0_prog_clk mem_right_track_16.DFFR_1_.Q _0097_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_16.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1201_ mux_bottom_track_19.INVTX1_0_.out _0315_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_0580_ mem_right_track_16.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__inv_2
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1132_ mux_left_track_1.INVTX1_5_.out _0246_ vssd1 vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1063_ mux_right_track_8.INVTX1_1_.out _0177_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_33_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0916_ clknet_4_14_0_prog_clk mem_bottom_track_5.DFFR_5_.Q _0029_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_7.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_1
X_0847_ clknet_4_14_0_prog_clk mem_right_track_0.DFFR_2_.Q _0080_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_0.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_2
X_0778_ _0123_ vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__inv_2
XFILLER_56_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0632_ net54 vssd1 vssd1 vccd1 vccd1 mux_left_track_17.INVTX1_3_.out sky130_fd_sc_hd__inv_2
X_0701_ net57 vssd1 vssd1 vccd1 vccd1 mux_left_track_1.INVTX1_3_.out sky130_fd_sc_hd__inv_2
X_0563_ mem_right_track_24.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__inv_2
XFILLER_38_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0494_ mem_bottom_track_3.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__inv_2
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1115_ mux_left_track_17.INVTX1_4_.out _0229_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1046_ mux_bottom_track_21.INVTX1_1_.out _0160_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_0_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0546_ mem_left_track_17.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__inv_2
XFILLER_7_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0615_ net83 vssd1 vssd1 vccd1 vccd1 mux_right_track_16.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0477_ _0151_ vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1029_ net27 vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__clkbuf_1
XFILLER_30_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0400_ mem_left_track_1.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__inv_2
XFILLER_35_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0529_ mem_left_track_25.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__inv_2
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 chanx_right_out[12] sky130_fd_sc_hd__buf_2
XFILLER_9_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0880_ clknet_4_14_0_prog_clk mem_left_track_9.DFFR_1_.Q _0113_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_9.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_2
XFILLER_13_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 chanx_right_out[5] sky130_fd_sc_hd__buf_2
Xoutput129 net129 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[15] sky130_fd_sc_hd__buf_2
XFILLER_23_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0932_ clknet_4_7_0_prog_clk mem_bottom_track_11.DFFR_0_.D _0045_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_11.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0794_ _0124_ vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__inv_2
X_0863_ clknet_4_7_0_prog_clk mem_right_track_16.DFFR_2_.Q _0096_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_16.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_2
XFILLER_51_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1200_ mux_bottom_track_19.INVTX1_2_.out _0314_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_1
X_1131_ mux_right_track_32.mux_2level_tapbuf_basis_input2_mem2_0_out _0245_ vssd1
+ vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out sky130_fd_sc_hd__ebufn_2
X_1062_ mux_bottom_track_13.INVTX1_1_.out _0176_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0915_ clknet_4_3_0_prog_clk mem_bottom_track_7.DFFR_0_.Q _0028_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_7.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
X_0846_ clknet_4_3_0_prog_clk mem_right_track_0.DFFR_3_.Q _0079_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_0.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0777_ _0155_ vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__buf_4
XFILLER_56_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0700_ net62 vssd1 vssd1 vccd1 vccd1 mux_left_track_1.INVTX1_4_.out sky130_fd_sc_hd__inv_2
X_0562_ mem_right_track_24.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__inv_2
X_0631_ net59 vssd1 vssd1 vccd1 vccd1 mux_left_track_17.INVTX1_4_.out sky130_fd_sc_hd__inv_2
XFILLER_53_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0493_ mem_bottom_track_5.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__inv_2
X_1114_ mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out _0228_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out sky130_fd_sc_hd__ebufn_4
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1045_ mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out _0159_ vssd1 vssd1
+ vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out sky130_fd_sc_hd__ebufn_4
X_1162__153 vssd1 vssd1 vccd1 vccd1 net153 _1162__153/LO sky130_fd_sc_hd__conb_1
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0829_ _0127_ vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__inv_2
XFILLER_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0476_ mem_bottom_track_11.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__clkbuf_1
X_0545_ mem_left_track_17.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__inv_2
X_0614_ mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out vssd1 vssd1 vccd1
+ vccd1 mux_right_track_16.out sky130_fd_sc_hd__inv_2
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1028_ net41 vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__clkbuf_2
XFILLER_29_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0528_ mem_left_track_25.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__inv_2
X_0459_ _0145_ vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__clkbuf_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 chanx_right_out[13] sky130_fd_sc_hd__buf_2
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 chanx_right_out[6] sky130_fd_sc_hd__buf_2
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 chanx_left_out[14] sky130_fd_sc_hd__buf_2
XFILLER_23_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0862_ clknet_4_0_0_prog_clk mem_right_track_16.DFFR_3_.Q _0095_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_16.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
X_0931_ clknet_4_1_0_prog_clk mem_bottom_track_11.DFFR_0_.Q _0044_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_11.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0793_ _0124_ vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__inv_2
XFILLER_51_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1172__155 vssd1 vssd1 vccd1 vccd1 net155 _1172__155/LO sky130_fd_sc_hd__conb_1
XFILLER_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1130_ mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out _0244_ vssd1
+ vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out sky130_fd_sc_hd__ebufn_2
X_1061_ mux_bottom_track_3.INVTX1_3_.out _0175_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_0914_ clknet_4_0_0_prog_clk mem_bottom_track_7.DFFR_1_.Q _0027_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_7.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_1
X_0845_ clknet_4_0_0_prog_clk mem_right_track_0.DFFR_4_.Q _0078_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_0.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
X_0776_ _0122_ vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__inv_2
XFILLER_17_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0630_ net46 vssd1 vssd1 vccd1 vccd1 mux_left_track_17.INVTX1_5_.out sky130_fd_sc_hd__inv_2
X_0492_ mem_bottom_track_5.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__inv_2
X_0561_ mem_right_track_24.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__inv_2
XFILLER_53_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1113_ mux_left_track_17.INVTX1_3_.out _0227_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1044_ mux_bottom_track_1.out vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__clkbuf_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1203__162 vssd1 vssd1 vccd1 vccd1 net162 _1203__162/LO sky130_fd_sc_hd__conb_1
X_0828_ _0127_ vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__inv_2
X_0759_ _0121_ vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__inv_2
XFILLER_56_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0613_ net77 vssd1 vssd1 vccd1 vccd1 mux_right_track_8.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_11_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0475_ mem_bottom_track_11.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__inv_2
X_0544_ mem_left_track_17.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__inv_2
X_1027_ net37 vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__clkbuf_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_8_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_8_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_4_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0527_ mem_left_track_25.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__inv_2
X_0458_ mem_bottom_track_17.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0145_ sky130_fd_sc_hd__clkbuf_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0389_ mem_left_track_33.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__inv_2
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1223__165 vssd1 vssd1 vccd1 vccd1 net165 _1223__165/LO sky130_fd_sc_hd__conb_1
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 chanx_right_out[14] sky130_fd_sc_hd__buf_2
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 chanx_left_out[15] sky130_fd_sc_hd__buf_2
XFILLER_36_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0930_ clknet_4_1_0_prog_clk mem_bottom_track_7.DFFR_5_.Q _0043_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_9.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_1
X_0861_ clknet_4_0_0_prog_clk mem_right_track_16.DFFR_4_.Q _0094_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_16.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0792_ _0124_ vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__inv_2
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1060_ mux_left_track_25.INVTX1_6_.out _0174_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_2_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0844_ clknet_4_0_0_prog_clk mem_right_track_0.DFFR_5_.Q _0077_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_0.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
X_0913_ clknet_4_1_0_prog_clk mem_bottom_track_7.DFFR_2_.Q _0026_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_7.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_1
X_0775_ _0122_ vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__inv_2
X_1189_ mux_bottom_track_21.INVTX1_1_.out _0303_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_21.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_10_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_10_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_3_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0560_ mem_left_track_9.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__inv_2
X_0491_ mem_bottom_track_5.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__inv_2
XFILLER_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1112_ mux_bottom_track_25.INVTX1_0_.out _0226_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1043_ mux_bottom_track_3.out vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__clkbuf_1
XFILLER_61_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0758_ _0121_ vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__inv_2
X_0827_ _0127_ vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__inv_2
X_0689_ mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_2_out vssd1 vssd1
+ vccd1 vccd1 mux_bottom_track_25.out sky130_fd_sc_hd__inv_2
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0612_ net82 vssd1 vssd1 vccd1 vccd1 mux_right_track_8.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0543_ mem_left_track_17.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__inv_2
X_0474_ mem_bottom_track_11.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__inv_2
XFILLER_53_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1026_ mux_bottom_track_37.out vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__clkbuf_1
XFILLER_61_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0526_ mem_left_track_25.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__inv_2
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0457_ mem_bottom_track_17.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__inv_2
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0388_ net84 vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__inv_2
X_1009_ mux_right_track_32.out vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__clkbuf_1
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 chanx_left_out[16] sky130_fd_sc_hd__buf_2
XFILLER_51_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0509_ mem_bottom_track_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__inv_2
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0791_ _0124_ vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__inv_2
X_0860_ clknet_4_0_0_prog_clk mem_right_track_16.DFFR_5_.Q _0093_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_16.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_36_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0989_ net32 vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__clkbuf_1
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0912_ clknet_4_4_0_prog_clk mem_bottom_track_7.DFFR_3_.Q _0025_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_7.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0774_ _0122_ vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__inv_2
X_0843_ clknet_4_0_0_prog_clk mem_right_track_0.DFFR_6_.Q _0076_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_0.DFFR_7_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1188_ net159 _0302_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_21.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0490_ mem_bottom_track_5.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__inv_2
XFILLER_2_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1042_ mux_bottom_track_5.out vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__clkbuf_1
X_1111_ mux_bottom_track_15.INVTX1_0_.out _0225_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_61_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0688_ net11 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_23.INVTX1_2_.out sky130_fd_sc_hd__inv_2
X_0757_ _0121_ vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__inv_2
X_0826_ _0127_ vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__inv_2
XFILLER_29_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0611_ mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out vssd1 vssd1 vccd1
+ vccd1 mux_right_track_8.out sky130_fd_sc_hd__inv_2
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0542_ mem_left_track_17.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__inv_2
XFILLER_7_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0473_ _0150_ vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1025_ mux_right_track_0.out vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__clkbuf_1
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0809_ _0125_ vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__inv_2
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0456_ mem_bottom_track_17.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__inv_2
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0525_ mem_left_track_25.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__inv_2
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0387_ mem_left_track_33.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__inv_2
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1008_ net13 vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__clkbuf_1
XFILLER_22_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 chanx_left_out[17] sky130_fd_sc_hd__buf_2
XFILLER_63_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0439_ mem_bottom_track_19.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0508_ mem_bottom_track_1.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__inv_2
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0790_ _0124_ vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__inv_2
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0988_ net33 vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__clkbuf_1
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0842_ _0128_ vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__inv_2
X_0911_ clknet_4_4_0_prog_clk mem_bottom_track_7.DFFR_4_.Q _0024_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_7.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0773_ _0122_ vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__inv_2
XFILLER_5_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1187_ mux_bottom_track_17.INVTX1_0_.out _0301_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1110_ mux_left_track_17.INVTX1_7_.out _0224_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_0_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1041_ mux_bottom_track_7.out vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__clkbuf_1
X_0825_ _0127_ vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__inv_2
X_0687_ net30 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_23.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0756_ _0121_ vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__inv_2
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1239_ mux_left_track_33.INVTX1_2_.out _0353_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0610_ net76 vssd1 vssd1 vccd1 vccd1 mux_right_track_0.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0541_ mem_left_track_17.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__inv_2
X_0472_ mem_bottom_track_13.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__clkbuf_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1024_ net6 vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__clkbuf_1
XFILLER_38_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0808_ _0125_ vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__inv_2
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0739_ _0158_ vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__inv_2
XFILLER_44_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_2 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0524_ mem_right_track_32.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__inv_2
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0455_ _0144_ vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0386_ mem_left_track_33.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__inv_2
X_1007_ net14 vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__clkbuf_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 chanx_left_out[18] sky130_fd_sc_hd__buf_2
XFILLER_49_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0438_ _0138_ vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0507_ mem_bottom_track_7.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__inv_2
XFILLER_54_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_7_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_7_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0772_ _0122_ vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__inv_2
X_0841_ _0128_ vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__inv_2
X_0910_ clknet_4_7_0_prog_clk mem_bottom_track_1.DFFR_0_.D _0023_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_1.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1186_ mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_0_out _0300_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1040_ mux_bottom_track_9.out vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__clkbuf_1
XFILLER_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0755_ _0155_ vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__buf_4
X_0824_ _0127_ vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__inv_2
X_0686_ net1 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_23.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1169_ mux_bottom_track_9.INVTX1_1_.out _0283_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1238_ mux_bottom_track_19.INVTX1_0_.out _0352_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0540_ mem_left_track_17.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__inv_2
X_0471_ _0149_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1023_ net16 vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__clkbuf_1
XFILLER_19_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0807_ _0125_ vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__inv_2
X_0738_ _0158_ vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__inv_2
X_0669_ net42 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_13.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_39_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0523_ mem_right_track_32.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__inv_2
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0454_ mem_bottom_track_21.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__clkbuf_1
X_0385_ mem_left_track_33.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__inv_2
XFILLER_22_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1006_ mux_left_track_1.out vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__clkbuf_1
XFILLER_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1071__144 vssd1 vssd1 vccd1 vccd1 net144 _1071__144/LO sky130_fd_sc_hd__conb_1
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 chanx_left_out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 ccff_tail sky130_fd_sc_hd__buf_2
XFILLER_63_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0506_ mem_bottom_track_7.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__inv_2
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0437_ mem_bottom_track_19.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0840_ _0128_ vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__inv_2
X_0771_ _0122_ vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__inv_2
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1185_ mux_bottom_track_17.INVTX1_1_.out _0299_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_24_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0685_ mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_2_out vssd1 vssd1
+ vccd1 vccd1 mux_bottom_track_23.out sky130_fd_sc_hd__inv_2
X_0754_ _0120_ vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__inv_2
X_0823_ _0127_ vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__inv_2
XFILLER_52_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1168_ net154 _0282_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1237_ mux_left_track_33.INVTX1_5_.out _0351_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1099_ mux_bottom_track_13.INVTX1_0_.out _0213_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_20_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0470_ mem_bottom_track_13.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__clkbuf_1
X_1022_ net17 vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__clkbuf_2
XFILLER_34_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0668_ mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_1_out vssd1 vssd1
+ vccd1 vccd1 mux_bottom_track_13.out sky130_fd_sc_hd__inv_2
X_0806_ _0125_ vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__inv_2
X_0737_ _0158_ vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__inv_2
X_0599_ mem_right_track_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__inv_2
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0522_ mem_right_track_32.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__inv_2
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0453_ _0143_ vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__clkbuf_1
X_0384_ mem_left_track_33.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__inv_2
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1129__149 vssd1 vssd1 vccd1 vccd1 net149 _1129__149/LO sky130_fd_sc_hd__conb_1
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1168__154 vssd1 vssd1 vccd1 vccd1 net154 _1168__154/LO sky130_fd_sc_hd__conb_1
X_1005_ net25 vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__clkbuf_1
XFILLER_22_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 chanx_left_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 chanx_left_out[0] sky130_fd_sc_hd__buf_2
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0436_ mem_bottom_track_19.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__inv_2
X_0505_ mem_bottom_track_7.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__inv_2
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

