magic
tech sky130A
magscale 1 2
timestamp 1674174156
<< obsli1 >>
rect 1104 2159 36892 37553
<< obsm1 >>
rect 14 1300 37430 37664
<< metal2 >>
rect 662 39200 718 39800
rect 2594 39200 2650 39800
rect 4526 39200 4582 39800
rect 5814 39200 5870 39800
rect 7746 39200 7802 39800
rect 9678 39200 9734 39800
rect 10966 39200 11022 39800
rect 12898 39200 12954 39800
rect 14830 39200 14886 39800
rect 16118 39200 16174 39800
rect 18050 39200 18106 39800
rect 19982 39200 20038 39800
rect 21270 39200 21326 39800
rect 23202 39200 23258 39800
rect 25134 39200 25190 39800
rect 26422 39200 26478 39800
rect 28354 39200 28410 39800
rect 30286 39200 30342 39800
rect 31574 39200 31630 39800
rect 33506 39200 33562 39800
rect 35438 39200 35494 39800
rect 36726 39200 36782 39800
rect 18 200 74 800
rect 1306 200 1362 800
rect 3238 200 3294 800
rect 4526 200 4582 800
rect 6458 200 6514 800
rect 8390 200 8446 800
rect 9678 200 9734 800
rect 11610 200 11666 800
rect 13542 200 13598 800
rect 14830 200 14886 800
rect 16762 200 16818 800
rect 18694 200 18750 800
rect 19982 200 20038 800
rect 21914 200 21970 800
rect 23846 200 23902 800
rect 25134 200 25190 800
rect 27066 200 27122 800
rect 28998 200 29054 800
rect 30286 200 30342 800
rect 32218 200 32274 800
rect 34150 200 34206 800
rect 35438 200 35494 800
rect 37370 200 37426 800
<< obsm2 >>
rect 20 39144 606 39545
rect 774 39144 2538 39545
rect 2706 39144 4470 39545
rect 4638 39144 5758 39545
rect 5926 39144 7690 39545
rect 7858 39144 9622 39545
rect 9790 39144 10910 39545
rect 11078 39144 12842 39545
rect 13010 39144 14774 39545
rect 14942 39144 16062 39545
rect 16230 39144 17994 39545
rect 18162 39144 19926 39545
rect 20094 39144 21214 39545
rect 21382 39144 23146 39545
rect 23314 39144 25078 39545
rect 25246 39144 26366 39545
rect 26534 39144 28298 39545
rect 28466 39144 30230 39545
rect 30398 39144 31518 39545
rect 31686 39144 33450 39545
rect 33618 39144 35382 39545
rect 35550 39144 36670 39545
rect 36838 39144 37424 39545
rect 20 856 37424 39144
rect 130 711 1250 856
rect 1418 711 3182 856
rect 3350 711 4470 856
rect 4638 711 6402 856
rect 6570 711 8334 856
rect 8502 711 9622 856
rect 9790 711 11554 856
rect 11722 711 13486 856
rect 13654 711 14774 856
rect 14942 711 16706 856
rect 16874 711 18638 856
rect 18806 711 19926 856
rect 20094 711 21858 856
rect 22026 711 23790 856
rect 23958 711 25078 856
rect 25246 711 27010 856
rect 27178 711 28942 856
rect 29110 711 30230 856
rect 30398 711 32162 856
rect 32330 711 34094 856
rect 34262 711 35382 856
rect 35550 711 37314 856
<< metal3 >>
rect 200 39448 800 39568
rect 37200 38768 37800 38888
rect 200 37408 800 37528
rect 37200 37408 37800 37528
rect 200 36048 800 36168
rect 37200 35368 37800 35488
rect 200 34008 800 34128
rect 37200 33328 37800 33448
rect 200 31968 800 32088
rect 37200 31968 37800 32088
rect 200 30608 800 30728
rect 37200 29928 37800 30048
rect 200 28568 800 28688
rect 37200 27888 37800 28008
rect 200 26528 800 26648
rect 37200 26528 37800 26648
rect 200 25168 800 25288
rect 37200 24488 37800 24608
rect 200 23128 800 23248
rect 37200 22448 37800 22568
rect 200 21088 800 21208
rect 37200 21088 37800 21208
rect 200 19728 800 19848
rect 37200 19048 37800 19168
rect 200 17688 800 17808
rect 37200 17008 37800 17128
rect 200 15648 800 15768
rect 37200 15648 37800 15768
rect 200 14288 800 14408
rect 37200 13608 37800 13728
rect 200 12248 800 12368
rect 37200 11568 37800 11688
rect 200 10208 800 10328
rect 37200 10208 37800 10328
rect 200 8848 800 8968
rect 37200 8168 37800 8288
rect 200 6808 800 6928
rect 37200 6128 37800 6248
rect 200 4768 800 4888
rect 37200 4768 37800 4888
rect 200 3408 800 3528
rect 37200 2728 37800 2848
rect 200 1368 800 1488
rect 37200 688 37800 808
<< obsm3 >>
rect 880 39368 37200 39541
rect 800 38968 37200 39368
rect 800 38688 37120 38968
rect 800 37608 37200 38688
rect 880 37328 37120 37608
rect 800 36248 37200 37328
rect 880 35968 37200 36248
rect 800 35568 37200 35968
rect 800 35288 37120 35568
rect 800 34208 37200 35288
rect 880 33928 37200 34208
rect 800 33528 37200 33928
rect 800 33248 37120 33528
rect 800 32168 37200 33248
rect 880 31888 37120 32168
rect 800 30808 37200 31888
rect 880 30528 37200 30808
rect 800 30128 37200 30528
rect 800 29848 37120 30128
rect 800 28768 37200 29848
rect 880 28488 37200 28768
rect 800 28088 37200 28488
rect 800 27808 37120 28088
rect 800 26728 37200 27808
rect 880 26448 37120 26728
rect 800 25368 37200 26448
rect 880 25088 37200 25368
rect 800 24688 37200 25088
rect 800 24408 37120 24688
rect 800 23328 37200 24408
rect 880 23048 37200 23328
rect 800 22648 37200 23048
rect 800 22368 37120 22648
rect 800 21288 37200 22368
rect 880 21008 37120 21288
rect 800 19928 37200 21008
rect 880 19648 37200 19928
rect 800 19248 37200 19648
rect 800 18968 37120 19248
rect 800 17888 37200 18968
rect 880 17608 37200 17888
rect 800 17208 37200 17608
rect 800 16928 37120 17208
rect 800 15848 37200 16928
rect 880 15568 37120 15848
rect 800 14488 37200 15568
rect 880 14208 37200 14488
rect 800 13808 37200 14208
rect 800 13528 37120 13808
rect 800 12448 37200 13528
rect 880 12168 37200 12448
rect 800 11768 37200 12168
rect 800 11488 37120 11768
rect 800 10408 37200 11488
rect 880 10128 37120 10408
rect 800 9048 37200 10128
rect 880 8768 37200 9048
rect 800 8368 37200 8768
rect 800 8088 37120 8368
rect 800 7008 37200 8088
rect 880 6728 37200 7008
rect 800 6328 37200 6728
rect 800 6048 37120 6328
rect 800 4968 37200 6048
rect 880 4688 37120 4968
rect 800 3608 37200 4688
rect 880 3328 37200 3608
rect 800 2928 37200 3328
rect 800 2648 37120 2928
rect 800 1568 37200 2648
rect 880 1288 37200 1568
rect 800 888 37200 1288
rect 800 715 37120 888
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< obsm4 >>
rect 5947 18803 10613 36005
<< labels >>
rlabel metal3 s 200 19728 800 19848 6 bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_
port 1 nsew signal output
rlabel metal3 s 37200 33328 37800 33448 6 bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_
port 2 nsew signal output
rlabel metal3 s 37200 8168 37800 8288 6 bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_
port 3 nsew signal output
rlabel metal2 s 27066 200 27122 800 6 bottom_grid_top_width_0_height_0_subtile_0__pin_clk_0_
port 4 nsew signal output
rlabel metal3 s 37200 31968 37800 32088 6 ccff_head
port 5 nsew signal input
rlabel metal3 s 37200 24488 37800 24608 6 ccff_tail
port 6 nsew signal output
rlabel metal2 s 16118 39200 16174 39800 6 chanx_left_in[0]
port 7 nsew signal input
rlabel metal2 s 14830 39200 14886 39800 6 chanx_left_in[10]
port 8 nsew signal input
rlabel metal3 s 37200 15648 37800 15768 6 chanx_left_in[11]
port 9 nsew signal input
rlabel metal2 s 662 39200 718 39800 6 chanx_left_in[12]
port 10 nsew signal input
rlabel metal3 s 200 4768 800 4888 6 chanx_left_in[13]
port 11 nsew signal input
rlabel metal3 s 200 36048 800 36168 6 chanx_left_in[14]
port 12 nsew signal input
rlabel metal2 s 13542 200 13598 800 6 chanx_left_in[15]
port 13 nsew signal input
rlabel metal3 s 37200 29928 37800 30048 6 chanx_left_in[16]
port 14 nsew signal input
rlabel metal3 s 200 28568 800 28688 6 chanx_left_in[17]
port 15 nsew signal input
rlabel metal3 s 37200 26528 37800 26648 6 chanx_left_in[18]
port 16 nsew signal input
rlabel metal2 s 8390 200 8446 800 6 chanx_left_in[1]
port 17 nsew signal input
rlabel metal2 s 35438 39200 35494 39800 6 chanx_left_in[2]
port 18 nsew signal input
rlabel metal3 s 200 30608 800 30728 6 chanx_left_in[3]
port 19 nsew signal input
rlabel metal3 s 200 14288 800 14408 6 chanx_left_in[4]
port 20 nsew signal input
rlabel metal2 s 25134 39200 25190 39800 6 chanx_left_in[5]
port 21 nsew signal input
rlabel metal2 s 34150 200 34206 800 6 chanx_left_in[6]
port 22 nsew signal input
rlabel metal2 s 35438 200 35494 800 6 chanx_left_in[7]
port 23 nsew signal input
rlabel metal2 s 23202 39200 23258 39800 6 chanx_left_in[8]
port 24 nsew signal input
rlabel metal3 s 37200 27888 37800 28008 6 chanx_left_in[9]
port 25 nsew signal input
rlabel metal2 s 5814 39200 5870 39800 6 chanx_left_out[0]
port 26 nsew signal output
rlabel metal3 s 200 23128 800 23248 6 chanx_left_out[10]
port 27 nsew signal output
rlabel metal3 s 37200 17008 37800 17128 6 chanx_left_out[11]
port 28 nsew signal output
rlabel metal2 s 19982 39200 20038 39800 6 chanx_left_out[12]
port 29 nsew signal output
rlabel metal3 s 37200 4768 37800 4888 6 chanx_left_out[13]
port 30 nsew signal output
rlabel metal2 s 26422 39200 26478 39800 6 chanx_left_out[14]
port 31 nsew signal output
rlabel metal3 s 200 3408 800 3528 6 chanx_left_out[15]
port 32 nsew signal output
rlabel metal3 s 200 10208 800 10328 6 chanx_left_out[16]
port 33 nsew signal output
rlabel metal3 s 200 1368 800 1488 6 chanx_left_out[17]
port 34 nsew signal output
rlabel metal2 s 18050 39200 18106 39800 6 chanx_left_out[18]
port 35 nsew signal output
rlabel metal3 s 37200 38768 37800 38888 6 chanx_left_out[1]
port 36 nsew signal output
rlabel metal3 s 200 21088 800 21208 6 chanx_left_out[2]
port 37 nsew signal output
rlabel metal3 s 37200 688 37800 808 6 chanx_left_out[3]
port 38 nsew signal output
rlabel metal3 s 37200 13608 37800 13728 6 chanx_left_out[4]
port 39 nsew signal output
rlabel metal3 s 200 39448 800 39568 6 chanx_left_out[5]
port 40 nsew signal output
rlabel metal2 s 30286 200 30342 800 6 chanx_left_out[6]
port 41 nsew signal output
rlabel metal2 s 14830 200 14886 800 6 chanx_left_out[7]
port 42 nsew signal output
rlabel metal3 s 200 6808 800 6928 6 chanx_left_out[8]
port 43 nsew signal output
rlabel metal3 s 37200 35368 37800 35488 6 chanx_left_out[9]
port 44 nsew signal output
rlabel metal3 s 200 8848 800 8968 6 chanx_right_in[0]
port 45 nsew signal input
rlabel metal2 s 3238 200 3294 800 6 chanx_right_in[10]
port 46 nsew signal input
rlabel metal2 s 9678 200 9734 800 6 chanx_right_in[11]
port 47 nsew signal input
rlabel metal2 s 32218 200 32274 800 6 chanx_right_in[12]
port 48 nsew signal input
rlabel metal3 s 37200 11568 37800 11688 6 chanx_right_in[13]
port 49 nsew signal input
rlabel metal3 s 37200 6128 37800 6248 6 chanx_right_in[14]
port 50 nsew signal input
rlabel metal2 s 23846 200 23902 800 6 chanx_right_in[15]
port 51 nsew signal input
rlabel metal3 s 200 37408 800 37528 6 chanx_right_in[16]
port 52 nsew signal input
rlabel metal2 s 37370 200 37426 800 6 chanx_right_in[17]
port 53 nsew signal input
rlabel metal2 s 9678 39200 9734 39800 6 chanx_right_in[18]
port 54 nsew signal input
rlabel metal3 s 37200 10208 37800 10328 6 chanx_right_in[1]
port 55 nsew signal input
rlabel metal3 s 200 25168 800 25288 6 chanx_right_in[2]
port 56 nsew signal input
rlabel metal2 s 28998 200 29054 800 6 chanx_right_in[3]
port 57 nsew signal input
rlabel metal3 s 200 17688 800 17808 6 chanx_right_in[4]
port 58 nsew signal input
rlabel metal3 s 200 31968 800 32088 6 chanx_right_in[5]
port 59 nsew signal input
rlabel metal2 s 12898 39200 12954 39800 6 chanx_right_in[6]
port 60 nsew signal input
rlabel metal2 s 18694 200 18750 800 6 chanx_right_in[7]
port 61 nsew signal input
rlabel metal2 s 18 200 74 800 6 chanx_right_in[8]
port 62 nsew signal input
rlabel metal2 s 21914 200 21970 800 6 chanx_right_in[9]
port 63 nsew signal input
rlabel metal2 s 10966 39200 11022 39800 6 chanx_right_out[0]
port 64 nsew signal output
rlabel metal2 s 21270 39200 21326 39800 6 chanx_right_out[10]
port 65 nsew signal output
rlabel metal2 s 33506 39200 33562 39800 6 chanx_right_out[11]
port 66 nsew signal output
rlabel metal3 s 200 26528 800 26648 6 chanx_right_out[12]
port 67 nsew signal output
rlabel metal2 s 4526 200 4582 800 6 chanx_right_out[13]
port 68 nsew signal output
rlabel metal2 s 1306 200 1362 800 6 chanx_right_out[14]
port 69 nsew signal output
rlabel metal2 s 36726 39200 36782 39800 6 chanx_right_out[15]
port 70 nsew signal output
rlabel metal2 s 28354 39200 28410 39800 6 chanx_right_out[16]
port 71 nsew signal output
rlabel metal2 s 16762 200 16818 800 6 chanx_right_out[17]
port 72 nsew signal output
rlabel metal3 s 37200 37408 37800 37528 6 chanx_right_out[18]
port 73 nsew signal output
rlabel metal3 s 37200 2728 37800 2848 6 chanx_right_out[1]
port 74 nsew signal output
rlabel metal2 s 4526 39200 4582 39800 6 chanx_right_out[2]
port 75 nsew signal output
rlabel metal3 s 37200 21088 37800 21208 6 chanx_right_out[3]
port 76 nsew signal output
rlabel metal2 s 6458 200 6514 800 6 chanx_right_out[4]
port 77 nsew signal output
rlabel metal2 s 11610 200 11666 800 6 chanx_right_out[5]
port 78 nsew signal output
rlabel metal3 s 200 15648 800 15768 6 chanx_right_out[6]
port 79 nsew signal output
rlabel metal3 s 37200 22448 37800 22568 6 chanx_right_out[7]
port 80 nsew signal output
rlabel metal2 s 19982 200 20038 800 6 chanx_right_out[8]
port 81 nsew signal output
rlabel metal2 s 31574 39200 31630 39800 6 chanx_right_out[9]
port 82 nsew signal output
rlabel metal2 s 30286 39200 30342 39800 6 pReset
port 83 nsew signal input
rlabel metal2 s 2594 39200 2650 39800 6 prog_clk
port 84 nsew signal input
rlabel metal2 s 7746 39200 7802 39800 6 top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_
port 85 nsew signal output
rlabel metal2 s 25134 200 25190 800 6 top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_
port 86 nsew signal output
rlabel metal3 s 200 12248 800 12368 6 top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_
port 87 nsew signal output
rlabel metal3 s 200 34008 800 34128 6 vccd1
port 88 nsew signal bidirectional
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 88 nsew signal bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 88 nsew signal bidirectional
rlabel metal3 s 37200 19048 37800 19168 6 vssd1
port 89 nsew signal bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 89 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 38000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1339430
string GDS_FILE /home/baungarten/Proyectos_caravel/FPGA_3/openlane/cbx_1__1_/runs/23_01_19_18_22/results/signoff/cbx_1__1_.magic.gds
string GDS_START 134360
<< end >>

