magic
tech sky130A
magscale 1 2
timestamp 1674174268
<< viali >>
rect 38301 37417 38335 37451
rect 16037 37349 16071 37383
rect 23397 37349 23431 37383
rect 5733 37281 5767 37315
rect 7113 37281 7147 37315
rect 8585 37281 8619 37315
rect 13185 37281 13219 37315
rect 20177 37281 20211 37315
rect 23949 37281 23983 37315
rect 29101 37281 29135 37315
rect 35081 37281 35115 37315
rect 35541 37281 35575 37315
rect 1685 37213 1719 37247
rect 6009 37213 6043 37247
rect 6837 37213 6871 37247
rect 9413 37213 9447 37247
rect 13461 37213 13495 37247
rect 14289 37213 14323 37247
rect 17141 37213 17175 37247
rect 17785 37213 17819 37247
rect 18429 37213 18463 37247
rect 19441 37213 19475 37247
rect 20913 37213 20947 37247
rect 21373 37213 21407 37247
rect 22017 37213 22051 37247
rect 22753 37213 22787 37247
rect 24593 37213 24627 37247
rect 25329 37213 25363 37247
rect 27169 37213 27203 37247
rect 29745 37213 29779 37247
rect 30665 37213 30699 37247
rect 31125 37213 31159 37247
rect 32321 37213 32355 37247
rect 33885 37213 33919 37247
rect 35817 37213 35851 37247
rect 37473 37213 37507 37247
rect 1961 37145 1995 37179
rect 9689 37145 9723 37179
rect 14565 37145 14599 37179
rect 3433 37077 3467 37111
rect 4261 37077 4295 37111
rect 11161 37077 11195 37111
rect 11713 37077 11747 37111
rect 16957 37077 16991 37111
rect 17693 37077 17727 37111
rect 18245 37077 18279 37111
rect 19625 37077 19659 37111
rect 20729 37077 20763 37111
rect 22201 37077 22235 37111
rect 22845 37077 22879 37111
rect 24777 37077 24811 37111
rect 25513 37077 25547 37111
rect 26525 37077 26559 37111
rect 27353 37077 27387 37111
rect 27997 37077 28031 37111
rect 28457 37077 28491 37111
rect 29929 37077 29963 37111
rect 30481 37077 30515 37111
rect 32505 37077 32539 37111
rect 33701 37077 33735 37111
rect 36829 37077 36863 37111
rect 37657 37077 37691 37111
rect 6009 36873 6043 36907
rect 16957 36873 16991 36907
rect 26065 36873 26099 36907
rect 3525 36805 3559 36839
rect 11989 36805 12023 36839
rect 22109 36805 22143 36839
rect 38209 36805 38243 36839
rect 3801 36737 3835 36771
rect 4261 36737 4295 36771
rect 17141 36737 17175 36771
rect 17601 36737 17635 36771
rect 18705 36737 18739 36771
rect 19625 36737 19659 36771
rect 20453 36737 20487 36771
rect 21373 36737 21407 36771
rect 21465 36737 21499 36771
rect 22201 36737 22235 36771
rect 22661 36737 22695 36771
rect 23949 36737 23983 36771
rect 25881 36737 25915 36771
rect 27353 36737 27387 36771
rect 27445 36737 27479 36771
rect 2053 36669 2087 36703
rect 4537 36669 4571 36703
rect 6837 36669 6871 36703
rect 7113 36669 7147 36703
rect 8861 36669 8895 36703
rect 9321 36669 9355 36703
rect 9597 36669 9631 36703
rect 11713 36669 11747 36703
rect 14013 36669 14047 36703
rect 19349 36669 19383 36703
rect 20177 36669 20211 36703
rect 23305 36669 23339 36703
rect 24041 36669 24075 36703
rect 26525 36669 26559 36703
rect 29653 36669 29687 36703
rect 17785 36601 17819 36635
rect 38025 36601 38059 36635
rect 11069 36533 11103 36567
rect 13461 36533 13495 36567
rect 14276 36533 14310 36567
rect 15761 36533 15795 36567
rect 16313 36533 16347 36567
rect 18613 36533 18647 36567
rect 22753 36533 22787 36567
rect 24685 36533 24719 36567
rect 25145 36533 25179 36567
rect 28089 36533 28123 36567
rect 28549 36533 28583 36567
rect 29101 36533 29135 36567
rect 37565 36533 37599 36567
rect 4077 36329 4111 36363
rect 6377 36329 6411 36363
rect 8585 36329 8619 36363
rect 17417 36329 17451 36363
rect 23857 36329 23891 36363
rect 37381 36329 37415 36363
rect 38209 36329 38243 36363
rect 3433 36261 3467 36295
rect 19533 36261 19567 36295
rect 26801 36261 26835 36295
rect 1961 36193 1995 36227
rect 4629 36193 4663 36227
rect 6837 36193 6871 36227
rect 9413 36193 9447 36227
rect 11621 36193 11655 36227
rect 13093 36193 13127 36227
rect 16037 36193 16071 36227
rect 18797 36193 18831 36227
rect 22109 36193 22143 36227
rect 22753 36193 22787 36227
rect 1685 36125 1719 36159
rect 3985 36125 4019 36159
rect 9137 36125 9171 36159
rect 11345 36125 11379 36159
rect 13737 36125 13771 36159
rect 16589 36125 16623 36159
rect 17233 36125 17267 36159
rect 17877 36125 17911 36159
rect 18889 36125 18923 36159
rect 19625 36125 19659 36159
rect 20085 36125 20119 36159
rect 21649 36125 21683 36159
rect 37565 36125 37599 36159
rect 38025 36125 38059 36159
rect 4905 36057 4939 36091
rect 7113 36057 7147 36091
rect 15761 36057 15795 36091
rect 20361 36057 20395 36091
rect 22661 36057 22695 36091
rect 10885 35989 10919 36023
rect 13553 35989 13587 36023
rect 14289 35989 14323 36023
rect 16681 35989 16715 36023
rect 17969 35989 18003 36023
rect 21557 35989 21591 36023
rect 23305 35989 23339 36023
rect 24685 35989 24719 36023
rect 25145 35989 25179 36023
rect 25697 35989 25731 36023
rect 26249 35989 26283 36023
rect 27353 35989 27387 36023
rect 27905 35989 27939 36023
rect 28457 35989 28491 36023
rect 29009 35989 29043 36023
rect 6929 35785 6963 35819
rect 10517 35785 10551 35819
rect 18797 35785 18831 35819
rect 5733 35717 5767 35751
rect 11989 35717 12023 35751
rect 15393 35717 15427 35751
rect 16221 35717 16255 35751
rect 19625 35717 19659 35751
rect 27169 35717 27203 35751
rect 2053 35649 2087 35683
rect 6009 35649 6043 35683
rect 7113 35649 7147 35683
rect 9597 35649 9631 35683
rect 10701 35649 10735 35683
rect 16313 35649 16347 35683
rect 17049 35649 17083 35683
rect 17969 35649 18003 35683
rect 18613 35649 18647 35683
rect 19717 35649 19751 35683
rect 20361 35649 20395 35683
rect 21005 35649 21039 35683
rect 22201 35649 22235 35683
rect 38025 35649 38059 35683
rect 2329 35581 2363 35615
rect 7573 35581 7607 35615
rect 9321 35581 9355 35615
rect 11713 35581 11747 35615
rect 13921 35581 13955 35615
rect 15669 35581 15703 35615
rect 20913 35581 20947 35615
rect 23213 35581 23247 35615
rect 3801 35513 3835 35547
rect 27721 35513 27755 35547
rect 28273 35513 28307 35547
rect 28825 35513 28859 35547
rect 4261 35445 4295 35479
rect 13461 35445 13495 35479
rect 16957 35445 16991 35479
rect 18061 35445 18095 35479
rect 20269 35445 20303 35479
rect 22109 35445 22143 35479
rect 22753 35445 22787 35479
rect 23765 35445 23799 35479
rect 24317 35445 24351 35479
rect 24869 35445 24903 35479
rect 25421 35445 25455 35479
rect 25973 35445 26007 35479
rect 26525 35445 26559 35479
rect 37473 35445 37507 35479
rect 38209 35445 38243 35479
rect 6837 35241 6871 35275
rect 24593 35241 24627 35275
rect 25697 35241 25731 35275
rect 26249 35241 26283 35275
rect 26801 35241 26835 35275
rect 27353 35241 27387 35275
rect 27905 35241 27939 35275
rect 18797 35173 18831 35207
rect 22937 35173 22971 35207
rect 3433 35105 3467 35139
rect 4629 35105 4663 35139
rect 10701 35105 10735 35139
rect 20085 35105 20119 35139
rect 21005 35105 21039 35139
rect 25145 35105 25179 35139
rect 3985 35037 4019 35071
rect 8585 35037 8619 35071
rect 9137 35037 9171 35071
rect 9413 35037 9447 35071
rect 13277 35037 13311 35071
rect 15025 35037 15059 35071
rect 15485 35037 15519 35071
rect 16313 35037 16347 35071
rect 17233 35037 17267 35071
rect 17325 35037 17359 35071
rect 17877 35037 17911 35071
rect 17969 35037 18003 35071
rect 18889 35037 18923 35071
rect 19901 35037 19935 35071
rect 20821 35037 20855 35071
rect 3157 34969 3191 35003
rect 4905 34969 4939 35003
rect 8309 34969 8343 35003
rect 10977 34969 11011 35003
rect 16221 34969 16255 35003
rect 1685 34901 1719 34935
rect 4077 34901 4111 34935
rect 6377 34901 6411 34935
rect 12449 34901 12483 34935
rect 13093 34901 13127 34935
rect 14289 34901 14323 34935
rect 14933 34901 14967 34935
rect 15577 34901 15611 34935
rect 21741 34901 21775 34935
rect 22385 34901 22419 34935
rect 23489 34901 23523 34935
rect 24041 34901 24075 34935
rect 10425 34697 10459 34731
rect 11069 34697 11103 34731
rect 18245 34697 18279 34731
rect 21373 34697 21407 34731
rect 25329 34697 25363 34731
rect 26525 34697 26559 34731
rect 9781 34629 9815 34663
rect 17417 34629 17451 34663
rect 17509 34629 17543 34663
rect 22569 34629 22603 34663
rect 23213 34629 23247 34663
rect 2605 34561 2639 34595
rect 5549 34561 5583 34595
rect 6561 34561 6595 34595
rect 9873 34561 9907 34595
rect 10517 34561 10551 34595
rect 11161 34561 11195 34595
rect 13461 34561 13495 34595
rect 13921 34561 13955 34595
rect 14841 34561 14875 34595
rect 15577 34561 15611 34595
rect 16865 34561 16899 34595
rect 18337 34561 18371 34595
rect 18981 34561 19015 34595
rect 19901 34561 19935 34595
rect 22017 34561 22051 34595
rect 2881 34493 2915 34527
rect 3801 34493 3835 34527
rect 6653 34493 6687 34527
rect 7205 34493 7239 34527
rect 8953 34493 8987 34527
rect 9229 34493 9263 34527
rect 13185 34493 13219 34527
rect 14749 34493 14783 34527
rect 15485 34493 15519 34527
rect 16037 34493 16071 34527
rect 18889 34493 18923 34527
rect 20177 34493 20211 34527
rect 24317 34493 24351 34527
rect 24777 34425 24811 34459
rect 25881 34425 25915 34459
rect 27169 34425 27203 34459
rect 5285 34357 5319 34391
rect 11713 34357 11747 34391
rect 14105 34357 14139 34391
rect 20821 34357 20855 34391
rect 23673 34357 23707 34391
rect 1948 34153 1982 34187
rect 4813 34153 4847 34187
rect 9229 34153 9263 34187
rect 9781 34153 9815 34187
rect 23213 34153 23247 34187
rect 25697 34153 25731 34187
rect 26249 34153 26283 34187
rect 21465 34085 21499 34119
rect 1685 34017 1719 34051
rect 5365 34017 5399 34051
rect 7389 34017 7423 34051
rect 12173 34017 12207 34051
rect 19533 34017 19567 34051
rect 20177 34017 20211 34051
rect 3985 33949 4019 33983
rect 4629 33949 4663 33983
rect 7849 33949 7883 33983
rect 9321 33949 9355 33983
rect 13093 33949 13127 33983
rect 14841 33949 14875 33983
rect 17049 33949 17083 33983
rect 19993 33949 20027 33983
rect 24593 33949 24627 33983
rect 7113 33881 7147 33915
rect 11897 33881 11931 33915
rect 14749 33881 14783 33915
rect 15393 33881 15427 33915
rect 15485 33881 15519 33915
rect 16037 33881 16071 33915
rect 16497 33881 16531 33915
rect 17141 33881 17175 33915
rect 18153 33881 18187 33915
rect 18245 33881 18279 33915
rect 18797 33881 18831 33915
rect 25145 33881 25179 33915
rect 3433 33813 3467 33847
rect 4077 33813 4111 33847
rect 7941 33813 7975 33847
rect 8585 33813 8619 33847
rect 10425 33813 10459 33847
rect 13185 33813 13219 33847
rect 20913 33813 20947 33847
rect 22109 33813 22143 33847
rect 22569 33813 22603 33847
rect 23673 33813 23707 33847
rect 3065 33609 3099 33643
rect 19533 33609 19567 33643
rect 22661 33609 22695 33643
rect 25329 33609 25363 33643
rect 5273 33541 5307 33575
rect 7297 33541 7331 33575
rect 16037 33541 16071 33575
rect 16129 33541 16163 33575
rect 21097 33541 21131 33575
rect 2421 33473 2455 33507
rect 2973 33473 3007 33507
rect 5549 33473 5583 33507
rect 7021 33473 7055 33507
rect 9321 33473 9355 33507
rect 11713 33473 11747 33507
rect 14657 33473 14691 33507
rect 16865 33473 16899 33507
rect 17969 33473 18003 33507
rect 18981 33473 19015 33507
rect 19625 33473 19659 33507
rect 20637 33473 20671 33507
rect 24869 33473 24903 33507
rect 26433 33473 26467 33507
rect 37565 33473 37599 33507
rect 38209 33473 38243 33507
rect 2145 33405 2179 33439
rect 9597 33405 9631 33439
rect 11989 33405 12023 33439
rect 13737 33405 13771 33439
rect 15853 33405 15887 33439
rect 18889 33405 18923 33439
rect 23673 33405 23707 33439
rect 20545 33337 20579 33371
rect 23121 33337 23155 33371
rect 25881 33337 25915 33371
rect 38025 33337 38059 33371
rect 3801 33269 3835 33303
rect 8769 33269 8803 33303
rect 11069 33269 11103 33303
rect 14565 33269 14599 33303
rect 16957 33269 16991 33303
rect 18061 33269 18095 33303
rect 22109 33269 22143 33303
rect 24225 33269 24259 33303
rect 1948 33065 1982 33099
rect 3433 33065 3467 33099
rect 19533 33065 19567 33099
rect 20729 33065 20763 33099
rect 21741 33065 21775 33099
rect 22937 33065 22971 33099
rect 23489 33065 23523 33099
rect 25237 33065 25271 33099
rect 1685 32929 1719 32963
rect 4905 32929 4939 32963
rect 6929 32929 6963 32963
rect 11253 32929 11287 32963
rect 11529 32929 11563 32963
rect 15577 32929 15611 32963
rect 16589 32929 16623 32963
rect 16957 32929 16991 32963
rect 4261 32861 4295 32895
rect 7757 32861 7791 32895
rect 8585 32861 8619 32895
rect 9137 32861 9171 32895
rect 9873 32861 9907 32895
rect 10609 32861 10643 32895
rect 14381 32861 14415 32895
rect 18337 32861 18371 32895
rect 19625 32861 19659 32895
rect 21833 32861 21867 32895
rect 25697 32861 25731 32895
rect 6653 32793 6687 32827
rect 9965 32793 9999 32827
rect 13277 32793 13311 32827
rect 14933 32793 14967 32827
rect 15025 32793 15059 32827
rect 16681 32793 16715 32827
rect 4353 32725 4387 32759
rect 7665 32725 7699 32759
rect 8493 32725 8527 32759
rect 9229 32725 9263 32759
rect 10701 32725 10735 32759
rect 18429 32725 18463 32759
rect 20177 32725 20211 32759
rect 22293 32725 22327 32759
rect 24041 32725 24075 32759
rect 24593 32725 24627 32759
rect 1777 32521 1811 32555
rect 3065 32521 3099 32555
rect 5917 32521 5951 32555
rect 11805 32521 11839 32555
rect 20177 32521 20211 32555
rect 22109 32521 22143 32555
rect 8493 32453 8527 32487
rect 9689 32453 9723 32487
rect 17417 32453 17451 32487
rect 18337 32453 18371 32487
rect 18429 32453 18463 32487
rect 18981 32453 19015 32487
rect 1685 32385 1719 32419
rect 2605 32385 2639 32419
rect 5457 32385 5491 32419
rect 19625 32385 19659 32419
rect 20269 32385 20303 32419
rect 22201 32385 22235 32419
rect 38025 32385 38059 32419
rect 5181 32317 5215 32351
rect 6745 32317 6779 32351
rect 8769 32317 8803 32351
rect 9413 32317 9447 32351
rect 13277 32317 13311 32351
rect 13553 32317 13587 32351
rect 15577 32317 15611 32351
rect 15853 32317 15887 32351
rect 17509 32317 17543 32351
rect 19533 32317 19567 32351
rect 20729 32317 20763 32351
rect 22661 32317 22695 32351
rect 23765 32317 23799 32351
rect 24317 32317 24351 32351
rect 2421 32249 2455 32283
rect 3709 32249 3743 32283
rect 11161 32249 11195 32283
rect 16957 32249 16991 32283
rect 14105 32181 14139 32215
rect 21373 32181 21407 32215
rect 23213 32181 23247 32215
rect 38209 32181 38243 32215
rect 1685 31977 1719 32011
rect 4813 31977 4847 32011
rect 13001 31977 13035 32011
rect 19533 31977 19567 32011
rect 21741 31977 21775 32011
rect 22293 31977 22327 32011
rect 23397 31977 23431 32011
rect 9505 31909 9539 31943
rect 16405 31909 16439 31943
rect 22845 31909 22879 31943
rect 3157 31841 3191 31875
rect 7389 31841 7423 31875
rect 7849 31841 7883 31875
rect 10793 31841 10827 31875
rect 12541 31841 12575 31875
rect 14381 31841 14415 31875
rect 15393 31841 15427 31875
rect 15761 31841 15795 31875
rect 21189 31841 21223 31875
rect 3433 31773 3467 31807
rect 4261 31773 4295 31807
rect 4721 31773 4755 31807
rect 8401 31773 8435 31807
rect 8493 31773 8527 31807
rect 9413 31773 9447 31807
rect 10057 31773 10091 31807
rect 10149 31773 10183 31807
rect 13645 31773 13679 31807
rect 13737 31773 13771 31807
rect 14289 31773 14323 31807
rect 18797 31773 18831 31807
rect 18889 31773 18923 31807
rect 19625 31773 19659 31807
rect 20269 31773 20303 31807
rect 21281 31773 21315 31807
rect 5365 31705 5399 31739
rect 7113 31705 7147 31739
rect 12265 31705 12299 31739
rect 15669 31705 15703 31739
rect 16865 31705 16899 31739
rect 16957 31705 16991 31739
rect 17601 31705 17635 31739
rect 17693 31705 17727 31739
rect 18245 31705 18279 31739
rect 20177 31705 20211 31739
rect 4169 31637 4203 31671
rect 5917 31433 5951 31467
rect 20913 31433 20947 31467
rect 22109 31433 22143 31467
rect 22569 31433 22603 31467
rect 23213 31433 23247 31467
rect 3249 31365 3283 31399
rect 15025 31365 15059 31399
rect 17325 31365 17359 31399
rect 17877 31365 17911 31399
rect 18521 31365 18555 31399
rect 19073 31365 19107 31399
rect 1685 31297 1719 31331
rect 2513 31297 2547 31331
rect 5825 31297 5859 31331
rect 6745 31297 6779 31331
rect 9413 31297 9447 31331
rect 10333 31297 10367 31331
rect 10977 31297 11011 31331
rect 14197 31297 14231 31331
rect 16037 31297 16071 31331
rect 19717 31297 19751 31331
rect 20361 31297 20395 31331
rect 20821 31297 20855 31331
rect 2973 31229 3007 31263
rect 4997 31229 5031 31263
rect 7389 31229 7423 31263
rect 9137 31229 9171 31263
rect 13277 31229 13311 31263
rect 13553 31229 13587 31263
rect 14933 31229 14967 31263
rect 15209 31229 15243 31263
rect 17233 31229 17267 31263
rect 18429 31229 18463 31263
rect 1869 31161 1903 31195
rect 20269 31161 20303 31195
rect 2329 31093 2363 31127
rect 6837 31093 6871 31127
rect 10425 31093 10459 31127
rect 11069 31093 11103 31127
rect 11805 31093 11839 31127
rect 14289 31093 14323 31127
rect 16129 31093 16163 31127
rect 19625 31093 19659 31127
rect 9229 30889 9263 30923
rect 10425 30889 10459 30923
rect 20177 30889 20211 30923
rect 20729 30889 20763 30923
rect 16221 30821 16255 30855
rect 19533 30821 19567 30855
rect 21741 30821 21775 30855
rect 31125 30821 31159 30855
rect 4261 30753 4295 30787
rect 8585 30753 8619 30787
rect 15025 30753 15059 30787
rect 3433 30685 3467 30719
rect 3985 30685 4019 30719
rect 6009 30685 6043 30719
rect 9689 30685 9723 30719
rect 10333 30685 10367 30719
rect 10977 30685 11011 30719
rect 13001 30685 13035 30719
rect 13553 30685 13587 30719
rect 14289 30685 14323 30719
rect 18613 30685 18647 30719
rect 19441 30685 19475 30719
rect 20269 30685 20303 30719
rect 21833 30685 21867 30719
rect 22477 30685 22511 30719
rect 30941 30685 30975 30719
rect 31585 30685 31619 30719
rect 3157 30617 3191 30651
rect 6561 30617 6595 30651
rect 8309 30617 8343 30651
rect 9781 30617 9815 30651
rect 12725 30617 12759 30651
rect 15117 30617 15151 30651
rect 15669 30617 15703 30651
rect 16681 30617 16715 30651
rect 16773 30617 16807 30651
rect 17325 30617 17359 30651
rect 17877 30617 17911 30651
rect 17969 30617 18003 30651
rect 18521 30617 18555 30651
rect 1685 30549 1719 30583
rect 13645 30549 13679 30583
rect 14381 30549 14415 30583
rect 22385 30549 22419 30583
rect 9413 30345 9447 30379
rect 3157 30277 3191 30311
rect 5365 30277 5399 30311
rect 14933 30277 14967 30311
rect 16129 30277 16163 30311
rect 17049 30277 17083 30311
rect 18061 30209 18095 30243
rect 18981 30209 19015 30243
rect 19625 30209 19659 30243
rect 20269 30209 20303 30243
rect 29561 30209 29595 30243
rect 38025 30209 38059 30243
rect 3433 30141 3467 30175
rect 5641 30141 5675 30175
rect 7021 30141 7055 30175
rect 7297 30141 7331 30175
rect 10885 30141 10919 30175
rect 11161 30141 11195 30175
rect 11713 30141 11747 30175
rect 13185 30141 13219 30175
rect 13461 30141 13495 30175
rect 14381 30141 14415 30175
rect 15025 30141 15059 30175
rect 15945 30141 15979 30175
rect 16221 30141 16255 30175
rect 16957 30141 16991 30175
rect 17417 30141 17451 30175
rect 22109 30141 22143 30175
rect 30113 30141 30147 30175
rect 1685 30073 1719 30107
rect 20177 30073 20211 30107
rect 20821 30073 20855 30107
rect 22569 30073 22603 30107
rect 3893 30005 3927 30039
rect 8769 30005 8803 30039
rect 18153 30005 18187 30039
rect 18889 30005 18923 30039
rect 19533 30005 19567 30039
rect 21281 30005 21315 30039
rect 29469 30005 29503 30039
rect 38209 30005 38243 30039
rect 1948 29801 1982 29835
rect 3985 29801 4019 29835
rect 20177 29801 20211 29835
rect 20821 29801 20855 29835
rect 21465 29801 21499 29835
rect 22569 29801 22603 29835
rect 38025 29801 38059 29835
rect 9781 29733 9815 29767
rect 1685 29665 1719 29699
rect 8493 29665 8527 29699
rect 10609 29665 10643 29699
rect 10885 29665 10919 29699
rect 13645 29665 13679 29699
rect 14565 29665 14599 29699
rect 15577 29665 15611 29699
rect 5733 29597 5767 29631
rect 17141 29597 17175 29631
rect 19441 29597 19475 29631
rect 20269 29597 20303 29631
rect 20729 29597 20763 29631
rect 37841 29597 37875 29631
rect 5457 29529 5491 29563
rect 8217 29529 8251 29563
rect 9229 29529 9263 29563
rect 9321 29529 9355 29563
rect 13001 29529 13035 29563
rect 13093 29529 13127 29563
rect 14657 29529 14691 29563
rect 16497 29529 16531 29563
rect 16589 29529 16623 29563
rect 18153 29529 18187 29563
rect 18245 29529 18279 29563
rect 18797 29529 18831 29563
rect 21925 29529 21959 29563
rect 3433 29461 3467 29495
rect 6745 29461 6779 29495
rect 12357 29461 12391 29495
rect 19533 29461 19567 29495
rect 37381 29461 37415 29495
rect 2697 29257 2731 29291
rect 5917 29257 5951 29291
rect 19625 29257 19659 29291
rect 1685 29189 1719 29223
rect 8217 29189 8251 29223
rect 8769 29189 8803 29223
rect 9413 29189 9447 29223
rect 10609 29189 10643 29223
rect 11989 29189 12023 29223
rect 14197 29189 14231 29223
rect 15393 29189 15427 29223
rect 15945 29189 15979 29223
rect 17509 29189 17543 29223
rect 17601 29189 17635 29223
rect 18337 29189 18371 29223
rect 2605 29121 2639 29155
rect 5825 29121 5859 29155
rect 7113 29121 7147 29155
rect 11161 29121 11195 29155
rect 11713 29121 11747 29155
rect 19441 29121 19475 29155
rect 20269 29121 20303 29155
rect 20913 29121 20947 29155
rect 21373 29121 21407 29155
rect 38025 29121 38059 29155
rect 3249 29053 3283 29087
rect 4997 29053 5031 29087
rect 6929 29053 6963 29087
rect 8125 29053 8159 29087
rect 9321 29053 9355 29087
rect 10517 29053 10551 29087
rect 14106 29053 14140 29087
rect 15301 29053 15335 29087
rect 17325 29053 17359 29087
rect 18245 29053 18279 29087
rect 18521 29053 18555 29087
rect 22017 29053 22051 29087
rect 1869 28985 1903 29019
rect 9873 28985 9907 29019
rect 13461 28985 13495 29019
rect 14657 28985 14691 29019
rect 20821 28985 20855 29019
rect 38209 28985 38243 29019
rect 4739 28917 4773 28951
rect 7573 28917 7607 28951
rect 20177 28917 20211 28951
rect 2697 28713 2731 28747
rect 33977 28713 34011 28747
rect 3341 28645 3375 28679
rect 9965 28645 9999 28679
rect 20821 28645 20855 28679
rect 30941 28645 30975 28679
rect 2053 28577 2087 28611
rect 6561 28577 6595 28611
rect 7941 28577 7975 28611
rect 10517 28577 10551 28611
rect 13461 28577 13495 28611
rect 14933 28577 14967 28611
rect 16037 28577 16071 28611
rect 16313 28577 16347 28611
rect 16957 28577 16991 28611
rect 2145 28509 2179 28543
rect 2605 28509 2639 28543
rect 3433 28509 3467 28543
rect 7389 28509 7423 28543
rect 20913 28509 20947 28543
rect 21373 28509 21407 28543
rect 30757 28509 30791 28543
rect 31401 28509 31435 28543
rect 34161 28509 34195 28543
rect 34897 28509 34931 28543
rect 4077 28441 4111 28475
rect 4169 28441 4203 28475
rect 4721 28441 4755 28475
rect 5549 28441 5583 28475
rect 5641 28441 5675 28475
rect 8033 28441 8067 28475
rect 8585 28441 8619 28475
rect 9413 28441 9447 28475
rect 9505 28441 9539 28475
rect 11437 28441 11471 28475
rect 11529 28441 11563 28475
rect 12541 28441 12575 28475
rect 12633 28441 12667 28475
rect 14289 28441 14323 28475
rect 14841 28441 14875 28475
rect 16221 28441 16255 28475
rect 17049 28441 17083 28475
rect 17601 28441 17635 28475
rect 18153 28441 18187 28475
rect 18705 28441 18739 28475
rect 18797 28441 18831 28475
rect 7297 28373 7331 28407
rect 19625 28373 19659 28407
rect 20085 28373 20119 28407
rect 2697 28169 2731 28203
rect 4537 28169 4571 28203
rect 5273 28169 5307 28203
rect 16221 28169 16255 28203
rect 18245 28169 18279 28203
rect 21097 28169 21131 28203
rect 7757 28101 7791 28135
rect 9413 28101 9447 28135
rect 10609 28101 10643 28135
rect 12909 28101 12943 28135
rect 13461 28101 13495 28135
rect 14289 28101 14323 28135
rect 17049 28101 17083 28135
rect 18981 28101 19015 28135
rect 22109 28101 22143 28135
rect 1869 28033 1903 28067
rect 2513 28033 2547 28067
rect 3341 28033 3375 28067
rect 3985 28033 4019 28067
rect 4537 28033 4571 28067
rect 5181 28033 5215 28067
rect 5825 28033 5859 28067
rect 5917 28033 5951 28067
rect 6929 28033 6963 28067
rect 9965 28033 9999 28067
rect 12265 28033 12299 28067
rect 15485 28033 15519 28067
rect 16129 28033 16163 28067
rect 18337 28033 18371 28067
rect 19993 28033 20027 28067
rect 3249 27965 3283 27999
rect 7665 27965 7699 27999
rect 8309 27965 8343 27999
rect 9321 27965 9355 27999
rect 10517 27965 10551 27999
rect 12817 27965 12851 27999
rect 14197 27965 14231 27999
rect 14657 27965 14691 27999
rect 16957 27965 16991 27999
rect 17233 27965 17267 27999
rect 18889 27965 18923 27999
rect 20177 27965 20211 27999
rect 1685 27897 1719 27931
rect 3893 27897 3927 27931
rect 11069 27897 11103 27931
rect 19441 27897 19475 27931
rect 7021 27829 7055 27863
rect 12173 27829 12207 27863
rect 15393 27829 15427 27863
rect 20361 27829 20395 27863
rect 8493 27625 8527 27659
rect 18889 27625 18923 27659
rect 22385 27625 22419 27659
rect 22845 27625 22879 27659
rect 1961 27557 1995 27591
rect 2697 27557 2731 27591
rect 14657 27557 14691 27591
rect 3341 27489 3375 27523
rect 5365 27489 5399 27523
rect 6561 27489 6595 27523
rect 12081 27489 12115 27523
rect 15209 27489 15243 27523
rect 15853 27489 15887 27523
rect 17693 27489 17727 27523
rect 18429 27489 18463 27523
rect 19993 27489 20027 27523
rect 20453 27489 20487 27523
rect 24685 27489 24719 27523
rect 1869 27421 1903 27455
rect 2789 27421 2823 27455
rect 3249 27421 3283 27455
rect 4537 27421 4571 27455
rect 6009 27421 6043 27455
rect 6469 27421 6503 27455
rect 7113 27421 7147 27455
rect 7749 27421 7783 27455
rect 8401 27421 8435 27455
rect 9137 27421 9171 27455
rect 9321 27421 9355 27455
rect 13737 27421 13771 27455
rect 17601 27421 17635 27455
rect 18245 27421 18279 27455
rect 21281 27421 21315 27455
rect 21741 27421 21775 27455
rect 24777 27421 24811 27455
rect 4629 27353 4663 27387
rect 7849 27353 7883 27387
rect 10241 27353 10275 27387
rect 11161 27353 11195 27387
rect 11253 27353 11287 27387
rect 12173 27353 12207 27387
rect 13093 27353 13127 27387
rect 15117 27353 15151 27387
rect 15945 27353 15979 27387
rect 16865 27353 16899 27387
rect 20085 27353 20119 27387
rect 25329 27353 25363 27387
rect 3985 27285 4019 27319
rect 5917 27285 5951 27319
rect 7205 27285 7239 27319
rect 9781 27285 9815 27319
rect 13553 27285 13587 27319
rect 21189 27285 21223 27319
rect 2421 27081 2455 27115
rect 3065 27081 3099 27115
rect 16221 27081 16255 27115
rect 20361 27081 20395 27115
rect 22109 27081 22143 27115
rect 23765 27081 23799 27115
rect 3985 27013 4019 27047
rect 8033 27013 8067 27047
rect 8125 27013 8159 27047
rect 9229 27013 9263 27047
rect 10425 27013 10459 27047
rect 10977 27013 11011 27047
rect 11897 27013 11931 27047
rect 12817 27013 12851 27047
rect 14381 27013 14415 27047
rect 14933 27013 14967 27047
rect 16957 27013 16991 27047
rect 17049 27013 17083 27047
rect 18337 27013 18371 27047
rect 19441 27013 19475 27047
rect 22569 27013 22603 27047
rect 38025 27013 38059 27047
rect 1869 26945 1903 26979
rect 2513 26945 2547 26979
rect 2973 26945 3007 26979
rect 3893 26945 3927 26979
rect 4537 26945 4571 26979
rect 5181 26945 5215 26979
rect 5833 26951 5867 26985
rect 6837 26945 6871 26979
rect 7481 26945 7515 26979
rect 13737 26945 13771 26979
rect 15577 26945 15611 26979
rect 16129 26945 16163 26979
rect 18245 26945 18279 26979
rect 20453 26945 20487 26979
rect 20913 26945 20947 26979
rect 23581 26945 23615 26979
rect 24225 26945 24259 26979
rect 37565 26945 37599 26979
rect 38209 26945 38243 26979
rect 4629 26877 4663 26911
rect 9137 26877 9171 26911
rect 10333 26877 10367 26911
rect 11805 26877 11839 26911
rect 14289 26877 14323 26911
rect 18889 26877 18923 26911
rect 19533 26877 19567 26911
rect 5917 26809 5951 26843
rect 9689 26809 9723 26843
rect 17509 26809 17543 26843
rect 1685 26741 1719 26775
rect 5273 26741 5307 26775
rect 6929 26741 6963 26775
rect 13645 26741 13679 26775
rect 15485 26741 15519 26775
rect 1961 26537 1995 26571
rect 9505 26537 9539 26571
rect 15117 26537 15151 26571
rect 17141 26537 17175 26571
rect 18889 26537 18923 26571
rect 19533 26537 19567 26571
rect 20821 26537 20855 26571
rect 2605 26469 2639 26503
rect 7297 26469 7331 26503
rect 11253 26469 11287 26503
rect 12081 26469 12115 26503
rect 4721 26401 4755 26435
rect 10149 26401 10183 26435
rect 10793 26401 10827 26435
rect 13737 26401 13771 26435
rect 15301 26401 15335 26435
rect 15485 26401 15519 26435
rect 18245 26401 18279 26435
rect 19993 26401 20027 26435
rect 21925 26401 21959 26435
rect 30481 26401 30515 26435
rect 1869 26333 1903 26367
rect 2513 26333 2547 26367
rect 3249 26333 3283 26367
rect 3985 26333 4019 26367
rect 4077 26333 4111 26367
rect 4629 26333 4663 26367
rect 5273 26333 5307 26367
rect 5917 26333 5951 26367
rect 6653 26333 6687 26367
rect 6745 26333 6779 26367
rect 7205 26333 7239 26367
rect 9965 26333 9999 26367
rect 10609 26333 10643 26367
rect 11713 26333 11747 26367
rect 11897 26333 11931 26367
rect 14381 26333 14415 26367
rect 16129 26333 16163 26367
rect 16957 26333 16991 26367
rect 17601 26333 17635 26367
rect 18429 26333 18463 26367
rect 20177 26333 20211 26367
rect 21373 26333 21407 26367
rect 29837 26333 29871 26367
rect 29929 26333 29963 26367
rect 30573 26333 30607 26367
rect 31125 26333 31159 26367
rect 3341 26265 3375 26299
rect 5365 26265 5399 26299
rect 6009 26265 6043 26299
rect 7941 26265 7975 26299
rect 8033 26265 8067 26299
rect 8585 26265 8619 26299
rect 13093 26265 13127 26299
rect 13185 26265 13219 26299
rect 16037 26265 16071 26299
rect 17693 26265 17727 26299
rect 38209 26197 38243 26231
rect 1961 25993 1995 26027
rect 4077 25993 4111 26027
rect 4629 25993 4663 26027
rect 6745 25993 6779 26027
rect 13737 25993 13771 26027
rect 17233 25993 17267 26027
rect 19165 25993 19199 26027
rect 21097 25993 21131 26027
rect 37841 25993 37875 26027
rect 3249 25925 3283 25959
rect 7481 25925 7515 25959
rect 9045 25925 9079 25959
rect 9873 25925 9907 25959
rect 13093 25925 13127 25959
rect 13185 25925 13219 25959
rect 22569 25925 22603 25959
rect 1869 25857 1903 25891
rect 2513 25857 2547 25891
rect 3157 25857 3191 25891
rect 3985 25857 4019 25891
rect 5181 25857 5215 25891
rect 5825 25857 5859 25891
rect 6653 25857 6687 25891
rect 10977 25857 11011 25891
rect 11897 25857 11931 25891
rect 14381 25857 14415 25891
rect 15025 25857 15059 25891
rect 15669 25857 15703 25891
rect 16313 25857 16347 25891
rect 17141 25857 17175 25891
rect 17969 25857 18003 25891
rect 19257 25857 19291 25891
rect 21189 25857 21223 25891
rect 38025 25857 38059 25891
rect 7389 25789 7423 25823
rect 8493 25789 8527 25823
rect 9137 25789 9171 25823
rect 9781 25789 9815 25823
rect 14197 25789 14231 25823
rect 17785 25789 17819 25823
rect 19901 25789 19935 25823
rect 20085 25789 20119 25823
rect 2605 25721 2639 25755
rect 5273 25721 5307 25755
rect 7941 25721 7975 25755
rect 10333 25721 10367 25755
rect 12633 25721 12667 25755
rect 16221 25721 16255 25755
rect 18429 25721 18463 25755
rect 20269 25721 20303 25755
rect 5917 25653 5951 25687
rect 11069 25653 11103 25687
rect 11989 25653 12023 25687
rect 14933 25653 14967 25687
rect 15577 25653 15611 25687
rect 22017 25653 22051 25687
rect 2605 25449 2639 25483
rect 3249 25449 3283 25483
rect 4077 25449 4111 25483
rect 6193 25449 6227 25483
rect 7941 25449 7975 25483
rect 13737 25449 13771 25483
rect 17509 25449 17543 25483
rect 21097 25449 21131 25483
rect 1961 25381 1995 25415
rect 4905 25381 4939 25415
rect 14933 25381 14967 25415
rect 18797 25381 18831 25415
rect 20453 25381 20487 25415
rect 5641 25313 5675 25347
rect 7573 25313 7607 25347
rect 8585 25313 8619 25347
rect 9965 25313 9999 25347
rect 11345 25313 11379 25347
rect 12449 25313 12483 25347
rect 14381 25313 14415 25347
rect 16221 25313 16255 25347
rect 18245 25313 18279 25347
rect 1869 25245 1903 25279
rect 2513 25245 2547 25279
rect 3157 25245 3191 25279
rect 4169 25245 4203 25279
rect 4813 25245 4847 25279
rect 6101 25245 6135 25279
rect 6745 25245 6779 25279
rect 7389 25245 7423 25279
rect 11529 25245 11563 25279
rect 16405 25245 16439 25279
rect 17049 25245 17083 25279
rect 17693 25245 17727 25279
rect 21189 25245 21223 25279
rect 21649 25245 21683 25279
rect 28365 25245 28399 25279
rect 29745 25245 29779 25279
rect 37841 25245 37875 25279
rect 6837 25177 6871 25211
rect 9689 25177 9723 25211
rect 9781 25177 9815 25211
rect 13001 25177 13035 25211
rect 13093 25177 13127 25211
rect 14473 25177 14507 25211
rect 18337 25177 18371 25211
rect 19901 25177 19935 25211
rect 19993 25177 20027 25211
rect 28457 25177 28491 25211
rect 10793 25109 10827 25143
rect 11989 25109 12023 25143
rect 15761 25109 15795 25143
rect 16957 25109 16991 25143
rect 29837 25109 29871 25143
rect 38025 25109 38059 25143
rect 7941 24905 7975 24939
rect 10609 24837 10643 24871
rect 12357 24837 12391 24871
rect 15761 24837 15795 24871
rect 19809 24837 19843 24871
rect 1869 24769 1903 24803
rect 2329 24769 2363 24803
rect 2973 24769 3007 24803
rect 3709 24769 3743 24803
rect 3801 24769 3835 24803
rect 4813 24769 4847 24803
rect 5825 24769 5859 24803
rect 5917 24769 5951 24803
rect 6745 24769 6779 24803
rect 7849 24769 7883 24803
rect 8493 24769 8527 24803
rect 8585 24769 8619 24803
rect 9781 24769 9815 24803
rect 12909 24769 12943 24803
rect 13461 24769 13495 24803
rect 14565 24769 14599 24803
rect 14749 24769 14783 24803
rect 17969 24769 18003 24803
rect 18613 24769 18647 24803
rect 18705 24769 18739 24803
rect 38025 24769 38059 24803
rect 3065 24701 3099 24735
rect 7389 24701 7423 24735
rect 9137 24701 9171 24735
rect 9321 24701 9355 24735
rect 10517 24701 10551 24735
rect 12265 24701 12299 24735
rect 15669 24701 15703 24735
rect 16865 24701 16899 24735
rect 19901 24701 19935 24735
rect 20453 24701 20487 24735
rect 11069 24633 11103 24667
rect 14381 24633 14415 24667
rect 16221 24633 16255 24667
rect 19349 24633 19383 24667
rect 1685 24565 1719 24599
rect 2421 24565 2455 24599
rect 5365 24565 5399 24599
rect 6653 24565 6687 24599
rect 13553 24565 13587 24599
rect 18061 24565 18095 24599
rect 38209 24565 38243 24599
rect 1961 24361 1995 24395
rect 2605 24361 2639 24395
rect 3985 24361 4019 24395
rect 5457 24361 5491 24395
rect 7849 24361 7883 24395
rect 12909 24361 12943 24395
rect 17509 24361 17543 24395
rect 18061 24361 18095 24395
rect 18705 24361 18739 24395
rect 19625 24361 19659 24395
rect 20177 24361 20211 24395
rect 6469 24293 6503 24327
rect 9689 24225 9723 24259
rect 12449 24225 12483 24259
rect 15669 24225 15703 24259
rect 16313 24225 16347 24259
rect 1869 24157 1903 24191
rect 2513 24157 2547 24191
rect 3157 24157 3191 24191
rect 6653 24157 6687 24191
rect 7113 24157 7147 24191
rect 7757 24157 7791 24191
rect 8401 24157 8435 24191
rect 8493 24157 8527 24191
rect 10701 24157 10735 24191
rect 10885 24157 10919 24191
rect 12265 24157 12299 24191
rect 13553 24157 13587 24191
rect 14381 24157 14415 24191
rect 15025 24157 15059 24191
rect 16957 24157 16991 24191
rect 17601 24157 17635 24191
rect 18613 24157 18647 24191
rect 19533 24157 19567 24191
rect 6009 24089 6043 24123
rect 9229 24089 9263 24123
rect 9321 24089 9355 24123
rect 14565 24089 14599 24123
rect 15761 24089 15795 24123
rect 4813 24021 4847 24055
rect 7205 24021 7239 24055
rect 11345 24021 11379 24055
rect 13645 24021 13679 24055
rect 16865 24021 16899 24055
rect 1961 23817 1995 23851
rect 3249 23817 3283 23851
rect 4261 23817 4295 23851
rect 5089 23817 5123 23851
rect 7849 23817 7883 23851
rect 11713 23817 11747 23851
rect 16957 23817 16991 23851
rect 5917 23749 5951 23783
rect 9689 23749 9723 23783
rect 10517 23749 10551 23783
rect 11069 23749 11103 23783
rect 13461 23749 13495 23783
rect 15669 23749 15703 23783
rect 18153 23749 18187 23783
rect 18705 23749 18739 23783
rect 2053 23681 2087 23715
rect 7113 23681 7147 23715
rect 7757 23681 7791 23715
rect 8401 23681 8435 23715
rect 8493 23681 8527 23715
rect 9229 23681 9263 23715
rect 12357 23681 12391 23715
rect 14473 23681 14507 23715
rect 17049 23681 17083 23715
rect 38025 23681 38059 23715
rect 9045 23613 9079 23647
rect 10425 23613 10459 23647
rect 12173 23613 12207 23647
rect 13369 23613 13403 23647
rect 15761 23613 15795 23647
rect 18061 23613 18095 23647
rect 19165 23613 19199 23647
rect 7205 23545 7239 23579
rect 13921 23545 13955 23579
rect 15209 23545 15243 23579
rect 19717 23545 19751 23579
rect 2605 23477 2639 23511
rect 6653 23477 6687 23511
rect 14565 23477 14599 23511
rect 38209 23477 38243 23511
rect 2973 23273 3007 23307
rect 3985 23273 4019 23307
rect 4629 23273 4663 23307
rect 5181 23273 5215 23307
rect 5733 23273 5767 23307
rect 6745 23273 6779 23307
rect 9689 23273 9723 23307
rect 12081 23273 12115 23307
rect 17785 23273 17819 23307
rect 27261 23273 27295 23307
rect 27997 23273 28031 23307
rect 8493 23205 8527 23239
rect 14381 23205 14415 23239
rect 18429 23205 18463 23239
rect 7941 23137 7975 23171
rect 10793 23137 10827 23171
rect 16681 23137 16715 23171
rect 1961 23069 1995 23103
rect 2421 23069 2455 23103
rect 7205 23069 7239 23103
rect 8401 23069 8435 23103
rect 9597 23069 9631 23103
rect 11437 23069 11471 23103
rect 12541 23069 12575 23103
rect 12725 23069 12759 23103
rect 13461 23069 13495 23103
rect 17325 23069 17359 23103
rect 27905 23069 27939 23103
rect 10333 23001 10367 23035
rect 10425 23001 10459 23035
rect 14841 23001 14875 23035
rect 14933 23001 14967 23035
rect 16037 23001 16071 23035
rect 16129 23001 16163 23035
rect 1777 22933 1811 22967
rect 11529 22933 11563 22967
rect 13369 22933 13403 22967
rect 17233 22933 17267 22967
rect 3433 22729 3467 22763
rect 3985 22729 4019 22763
rect 4905 22729 4939 22763
rect 6561 22729 6595 22763
rect 7297 22729 7331 22763
rect 9045 22729 9079 22763
rect 5365 22661 5399 22695
rect 8401 22661 8435 22695
rect 9689 22661 9723 22695
rect 13001 22661 13035 22695
rect 14197 22661 14231 22695
rect 17141 22661 17175 22695
rect 18429 22661 18463 22695
rect 19165 22661 19199 22695
rect 1869 22593 1903 22627
rect 8309 22593 8343 22627
rect 8953 22593 8987 22627
rect 9597 22593 9631 22627
rect 10241 22593 10275 22627
rect 11069 22593 11103 22627
rect 11713 22593 11747 22627
rect 15209 22593 15243 22627
rect 15393 22593 15427 22627
rect 18337 22593 18371 22627
rect 6009 22525 6043 22559
rect 7849 22525 7883 22559
rect 11897 22525 11931 22559
rect 12909 22525 12943 22559
rect 14105 22525 14139 22559
rect 17049 22525 17083 22559
rect 17325 22525 17359 22559
rect 19073 22525 19107 22559
rect 19349 22525 19383 22559
rect 1685 22457 1719 22491
rect 13461 22457 13495 22491
rect 14657 22457 14691 22491
rect 15577 22457 15611 22491
rect 2697 22389 2731 22423
rect 10333 22389 10367 22423
rect 10977 22389 11011 22423
rect 12173 22389 12207 22423
rect 5181 22185 5215 22219
rect 6009 22185 6043 22219
rect 6469 22185 6503 22219
rect 8585 22185 8619 22219
rect 2237 22049 2271 22083
rect 4629 22049 4663 22083
rect 7113 22049 7147 22083
rect 10425 22049 10459 22083
rect 11345 22049 11379 22083
rect 12817 22049 12851 22083
rect 14565 22049 14599 22083
rect 15025 22049 15059 22083
rect 15761 22049 15795 22083
rect 1685 21981 1719 22015
rect 3433 21981 3467 22015
rect 7573 21981 7607 22015
rect 12633 21981 12667 22015
rect 15209 21981 15243 22015
rect 15853 21981 15887 22015
rect 16497 21981 16531 22015
rect 10609 21913 10643 21947
rect 10701 21913 10735 21947
rect 11437 21913 11471 21947
rect 11989 21913 12023 21947
rect 17049 21913 17083 21947
rect 18337 21913 18371 21947
rect 2881 21845 2915 21879
rect 4077 21845 4111 21879
rect 9597 21845 9631 21879
rect 13277 21845 13311 21879
rect 16405 21845 16439 21879
rect 17785 21845 17819 21879
rect 2421 21641 2455 21675
rect 3801 21641 3835 21675
rect 4997 21641 5031 21675
rect 5825 21641 5859 21675
rect 6561 21641 6595 21675
rect 11161 21641 11195 21675
rect 12173 21641 12207 21675
rect 3249 21573 3283 21607
rect 14105 21573 14139 21607
rect 1685 21505 1719 21539
rect 1869 21505 1903 21539
rect 10517 21505 10551 21539
rect 13461 21505 13495 21539
rect 14381 21505 14415 21539
rect 15669 21505 15703 21539
rect 38025 21505 38059 21539
rect 9505 21437 9539 21471
rect 10701 21437 10735 21471
rect 12633 21437 12667 21471
rect 12817 21437 12851 21471
rect 15853 21437 15887 21471
rect 17325 21437 17359 21471
rect 17509 21437 17543 21471
rect 15485 21369 15519 21403
rect 4445 21301 4479 21335
rect 10057 21301 10091 21335
rect 13553 21301 13587 21335
rect 16865 21301 16899 21335
rect 38209 21301 38243 21335
rect 1593 21097 1627 21131
rect 3157 21097 3191 21131
rect 4077 21097 4111 21131
rect 4629 21097 4663 21131
rect 5181 21097 5215 21131
rect 11621 21097 11655 21131
rect 16681 21097 16715 21131
rect 17969 21097 18003 21131
rect 2697 21029 2731 21063
rect 12449 21029 12483 21063
rect 10977 20961 11011 20995
rect 12909 20961 12943 20995
rect 14289 20961 14323 20995
rect 17325 20961 17359 20995
rect 10885 20893 10919 20927
rect 11529 20893 11563 20927
rect 13093 20893 13127 20927
rect 16589 20893 16623 20927
rect 17417 20893 17451 20927
rect 12265 20825 12299 20859
rect 14841 20825 14875 20859
rect 14933 20825 14967 20859
rect 15669 20825 15703 20859
rect 5641 20757 5675 20791
rect 10425 20757 10459 20791
rect 13553 20757 13587 20791
rect 15577 20757 15611 20791
rect 1593 20553 1627 20587
rect 2237 20553 2271 20587
rect 3617 20553 3651 20587
rect 4169 20553 4203 20587
rect 5273 20553 5307 20587
rect 10425 20553 10459 20587
rect 11069 20553 11103 20587
rect 13185 20553 13219 20587
rect 16957 20553 16991 20587
rect 2789 20485 2823 20519
rect 4721 20485 4755 20519
rect 12265 20485 12299 20519
rect 13829 20485 13863 20519
rect 16037 20485 16071 20519
rect 16129 20485 16163 20519
rect 9873 20417 9907 20451
rect 10517 20417 10551 20451
rect 11161 20417 11195 20451
rect 13093 20417 13127 20451
rect 13737 20417 13771 20451
rect 14841 20417 14875 20451
rect 11713 20349 11747 20383
rect 12357 20349 12391 20383
rect 14381 20349 14415 20383
rect 15025 20349 15059 20383
rect 15577 20281 15611 20315
rect 1685 20009 1719 20043
rect 2237 20009 2271 20043
rect 2881 20009 2915 20043
rect 3341 20009 3375 20043
rect 4077 20009 4111 20043
rect 12265 20009 12299 20043
rect 13001 20009 13035 20043
rect 13645 20009 13679 20043
rect 16681 20009 16715 20043
rect 15393 19873 15427 19907
rect 16037 19873 16071 19907
rect 38025 19873 38059 19907
rect 12357 19805 12391 19839
rect 13093 19805 13127 19839
rect 13737 19805 13771 19839
rect 14473 19805 14507 19839
rect 38301 19805 38335 19839
rect 15945 19737 15979 19771
rect 10609 19669 10643 19703
rect 11253 19669 11287 19703
rect 14289 19669 14323 19703
rect 11989 19465 12023 19499
rect 12725 19465 12759 19499
rect 14749 19465 14783 19499
rect 38301 19465 38335 19499
rect 1685 19329 1719 19363
rect 2329 19261 2363 19295
rect 13277 19261 13311 19295
rect 15209 19261 15243 19295
rect 1869 19193 1903 19227
rect 14013 19193 14047 19227
rect 2881 19125 2915 19159
rect 16313 19125 16347 19159
rect 1593 18921 1627 18955
rect 2237 18921 2271 18955
rect 4997 18921 5031 18955
rect 13553 18921 13587 18955
rect 19533 18921 19567 18955
rect 4445 18717 4479 18751
rect 19625 18717 19659 18751
rect 4261 18581 4295 18615
rect 20177 18581 20211 18615
rect 1869 18241 1903 18275
rect 29469 18241 29503 18275
rect 1685 18037 1719 18071
rect 29377 18037 29411 18071
rect 19809 17289 19843 17323
rect 6837 17153 6871 17187
rect 19901 17153 19935 17187
rect 6745 16949 6779 16983
rect 20453 16949 20487 16983
rect 1869 16065 1903 16099
rect 38025 16065 38059 16099
rect 38301 15997 38335 16031
rect 1685 15861 1719 15895
rect 38301 15657 38335 15691
rect 7113 15453 7147 15487
rect 7021 15317 7055 15351
rect 2513 14569 2547 14603
rect 38025 14433 38059 14467
rect 1961 14365 1995 14399
rect 38301 14365 38335 14399
rect 1777 14229 1811 14263
rect 38301 14025 38335 14059
rect 1869 13957 1903 13991
rect 1685 13889 1719 13923
rect 2513 13889 2547 13923
rect 2421 13821 2455 13855
rect 1593 13481 1627 13515
rect 1869 12801 1903 12835
rect 37565 12801 37599 12835
rect 38209 12801 38243 12835
rect 38025 12665 38059 12699
rect 1685 12597 1719 12631
rect 15577 12393 15611 12427
rect 15669 12189 15703 12223
rect 37841 12189 37875 12223
rect 16129 12053 16163 12087
rect 38025 12053 38059 12087
rect 10793 11101 10827 11135
rect 11437 11101 11471 11135
rect 38025 11101 38059 11135
rect 10885 11033 10919 11067
rect 37565 11033 37599 11067
rect 38209 11033 38243 11067
rect 8953 10761 8987 10795
rect 11805 10761 11839 10795
rect 25421 10761 25455 10795
rect 1869 10625 1903 10659
rect 8861 10625 8895 10659
rect 11897 10625 11931 10659
rect 18981 10625 19015 10659
rect 19625 10625 19659 10659
rect 25513 10625 25547 10659
rect 25973 10625 26007 10659
rect 19073 10489 19107 10523
rect 1685 10421 1719 10455
rect 12449 10421 12483 10455
rect 16865 10217 16899 10251
rect 16129 10013 16163 10047
rect 16221 9945 16255 9979
rect 16313 9061 16347 9095
rect 14749 8925 14783 8959
rect 15393 8925 15427 8959
rect 16129 8925 16163 8959
rect 16773 8925 16807 8959
rect 38025 8925 38059 8959
rect 1685 8857 1719 8891
rect 1777 8789 1811 8823
rect 14933 8789 14967 8823
rect 38209 8789 38243 8823
rect 1685 8585 1719 8619
rect 38025 7429 38059 7463
rect 22385 7361 22419 7395
rect 23029 7361 23063 7395
rect 37565 7361 37599 7395
rect 38209 7361 38243 7395
rect 1593 7293 1627 7327
rect 1869 7293 1903 7327
rect 22569 7157 22603 7191
rect 1593 6953 1627 6987
rect 24409 6273 24443 6307
rect 25053 6273 25087 6307
rect 24593 6069 24627 6103
rect 38117 5865 38151 5899
rect 37565 5593 37599 5627
rect 38209 5593 38243 5627
rect 1777 5321 1811 5355
rect 1685 5185 1719 5219
rect 1593 4777 1627 4811
rect 1685 3893 1719 3927
rect 38209 3893 38243 3927
rect 1869 3621 1903 3655
rect 1685 3485 1719 3519
rect 38025 3485 38059 3519
rect 37473 3349 37507 3383
rect 38209 3349 38243 3383
rect 12725 3145 12759 3179
rect 20729 3145 20763 3179
rect 34713 3145 34747 3179
rect 29745 3077 29779 3111
rect 38025 3077 38059 3111
rect 1869 3009 1903 3043
rect 8677 3009 8711 3043
rect 12265 3009 12299 3043
rect 18705 3009 18739 3043
rect 19349 3009 19383 3043
rect 21281 3009 21315 3043
rect 29009 3009 29043 3043
rect 36921 3009 36955 3043
rect 38209 3009 38243 3043
rect 2421 2941 2455 2975
rect 37473 2941 37507 2975
rect 12081 2873 12115 2907
rect 18889 2873 18923 2907
rect 1685 2805 1719 2839
rect 4537 2805 4571 2839
rect 8493 2805 8527 2839
rect 21373 2805 21407 2839
rect 29193 2805 29227 2839
rect 36369 2805 36403 2839
rect 4169 2601 4203 2635
rect 28549 2601 28583 2635
rect 33701 2601 33735 2635
rect 36001 2601 36035 2635
rect 2421 2533 2455 2567
rect 4629 2533 4663 2567
rect 11989 2533 12023 2567
rect 15209 2533 15243 2567
rect 32321 2533 32355 2567
rect 36645 2533 36679 2567
rect 10057 2465 10091 2499
rect 38025 2465 38059 2499
rect 1869 2397 1903 2431
rect 2605 2397 2639 2431
rect 3985 2397 4019 2431
rect 6837 2397 6871 2431
rect 8585 2397 8619 2431
rect 9321 2397 9355 2431
rect 9781 2397 9815 2431
rect 13001 2397 13035 2431
rect 16865 2397 16899 2431
rect 18153 2397 18187 2431
rect 20085 2397 20119 2431
rect 22017 2397 22051 2431
rect 23305 2397 23339 2431
rect 25237 2397 25271 2431
rect 27169 2397 27203 2431
rect 29745 2397 29779 2431
rect 34897 2397 34931 2431
rect 36185 2397 36219 2431
rect 38301 2397 38335 2431
rect 4813 2329 4847 2363
rect 11161 2329 11195 2363
rect 11805 2329 11839 2363
rect 14473 2329 14507 2363
rect 15025 2329 15059 2363
rect 27997 2329 28031 2363
rect 28641 2329 28675 2363
rect 32505 2329 32539 2363
rect 33149 2329 33183 2363
rect 33793 2329 33827 2363
rect 36829 2329 36863 2363
rect 1685 2261 1719 2295
rect 3341 2261 3375 2295
rect 6653 2261 6687 2295
rect 8401 2261 8435 2295
rect 13185 2261 13219 2295
rect 17049 2261 17083 2295
rect 18337 2261 18371 2295
rect 20269 2261 20303 2295
rect 22201 2261 22235 2295
rect 23489 2261 23523 2295
rect 25421 2261 25455 2295
rect 27353 2261 27387 2295
rect 29929 2261 29963 2295
rect 31769 2261 31803 2295
rect 35081 2261 35115 2295
<< metal1 >>
rect 14274 37680 14280 37732
rect 14332 37720 14338 37732
rect 21542 37720 21548 37732
rect 14332 37692 21548 37720
rect 14332 37680 14338 37692
rect 21542 37680 21548 37692
rect 21600 37680 21606 37732
rect 13170 37612 13176 37664
rect 13228 37652 13234 37664
rect 16114 37652 16120 37664
rect 13228 37624 16120 37652
rect 13228 37612 13234 37624
rect 16114 37612 16120 37624
rect 16172 37612 16178 37664
rect 16482 37612 16488 37664
rect 16540 37652 16546 37664
rect 18874 37652 18880 37664
rect 16540 37624 18880 37652
rect 16540 37612 16546 37624
rect 18874 37612 18880 37624
rect 18932 37612 18938 37664
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 8202 37408 8208 37460
rect 8260 37448 8266 37460
rect 22830 37448 22836 37460
rect 8260 37420 22836 37448
rect 8260 37408 8266 37420
rect 22830 37408 22836 37420
rect 22888 37408 22894 37460
rect 38194 37408 38200 37460
rect 38252 37448 38258 37460
rect 38289 37451 38347 37457
rect 38289 37448 38301 37451
rect 38252 37420 38301 37448
rect 38252 37408 38258 37420
rect 38289 37417 38301 37420
rect 38335 37448 38347 37451
rect 38654 37448 38660 37460
rect 38335 37420 38660 37448
rect 38335 37417 38347 37420
rect 38289 37411 38347 37417
rect 38654 37408 38660 37420
rect 38712 37408 38718 37460
rect 16022 37380 16028 37392
rect 8496 37352 9536 37380
rect 15983 37352 16028 37380
rect 14 37272 20 37324
rect 72 37312 78 37324
rect 2314 37312 2320 37324
rect 72 37284 2320 37312
rect 72 37272 78 37284
rect 2314 37272 2320 37284
rect 2372 37272 2378 37324
rect 5721 37315 5779 37321
rect 5721 37281 5733 37315
rect 5767 37312 5779 37315
rect 6546 37312 6552 37324
rect 5767 37284 6552 37312
rect 5767 37281 5779 37284
rect 5721 37275 5779 37281
rect 6546 37272 6552 37284
rect 6604 37272 6610 37324
rect 7101 37315 7159 37321
rect 7101 37281 7113 37315
rect 7147 37312 7159 37315
rect 8496 37312 8524 37352
rect 7147 37284 8524 37312
rect 8573 37315 8631 37321
rect 7147 37281 7159 37284
rect 7101 37275 7159 37281
rect 8573 37281 8585 37315
rect 8619 37312 8631 37315
rect 9508 37312 9536 37352
rect 16022 37340 16028 37352
rect 16080 37340 16086 37392
rect 16390 37340 16396 37392
rect 16448 37380 16454 37392
rect 16448 37352 18368 37380
rect 16448 37340 16454 37352
rect 11238 37312 11244 37324
rect 8619 37284 9076 37312
rect 9508 37284 11244 37312
rect 8619 37281 8631 37284
rect 8573 37275 8631 37281
rect 1670 37244 1676 37256
rect 1631 37216 1676 37244
rect 1670 37204 1676 37216
rect 1728 37204 1734 37256
rect 4614 37204 4620 37256
rect 4672 37204 4678 37256
rect 5997 37247 6055 37253
rect 5997 37213 6009 37247
rect 6043 37244 6055 37247
rect 6825 37247 6883 37253
rect 6825 37244 6837 37247
rect 6043 37216 6837 37244
rect 6043 37213 6055 37216
rect 5997 37207 6055 37213
rect 6825 37213 6837 37216
rect 6871 37213 6883 37247
rect 6825 37207 6883 37213
rect 1854 37136 1860 37188
rect 1912 37176 1918 37188
rect 1949 37179 2007 37185
rect 1949 37176 1961 37179
rect 1912 37148 1961 37176
rect 1912 37136 1918 37148
rect 1949 37145 1961 37148
rect 1995 37145 2007 37179
rect 1949 37139 2007 37145
rect 2682 37136 2688 37188
rect 2740 37136 2746 37188
rect 3878 37136 3884 37188
rect 3936 37176 3942 37188
rect 6012 37176 6040 37207
rect 8202 37204 8208 37256
rect 8260 37204 8266 37256
rect 3936 37148 4476 37176
rect 3936 37136 3942 37148
rect 3326 37068 3332 37120
rect 3384 37108 3390 37120
rect 3421 37111 3479 37117
rect 3421 37108 3433 37111
rect 3384 37080 3433 37108
rect 3384 37068 3390 37080
rect 3421 37077 3433 37080
rect 3467 37077 3479 37111
rect 4246 37108 4252 37120
rect 4207 37080 4252 37108
rect 3421 37071 3479 37077
rect 4246 37068 4252 37080
rect 4304 37068 4310 37120
rect 4448 37108 4476 37148
rect 5920 37148 6040 37176
rect 9048 37176 9076 37284
rect 11238 37272 11244 37284
rect 11296 37272 11302 37324
rect 13170 37312 13176 37324
rect 13131 37284 13176 37312
rect 13170 37272 13176 37284
rect 13228 37272 13234 37324
rect 14550 37272 14556 37324
rect 14608 37312 14614 37324
rect 14608 37284 16620 37312
rect 14608 37272 14614 37284
rect 9122 37204 9128 37256
rect 9180 37244 9186 37256
rect 9401 37247 9459 37253
rect 9401 37244 9413 37247
rect 9180 37216 9413 37244
rect 9180 37204 9186 37216
rect 9401 37213 9413 37216
rect 9447 37213 9459 37247
rect 9401 37207 9459 37213
rect 13449 37247 13507 37253
rect 13449 37213 13461 37247
rect 13495 37244 13507 37247
rect 13998 37244 14004 37256
rect 13495 37216 14004 37244
rect 13495 37213 13507 37216
rect 13449 37207 13507 37213
rect 13998 37204 14004 37216
rect 14056 37244 14062 37256
rect 14277 37247 14335 37253
rect 14277 37244 14289 37247
rect 14056 37216 14289 37244
rect 14056 37204 14062 37216
rect 14277 37213 14289 37216
rect 14323 37213 14335 37247
rect 16482 37244 16488 37256
rect 15686 37216 16488 37244
rect 14277 37207 14335 37213
rect 16482 37204 16488 37216
rect 16540 37204 16546 37256
rect 16592 37244 16620 37284
rect 16666 37272 16672 37324
rect 16724 37312 16730 37324
rect 18340 37312 18368 37352
rect 21542 37340 21548 37392
rect 21600 37380 21606 37392
rect 23385 37383 23443 37389
rect 23385 37380 23397 37383
rect 21600 37352 23397 37380
rect 21600 37340 21606 37352
rect 23385 37349 23397 37352
rect 23431 37349 23443 37383
rect 23385 37343 23443 37349
rect 19242 37312 19248 37324
rect 16724 37284 17264 37312
rect 18340 37284 19248 37312
rect 16724 37272 16730 37284
rect 16850 37244 16856 37256
rect 16592 37216 16856 37244
rect 16850 37204 16856 37216
rect 16908 37204 16914 37256
rect 17126 37244 17132 37256
rect 17087 37216 17132 37244
rect 17126 37204 17132 37216
rect 17184 37204 17190 37256
rect 17236 37244 17264 37284
rect 18432 37253 18460 37284
rect 19242 37272 19248 37284
rect 19300 37312 19306 37324
rect 20165 37315 20223 37321
rect 20165 37312 20177 37315
rect 19300 37284 20177 37312
rect 19300 37272 19306 37284
rect 20165 37281 20177 37284
rect 20211 37281 20223 37315
rect 23934 37312 23940 37324
rect 20165 37275 20223 37281
rect 20640 37284 21496 37312
rect 23895 37284 23940 37312
rect 17773 37247 17831 37253
rect 17773 37244 17785 37247
rect 17236 37216 17785 37244
rect 17773 37213 17785 37216
rect 17819 37244 17831 37247
rect 18417 37247 18475 37253
rect 17819 37216 18368 37244
rect 17819 37213 17831 37216
rect 17773 37207 17831 37213
rect 9582 37176 9588 37188
rect 9048 37148 9588 37176
rect 5920 37108 5948 37148
rect 9582 37136 9588 37148
rect 9640 37176 9646 37188
rect 9677 37179 9735 37185
rect 9677 37176 9689 37179
rect 9640 37148 9689 37176
rect 9640 37136 9646 37148
rect 9677 37145 9689 37148
rect 9723 37145 9735 37179
rect 9677 37139 9735 37145
rect 10686 37136 10692 37188
rect 10744 37136 10750 37188
rect 12710 37136 12716 37188
rect 12768 37136 12774 37188
rect 12894 37136 12900 37188
rect 12952 37176 12958 37188
rect 14182 37176 14188 37188
rect 12952 37148 14188 37176
rect 12952 37136 12958 37148
rect 14182 37136 14188 37148
rect 14240 37136 14246 37188
rect 14553 37179 14611 37185
rect 14553 37145 14565 37179
rect 14599 37176 14611 37179
rect 14642 37176 14648 37188
rect 14599 37148 14648 37176
rect 14599 37145 14611 37148
rect 14553 37139 14611 37145
rect 14642 37136 14648 37148
rect 14700 37136 14706 37188
rect 18340 37176 18368 37216
rect 18417 37213 18429 37247
rect 18463 37213 18475 37247
rect 19426 37244 19432 37256
rect 19387 37216 19432 37244
rect 18417 37207 18475 37213
rect 19426 37204 19432 37216
rect 19484 37204 19490 37256
rect 19978 37204 19984 37256
rect 20036 37244 20042 37256
rect 20640 37244 20668 37284
rect 20036 37216 20668 37244
rect 20036 37204 20042 37216
rect 20714 37204 20720 37256
rect 20772 37244 20778 37256
rect 20901 37247 20959 37253
rect 20901 37244 20913 37247
rect 20772 37216 20913 37244
rect 20772 37204 20778 37216
rect 20901 37213 20913 37216
rect 20947 37244 20959 37247
rect 21361 37247 21419 37253
rect 21361 37244 21373 37247
rect 20947 37216 21373 37244
rect 20947 37213 20959 37216
rect 20901 37207 20959 37213
rect 21361 37213 21373 37216
rect 21407 37213 21419 37247
rect 21468 37244 21496 37284
rect 23934 37272 23940 37284
rect 23992 37272 23998 37324
rect 29089 37315 29147 37321
rect 24504 37284 24716 37312
rect 22005 37247 22063 37253
rect 22005 37244 22017 37247
rect 21468 37216 22017 37244
rect 21361 37207 21419 37213
rect 22005 37213 22017 37216
rect 22051 37213 22063 37247
rect 22738 37244 22744 37256
rect 22699 37216 22744 37244
rect 22005 37207 22063 37213
rect 22738 37204 22744 37216
rect 22796 37204 22802 37256
rect 24504 37244 24532 37284
rect 23768 37216 24532 37244
rect 24581 37247 24639 37253
rect 15856 37148 18276 37176
rect 18340 37148 19748 37176
rect 4448 37080 5948 37108
rect 5994 37068 6000 37120
rect 6052 37108 6058 37120
rect 10962 37108 10968 37120
rect 6052 37080 10968 37108
rect 6052 37068 6058 37080
rect 10962 37068 10968 37080
rect 11020 37068 11026 37120
rect 11146 37108 11152 37120
rect 11107 37080 11152 37108
rect 11146 37068 11152 37080
rect 11204 37068 11210 37120
rect 11698 37108 11704 37120
rect 11659 37080 11704 37108
rect 11698 37068 11704 37080
rect 11756 37068 11762 37120
rect 12526 37068 12532 37120
rect 12584 37108 12590 37120
rect 15856 37108 15884 37148
rect 12584 37080 15884 37108
rect 12584 37068 12590 37080
rect 16022 37068 16028 37120
rect 16080 37108 16086 37120
rect 16574 37108 16580 37120
rect 16080 37080 16580 37108
rect 16080 37068 16086 37080
rect 16574 37068 16580 37080
rect 16632 37068 16638 37120
rect 16758 37068 16764 37120
rect 16816 37108 16822 37120
rect 16945 37111 17003 37117
rect 16945 37108 16957 37111
rect 16816 37080 16957 37108
rect 16816 37068 16822 37080
rect 16945 37077 16957 37080
rect 16991 37077 17003 37111
rect 17678 37108 17684 37120
rect 17639 37080 17684 37108
rect 16945 37071 17003 37077
rect 17678 37068 17684 37080
rect 17736 37068 17742 37120
rect 18248 37117 18276 37148
rect 18233 37111 18291 37117
rect 18233 37077 18245 37111
rect 18279 37077 18291 37111
rect 18233 37071 18291 37077
rect 18690 37068 18696 37120
rect 18748 37108 18754 37120
rect 19613 37111 19671 37117
rect 19613 37108 19625 37111
rect 18748 37080 19625 37108
rect 18748 37068 18754 37080
rect 19613 37077 19625 37080
rect 19659 37077 19671 37111
rect 19720 37108 19748 37148
rect 20438 37136 20444 37188
rect 20496 37176 20502 37188
rect 23768 37176 23796 37216
rect 24581 37213 24593 37247
rect 24627 37213 24639 37247
rect 24688 37244 24716 37284
rect 29089 37281 29101 37315
rect 29135 37312 29147 37315
rect 29178 37312 29184 37324
rect 29135 37284 29184 37312
rect 29135 37281 29147 37284
rect 29089 37275 29147 37281
rect 29178 37272 29184 37284
rect 29236 37272 29242 37324
rect 35069 37315 35127 37321
rect 35069 37281 35081 37315
rect 35115 37312 35127 37315
rect 35434 37312 35440 37324
rect 35115 37284 35440 37312
rect 35115 37281 35127 37284
rect 35069 37275 35127 37281
rect 35434 37272 35440 37284
rect 35492 37312 35498 37324
rect 35529 37315 35587 37321
rect 35529 37312 35541 37315
rect 35492 37284 35541 37312
rect 35492 37272 35498 37284
rect 35529 37281 35541 37284
rect 35575 37281 35587 37315
rect 35529 37275 35587 37281
rect 25314 37244 25320 37256
rect 24688 37216 24900 37244
rect 25275 37216 25320 37244
rect 24581 37207 24639 37213
rect 20496 37148 23796 37176
rect 20496 37136 20502 37148
rect 20717 37111 20775 37117
rect 20717 37108 20729 37111
rect 19720 37080 20729 37108
rect 19613 37071 19671 37077
rect 20717 37077 20729 37080
rect 20763 37077 20775 37111
rect 20717 37071 20775 37077
rect 21910 37068 21916 37120
rect 21968 37108 21974 37120
rect 22189 37111 22247 37117
rect 22189 37108 22201 37111
rect 21968 37080 22201 37108
rect 21968 37068 21974 37080
rect 22189 37077 22201 37080
rect 22235 37077 22247 37111
rect 22189 37071 22247 37077
rect 22646 37068 22652 37120
rect 22704 37108 22710 37120
rect 22833 37111 22891 37117
rect 22833 37108 22845 37111
rect 22704 37080 22845 37108
rect 22704 37068 22710 37080
rect 22833 37077 22845 37080
rect 22879 37077 22891 37111
rect 22833 37071 22891 37077
rect 22922 37068 22928 37120
rect 22980 37108 22986 37120
rect 24596 37108 24624 37207
rect 24872 37176 24900 37216
rect 25314 37204 25320 37216
rect 25372 37204 25378 37256
rect 26510 37204 26516 37256
rect 26568 37244 26574 37256
rect 27157 37247 27215 37253
rect 27157 37244 27169 37247
rect 26568 37216 27169 37244
rect 26568 37204 26574 37216
rect 27157 37213 27169 37216
rect 27203 37213 27215 37247
rect 29730 37244 29736 37256
rect 29691 37216 29736 37244
rect 27157 37207 27215 37213
rect 29730 37204 29736 37216
rect 29788 37204 29794 37256
rect 30374 37204 30380 37256
rect 30432 37244 30438 37256
rect 30653 37247 30711 37253
rect 30653 37244 30665 37247
rect 30432 37216 30665 37244
rect 30432 37204 30438 37216
rect 30653 37213 30665 37216
rect 30699 37244 30711 37247
rect 31113 37247 31171 37253
rect 31113 37244 31125 37247
rect 30699 37216 31125 37244
rect 30699 37213 30711 37216
rect 30653 37207 30711 37213
rect 31113 37213 31125 37216
rect 31159 37213 31171 37247
rect 32306 37244 32312 37256
rect 32267 37216 32312 37244
rect 31113 37207 31171 37213
rect 32306 37204 32312 37216
rect 32364 37204 32370 37256
rect 33873 37247 33931 37253
rect 33873 37213 33885 37247
rect 33919 37244 33931 37247
rect 33962 37244 33968 37256
rect 33919 37216 33968 37244
rect 33919 37213 33931 37216
rect 33873 37207 33931 37213
rect 33962 37204 33968 37216
rect 34020 37204 34026 37256
rect 35805 37247 35863 37253
rect 35805 37213 35817 37247
rect 35851 37213 35863 37247
rect 37461 37247 37519 37253
rect 37461 37244 37473 37247
rect 35805 37207 35863 37213
rect 36832 37216 37473 37244
rect 24872 37148 30512 37176
rect 24762 37108 24768 37120
rect 22980 37080 24624 37108
rect 24723 37080 24768 37108
rect 22980 37068 22986 37080
rect 24762 37068 24768 37080
rect 24820 37068 24826 37120
rect 25130 37068 25136 37120
rect 25188 37108 25194 37120
rect 25501 37111 25559 37117
rect 25501 37108 25513 37111
rect 25188 37080 25513 37108
rect 25188 37068 25194 37080
rect 25501 37077 25513 37080
rect 25547 37077 25559 37111
rect 26510 37108 26516 37120
rect 26471 37080 26516 37108
rect 25501 37071 25559 37077
rect 26510 37068 26516 37080
rect 26568 37068 26574 37120
rect 27062 37068 27068 37120
rect 27120 37108 27126 37120
rect 27341 37111 27399 37117
rect 27341 37108 27353 37111
rect 27120 37080 27353 37108
rect 27120 37068 27126 37080
rect 27341 37077 27353 37080
rect 27387 37077 27399 37111
rect 27341 37071 27399 37077
rect 27985 37111 28043 37117
rect 27985 37077 27997 37111
rect 28031 37108 28043 37111
rect 28442 37108 28448 37120
rect 28031 37080 28448 37108
rect 28031 37077 28043 37080
rect 27985 37071 28043 37077
rect 28442 37068 28448 37080
rect 28500 37068 28506 37120
rect 28994 37068 29000 37120
rect 29052 37108 29058 37120
rect 30484 37117 30512 37148
rect 30558 37136 30564 37188
rect 30616 37176 30622 37188
rect 35820 37176 35848 37207
rect 30616 37148 35848 37176
rect 30616 37136 30622 37148
rect 36832 37120 36860 37216
rect 37461 37213 37473 37216
rect 37507 37213 37519 37247
rect 37461 37207 37519 37213
rect 29917 37111 29975 37117
rect 29917 37108 29929 37111
rect 29052 37080 29929 37108
rect 29052 37068 29058 37080
rect 29917 37077 29929 37080
rect 29963 37077 29975 37111
rect 29917 37071 29975 37077
rect 30469 37111 30527 37117
rect 30469 37077 30481 37111
rect 30515 37077 30527 37111
rect 30469 37071 30527 37077
rect 32214 37068 32220 37120
rect 32272 37108 32278 37120
rect 32493 37111 32551 37117
rect 32493 37108 32505 37111
rect 32272 37080 32505 37108
rect 32272 37068 32278 37080
rect 32493 37077 32505 37080
rect 32539 37077 32551 37111
rect 32493 37071 32551 37077
rect 33502 37068 33508 37120
rect 33560 37108 33566 37120
rect 33689 37111 33747 37117
rect 33689 37108 33701 37111
rect 33560 37080 33701 37108
rect 33560 37068 33566 37080
rect 33689 37077 33701 37080
rect 33735 37077 33747 37111
rect 36814 37108 36820 37120
rect 36775 37080 36820 37108
rect 33689 37071 33747 37077
rect 36814 37068 36820 37080
rect 36872 37068 36878 37120
rect 37366 37068 37372 37120
rect 37424 37108 37430 37120
rect 37645 37111 37703 37117
rect 37645 37108 37657 37111
rect 37424 37080 37657 37108
rect 37424 37068 37430 37080
rect 37645 37077 37657 37080
rect 37691 37077 37703 37111
rect 37645 37071 37703 37077
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 1670 36864 1676 36916
rect 1728 36904 1734 36916
rect 3878 36904 3884 36916
rect 1728 36876 3884 36904
rect 1728 36864 1734 36876
rect 3878 36864 3884 36876
rect 3936 36864 3942 36916
rect 5902 36904 5908 36916
rect 4908 36876 5908 36904
rect 934 36796 940 36848
rect 992 36836 998 36848
rect 3513 36839 3571 36845
rect 992 36808 2346 36836
rect 992 36796 998 36808
rect 3513 36805 3525 36839
rect 3559 36836 3571 36839
rect 4908 36836 4936 36876
rect 5902 36864 5908 36876
rect 5960 36864 5966 36916
rect 5997 36907 6055 36913
rect 5997 36873 6009 36907
rect 6043 36904 6055 36907
rect 11882 36904 11888 36916
rect 6043 36876 11888 36904
rect 6043 36873 6055 36876
rect 5997 36867 6055 36873
rect 11882 36864 11888 36876
rect 11940 36864 11946 36916
rect 14550 36904 14556 36916
rect 11992 36876 14556 36904
rect 6270 36836 6276 36848
rect 3559 36808 4936 36836
rect 5750 36808 6276 36836
rect 3559 36805 3571 36808
rect 3513 36799 3571 36805
rect 6270 36796 6276 36808
rect 6328 36796 6334 36848
rect 9674 36836 9680 36848
rect 8326 36808 9680 36836
rect 9674 36796 9680 36808
rect 9732 36796 9738 36848
rect 10962 36836 10968 36848
rect 10810 36808 10968 36836
rect 10962 36796 10968 36808
rect 11020 36796 11026 36848
rect 11146 36796 11152 36848
rect 11204 36836 11210 36848
rect 11992 36845 12020 36876
rect 14550 36864 14556 36876
rect 14608 36864 14614 36916
rect 14660 36876 15700 36904
rect 11977 36839 12035 36845
rect 11977 36836 11989 36839
rect 11204 36808 11989 36836
rect 11204 36796 11210 36808
rect 11977 36805 11989 36808
rect 12023 36805 12035 36839
rect 14660 36836 14688 36876
rect 13202 36808 14688 36836
rect 15672 36836 15700 36876
rect 15746 36864 15752 36916
rect 15804 36904 15810 36916
rect 16945 36907 17003 36913
rect 16945 36904 16957 36907
rect 15804 36876 16957 36904
rect 15804 36864 15810 36876
rect 16945 36873 16957 36876
rect 16991 36873 17003 36907
rect 16945 36867 17003 36873
rect 17218 36864 17224 36916
rect 17276 36904 17282 36916
rect 22738 36904 22744 36916
rect 17276 36876 22744 36904
rect 17276 36864 17282 36876
rect 22738 36864 22744 36876
rect 22796 36864 22802 36916
rect 23842 36864 23848 36916
rect 23900 36904 23906 36916
rect 24762 36904 24768 36916
rect 23900 36876 24768 36904
rect 23900 36864 23906 36876
rect 24762 36864 24768 36876
rect 24820 36864 24826 36916
rect 26053 36907 26111 36913
rect 26053 36873 26065 36907
rect 26099 36904 26111 36907
rect 29730 36904 29736 36916
rect 26099 36876 29736 36904
rect 26099 36873 26111 36876
rect 26053 36867 26111 36873
rect 29730 36864 29736 36876
rect 29788 36864 29794 36916
rect 15672 36808 20576 36836
rect 11977 36799 12035 36805
rect 3789 36771 3847 36777
rect 3789 36737 3801 36771
rect 3835 36768 3847 36771
rect 3878 36768 3884 36780
rect 3835 36740 3884 36768
rect 3835 36737 3847 36740
rect 3789 36731 3847 36737
rect 3878 36728 3884 36740
rect 3936 36768 3942 36780
rect 4249 36771 4307 36777
rect 4249 36768 4261 36771
rect 3936 36740 4261 36768
rect 3936 36728 3942 36740
rect 4249 36737 4261 36740
rect 4295 36737 4307 36771
rect 11606 36768 11612 36780
rect 4249 36731 4307 36737
rect 10980 36740 11612 36768
rect 2041 36703 2099 36709
rect 2041 36669 2053 36703
rect 2087 36700 2099 36703
rect 4062 36700 4068 36712
rect 2087 36672 4068 36700
rect 2087 36669 2099 36672
rect 2041 36663 2099 36669
rect 4062 36660 4068 36672
rect 4120 36660 4126 36712
rect 4525 36703 4583 36709
rect 4525 36669 4537 36703
rect 4571 36700 4583 36703
rect 6362 36700 6368 36712
rect 4571 36672 6368 36700
rect 4571 36669 4583 36672
rect 4525 36663 4583 36669
rect 6362 36660 6368 36672
rect 6420 36660 6426 36712
rect 6822 36700 6828 36712
rect 6783 36672 6828 36700
rect 6822 36660 6828 36672
rect 6880 36660 6886 36712
rect 7101 36703 7159 36709
rect 7101 36669 7113 36703
rect 7147 36700 7159 36703
rect 7190 36700 7196 36712
rect 7147 36672 7196 36700
rect 7147 36669 7159 36672
rect 7101 36663 7159 36669
rect 7190 36660 7196 36672
rect 7248 36700 7254 36712
rect 8110 36700 8116 36712
rect 7248 36672 8116 36700
rect 7248 36660 7254 36672
rect 8110 36660 8116 36672
rect 8168 36660 8174 36712
rect 8849 36703 8907 36709
rect 8849 36669 8861 36703
rect 8895 36700 8907 36703
rect 9030 36700 9036 36712
rect 8895 36672 9036 36700
rect 8895 36669 8907 36672
rect 8849 36663 8907 36669
rect 9030 36660 9036 36672
rect 9088 36660 9094 36712
rect 9122 36660 9128 36712
rect 9180 36700 9186 36712
rect 9309 36703 9367 36709
rect 9309 36700 9321 36703
rect 9180 36672 9321 36700
rect 9180 36660 9186 36672
rect 9309 36669 9321 36672
rect 9355 36669 9367 36703
rect 9309 36663 9367 36669
rect 9585 36703 9643 36709
rect 9585 36669 9597 36703
rect 9631 36700 9643 36703
rect 10980 36700 11008 36740
rect 11606 36728 11612 36740
rect 11664 36728 11670 36780
rect 17034 36768 17040 36780
rect 15410 36740 17040 36768
rect 17034 36728 17040 36740
rect 17092 36728 17098 36780
rect 17129 36771 17187 36777
rect 17129 36737 17141 36771
rect 17175 36768 17187 36771
rect 17494 36768 17500 36780
rect 17175 36740 17500 36768
rect 17175 36737 17187 36740
rect 17129 36731 17187 36737
rect 17494 36728 17500 36740
rect 17552 36728 17558 36780
rect 17589 36771 17647 36777
rect 17589 36737 17601 36771
rect 17635 36768 17647 36771
rect 17862 36768 17868 36780
rect 17635 36740 17868 36768
rect 17635 36737 17647 36740
rect 17589 36731 17647 36737
rect 17862 36728 17868 36740
rect 17920 36728 17926 36780
rect 18693 36771 18751 36777
rect 18693 36737 18705 36771
rect 18739 36768 18751 36771
rect 18966 36768 18972 36780
rect 18739 36740 18972 36768
rect 18739 36737 18751 36740
rect 18693 36731 18751 36737
rect 18966 36728 18972 36740
rect 19024 36728 19030 36780
rect 19613 36771 19671 36777
rect 19613 36737 19625 36771
rect 19659 36768 19671 36771
rect 20438 36768 20444 36780
rect 19659 36740 20444 36768
rect 19659 36737 19671 36740
rect 19613 36731 19671 36737
rect 20438 36728 20444 36740
rect 20496 36728 20502 36780
rect 20548 36768 20576 36808
rect 20714 36796 20720 36848
rect 20772 36836 20778 36848
rect 22097 36839 22155 36845
rect 22097 36836 22109 36839
rect 20772 36808 22109 36836
rect 20772 36796 20778 36808
rect 22097 36805 22109 36808
rect 22143 36805 22155 36839
rect 22097 36799 22155 36805
rect 22554 36796 22560 36848
rect 22612 36836 22618 36848
rect 22612 36808 26004 36836
rect 22612 36796 22618 36808
rect 21361 36771 21419 36777
rect 21361 36768 21373 36771
rect 20548 36740 21373 36768
rect 21361 36737 21373 36740
rect 21407 36737 21419 36771
rect 21361 36731 21419 36737
rect 21453 36771 21511 36777
rect 21453 36737 21465 36771
rect 21499 36768 21511 36771
rect 22189 36771 22247 36777
rect 22189 36768 22201 36771
rect 21499 36740 22201 36768
rect 21499 36737 21511 36740
rect 21453 36731 21511 36737
rect 22189 36737 22201 36740
rect 22235 36768 22247 36771
rect 22649 36771 22707 36777
rect 22649 36768 22661 36771
rect 22235 36740 22661 36768
rect 22235 36737 22247 36740
rect 22189 36731 22247 36737
rect 22649 36737 22661 36740
rect 22695 36737 22707 36771
rect 22649 36731 22707 36737
rect 9631 36672 11008 36700
rect 9631 36669 9643 36672
rect 9585 36663 9643 36669
rect 11054 36660 11060 36712
rect 11112 36700 11118 36712
rect 11701 36703 11759 36709
rect 11701 36700 11713 36703
rect 11112 36672 11713 36700
rect 11112 36660 11118 36672
rect 11701 36669 11713 36672
rect 11747 36669 11759 36703
rect 13998 36700 14004 36712
rect 13959 36672 14004 36700
rect 11701 36663 11759 36669
rect 13998 36660 14004 36672
rect 14056 36660 14062 36712
rect 17218 36700 17224 36712
rect 14108 36672 17224 36700
rect 11606 36632 11612 36644
rect 10980 36604 11612 36632
rect 4246 36524 4252 36576
rect 4304 36564 4310 36576
rect 4982 36564 4988 36576
rect 4304 36536 4988 36564
rect 4304 36524 4310 36536
rect 4982 36524 4988 36536
rect 5040 36524 5046 36576
rect 6270 36524 6276 36576
rect 6328 36564 6334 36576
rect 10980 36564 11008 36604
rect 11606 36592 11612 36604
rect 11664 36592 11670 36644
rect 13078 36592 13084 36644
rect 13136 36632 13142 36644
rect 14108 36632 14136 36672
rect 17218 36660 17224 36672
rect 17276 36660 17282 36712
rect 18984 36700 19012 36728
rect 19337 36703 19395 36709
rect 19337 36700 19349 36703
rect 18984 36672 19349 36700
rect 19337 36669 19349 36672
rect 19383 36669 19395 36703
rect 20162 36700 20168 36712
rect 20123 36672 20168 36700
rect 19337 36663 19395 36669
rect 20162 36660 20168 36672
rect 20220 36660 20226 36712
rect 20622 36660 20628 36712
rect 20680 36700 20686 36712
rect 21468 36700 21496 36731
rect 23014 36728 23020 36780
rect 23072 36768 23078 36780
rect 23937 36771 23995 36777
rect 23937 36768 23949 36771
rect 23072 36740 23949 36768
rect 23072 36728 23078 36740
rect 23937 36737 23949 36740
rect 23983 36737 23995 36771
rect 25869 36771 25927 36777
rect 25869 36768 25881 36771
rect 23937 36731 23995 36737
rect 25792 36740 25881 36768
rect 25792 36712 25820 36740
rect 25869 36737 25881 36740
rect 25915 36737 25927 36771
rect 25976 36768 26004 36808
rect 27062 36796 27068 36848
rect 27120 36836 27126 36848
rect 36814 36836 36820 36848
rect 27120 36808 36820 36836
rect 27120 36796 27126 36808
rect 36814 36796 36820 36808
rect 36872 36796 36878 36848
rect 38194 36836 38200 36848
rect 38155 36808 38200 36836
rect 38194 36796 38200 36808
rect 38252 36796 38258 36848
rect 27341 36771 27399 36777
rect 27341 36768 27353 36771
rect 25976 36740 27353 36768
rect 25869 36731 25927 36737
rect 27341 36737 27353 36740
rect 27387 36737 27399 36771
rect 27341 36731 27399 36737
rect 27433 36771 27491 36777
rect 27433 36737 27445 36771
rect 27479 36768 27491 36771
rect 31588 36768 31708 36772
rect 32306 36768 32312 36780
rect 27479 36744 32312 36768
rect 27479 36740 31616 36744
rect 31680 36740 32312 36744
rect 27479 36737 27491 36740
rect 27433 36731 27491 36737
rect 32306 36728 32312 36740
rect 32364 36728 32370 36780
rect 20680 36672 21496 36700
rect 20680 36660 20686 36672
rect 22738 36660 22744 36712
rect 22796 36700 22802 36712
rect 23293 36703 23351 36709
rect 23293 36700 23305 36703
rect 22796 36672 23305 36700
rect 22796 36660 22802 36672
rect 23293 36669 23305 36672
rect 23339 36669 23351 36703
rect 24026 36700 24032 36712
rect 23939 36672 24032 36700
rect 23293 36663 23351 36669
rect 24026 36660 24032 36672
rect 24084 36700 24090 36712
rect 25682 36700 25688 36712
rect 24084 36672 25688 36700
rect 24084 36660 24090 36672
rect 25682 36660 25688 36672
rect 25740 36660 25746 36712
rect 25774 36660 25780 36712
rect 25832 36700 25838 36712
rect 26513 36703 26571 36709
rect 26513 36700 26525 36703
rect 25832 36672 26525 36700
rect 25832 36660 25838 36672
rect 26513 36669 26525 36672
rect 26559 36669 26571 36703
rect 29638 36700 29644 36712
rect 29599 36672 29644 36700
rect 26513 36663 26571 36669
rect 29638 36660 29644 36672
rect 29696 36660 29702 36712
rect 13136 36604 14136 36632
rect 17773 36635 17831 36641
rect 13136 36592 13142 36604
rect 17773 36601 17785 36635
rect 17819 36632 17831 36635
rect 27062 36632 27068 36644
rect 17819 36604 27068 36632
rect 17819 36601 17831 36604
rect 17773 36595 17831 36601
rect 27062 36592 27068 36604
rect 27120 36592 27126 36644
rect 38010 36632 38016 36644
rect 37971 36604 38016 36632
rect 38010 36592 38016 36604
rect 38068 36592 38074 36644
rect 6328 36536 11008 36564
rect 11057 36567 11115 36573
rect 6328 36524 6334 36536
rect 11057 36533 11069 36567
rect 11103 36564 11115 36567
rect 11790 36564 11796 36576
rect 11103 36536 11796 36564
rect 11103 36533 11115 36536
rect 11057 36527 11115 36533
rect 11790 36524 11796 36536
rect 11848 36524 11854 36576
rect 12986 36524 12992 36576
rect 13044 36564 13050 36576
rect 14274 36573 14280 36576
rect 13449 36567 13507 36573
rect 13449 36564 13461 36567
rect 13044 36536 13461 36564
rect 13044 36524 13050 36536
rect 13449 36533 13461 36536
rect 13495 36533 13507 36567
rect 13449 36527 13507 36533
rect 14264 36567 14280 36573
rect 14264 36533 14276 36567
rect 14264 36527 14280 36533
rect 14274 36524 14280 36527
rect 14332 36524 14338 36576
rect 15749 36567 15807 36573
rect 15749 36533 15761 36567
rect 15795 36564 15807 36567
rect 16114 36564 16120 36576
rect 15795 36536 16120 36564
rect 15795 36533 15807 36536
rect 15749 36527 15807 36533
rect 16114 36524 16120 36536
rect 16172 36524 16178 36576
rect 16298 36564 16304 36576
rect 16259 36536 16304 36564
rect 16298 36524 16304 36536
rect 16356 36564 16362 36576
rect 16666 36564 16672 36576
rect 16356 36536 16672 36564
rect 16356 36524 16362 36536
rect 16666 36524 16672 36536
rect 16724 36524 16730 36576
rect 18598 36564 18604 36576
rect 18559 36536 18604 36564
rect 18598 36524 18604 36536
rect 18656 36524 18662 36576
rect 19150 36524 19156 36576
rect 19208 36564 19214 36576
rect 22554 36564 22560 36576
rect 19208 36536 22560 36564
rect 19208 36524 19214 36536
rect 22554 36524 22560 36536
rect 22612 36524 22618 36576
rect 22741 36567 22799 36573
rect 22741 36533 22753 36567
rect 22787 36564 22799 36567
rect 22830 36564 22836 36576
rect 22787 36536 22836 36564
rect 22787 36533 22799 36536
rect 22741 36527 22799 36533
rect 22830 36524 22836 36536
rect 22888 36524 22894 36576
rect 24670 36564 24676 36576
rect 24631 36536 24676 36564
rect 24670 36524 24676 36536
rect 24728 36564 24734 36576
rect 25133 36567 25191 36573
rect 25133 36564 25145 36567
rect 24728 36536 25145 36564
rect 24728 36524 24734 36536
rect 25133 36533 25145 36536
rect 25179 36533 25191 36567
rect 25133 36527 25191 36533
rect 28077 36567 28135 36573
rect 28077 36533 28089 36567
rect 28123 36564 28135 36567
rect 28442 36564 28448 36576
rect 28123 36536 28448 36564
rect 28123 36533 28135 36536
rect 28077 36527 28135 36533
rect 28442 36524 28448 36536
rect 28500 36564 28506 36576
rect 28537 36567 28595 36573
rect 28537 36564 28549 36567
rect 28500 36536 28549 36564
rect 28500 36524 28506 36536
rect 28537 36533 28549 36536
rect 28583 36564 28595 36567
rect 29089 36567 29147 36573
rect 29089 36564 29101 36567
rect 28583 36536 29101 36564
rect 28583 36533 28595 36536
rect 28537 36527 28595 36533
rect 29089 36533 29101 36536
rect 29135 36533 29147 36567
rect 29089 36527 29147 36533
rect 37458 36524 37464 36576
rect 37516 36564 37522 36576
rect 37553 36567 37611 36573
rect 37553 36564 37565 36567
rect 37516 36536 37565 36564
rect 37516 36524 37522 36536
rect 37553 36533 37565 36536
rect 37599 36564 37611 36567
rect 37918 36564 37924 36576
rect 37599 36536 37924 36564
rect 37599 36533 37611 36536
rect 37553 36527 37611 36533
rect 37918 36524 37924 36536
rect 37976 36524 37982 36576
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 4065 36363 4123 36369
rect 4065 36329 4077 36363
rect 4111 36360 4123 36363
rect 4614 36360 4620 36372
rect 4111 36332 4620 36360
rect 4111 36329 4123 36332
rect 4065 36323 4123 36329
rect 4614 36320 4620 36332
rect 4672 36320 4678 36372
rect 6365 36363 6423 36369
rect 4724 36332 6316 36360
rect 3421 36295 3479 36301
rect 3421 36261 3433 36295
rect 3467 36292 3479 36295
rect 4724 36292 4752 36332
rect 3467 36264 4752 36292
rect 6288 36292 6316 36332
rect 6365 36329 6377 36363
rect 6411 36360 6423 36363
rect 7190 36360 7196 36372
rect 6411 36332 7196 36360
rect 6411 36329 6423 36332
rect 6365 36323 6423 36329
rect 7190 36320 7196 36332
rect 7248 36320 7254 36372
rect 8573 36363 8631 36369
rect 8573 36329 8585 36363
rect 8619 36360 8631 36363
rect 8619 36332 11468 36360
rect 8619 36329 8631 36332
rect 8573 36323 8631 36329
rect 6288 36264 6960 36292
rect 3467 36261 3479 36264
rect 3421 36255 3479 36261
rect 1949 36227 2007 36233
rect 1949 36193 1961 36227
rect 1995 36224 2007 36227
rect 3694 36224 3700 36236
rect 1995 36196 3700 36224
rect 1995 36193 2007 36196
rect 1949 36187 2007 36193
rect 3694 36184 3700 36196
rect 3752 36184 3758 36236
rect 3878 36184 3884 36236
rect 3936 36224 3942 36236
rect 4617 36227 4675 36233
rect 4617 36224 4629 36227
rect 3936 36196 4629 36224
rect 3936 36184 3942 36196
rect 4617 36193 4629 36196
rect 4663 36224 4675 36227
rect 6822 36224 6828 36236
rect 4663 36196 6828 36224
rect 4663 36193 4675 36196
rect 4617 36187 4675 36193
rect 6822 36184 6828 36196
rect 6880 36184 6886 36236
rect 6932 36224 6960 36264
rect 7742 36224 7748 36236
rect 6932 36196 7748 36224
rect 7742 36184 7748 36196
rect 7800 36224 7806 36236
rect 9401 36227 9459 36233
rect 7800 36196 8432 36224
rect 7800 36184 7806 36196
rect 1670 36156 1676 36168
rect 1631 36128 1676 36156
rect 1670 36116 1676 36128
rect 1728 36116 1734 36168
rect 3970 36156 3976 36168
rect 3931 36128 3976 36156
rect 3970 36116 3976 36128
rect 4028 36116 4034 36168
rect 8202 36116 8208 36168
rect 8260 36116 8266 36168
rect 2958 36048 2964 36100
rect 3016 36048 3022 36100
rect 4893 36091 4951 36097
rect 4893 36057 4905 36091
rect 4939 36088 4951 36091
rect 4982 36088 4988 36100
rect 4939 36060 4988 36088
rect 4939 36057 4951 36060
rect 4893 36051 4951 36057
rect 4982 36048 4988 36060
rect 5040 36048 5046 36100
rect 7101 36091 7159 36097
rect 6118 36060 7052 36088
rect 4062 35980 4068 36032
rect 4120 36020 4126 36032
rect 6914 36020 6920 36032
rect 4120 35992 6920 36020
rect 4120 35980 4126 35992
rect 6914 35980 6920 35992
rect 6972 35980 6978 36032
rect 7024 36020 7052 36060
rect 7101 36057 7113 36091
rect 7147 36088 7159 36091
rect 7190 36088 7196 36100
rect 7147 36060 7196 36088
rect 7147 36057 7159 36060
rect 7101 36051 7159 36057
rect 7190 36048 7196 36060
rect 7248 36048 7254 36100
rect 8404 36088 8432 36196
rect 9401 36193 9413 36227
rect 9447 36224 9459 36227
rect 10962 36224 10968 36236
rect 9447 36196 10968 36224
rect 9447 36193 9459 36196
rect 9401 36187 9459 36193
rect 10962 36184 10968 36196
rect 11020 36184 11026 36236
rect 11440 36224 11468 36332
rect 11606 36320 11612 36372
rect 11664 36360 11670 36372
rect 13722 36360 13728 36372
rect 11664 36332 13728 36360
rect 11664 36320 11670 36332
rect 13722 36320 13728 36332
rect 13780 36320 13786 36372
rect 17405 36363 17463 36369
rect 14752 36332 16988 36360
rect 12710 36252 12716 36304
rect 12768 36292 12774 36304
rect 14752 36292 14780 36332
rect 12768 36264 14780 36292
rect 12768 36252 12774 36264
rect 11606 36224 11612 36236
rect 11440 36196 11612 36224
rect 11606 36184 11612 36196
rect 11664 36184 11670 36236
rect 12618 36184 12624 36236
rect 12676 36224 12682 36236
rect 13078 36224 13084 36236
rect 12676 36196 13084 36224
rect 12676 36184 12682 36196
rect 13078 36184 13084 36196
rect 13136 36184 13142 36236
rect 14274 36184 14280 36236
rect 14332 36224 14338 36236
rect 16025 36227 16083 36233
rect 16025 36224 16037 36227
rect 14332 36196 16037 36224
rect 14332 36184 14338 36196
rect 16025 36193 16037 36196
rect 16071 36193 16083 36227
rect 16960 36224 16988 36332
rect 17405 36329 17417 36363
rect 17451 36360 17463 36363
rect 19426 36360 19432 36372
rect 17451 36332 19432 36360
rect 17451 36329 17463 36332
rect 17405 36323 17463 36329
rect 19426 36320 19432 36332
rect 19484 36320 19490 36372
rect 23014 36360 23020 36372
rect 21560 36332 23020 36360
rect 17034 36252 17040 36304
rect 17092 36292 17098 36304
rect 19521 36295 19579 36301
rect 19521 36292 19533 36295
rect 17092 36264 19533 36292
rect 17092 36252 17098 36264
rect 19521 36261 19533 36264
rect 19567 36261 19579 36295
rect 20714 36292 20720 36304
rect 19521 36255 19579 36261
rect 19628 36264 20720 36292
rect 18785 36227 18843 36233
rect 18785 36224 18797 36227
rect 16960 36196 18797 36224
rect 16025 36187 16083 36193
rect 18785 36193 18797 36196
rect 18831 36193 18843 36227
rect 18785 36187 18843 36193
rect 19058 36184 19064 36236
rect 19116 36224 19122 36236
rect 19628 36224 19656 36264
rect 20714 36252 20720 36264
rect 20772 36252 20778 36304
rect 21560 36224 21588 36332
rect 23014 36320 23020 36332
rect 23072 36320 23078 36372
rect 23842 36360 23848 36372
rect 23803 36332 23848 36360
rect 23842 36320 23848 36332
rect 23900 36320 23906 36372
rect 37182 36320 37188 36372
rect 37240 36360 37246 36372
rect 37369 36363 37427 36369
rect 37369 36360 37381 36363
rect 37240 36332 37381 36360
rect 37240 36320 37246 36332
rect 37369 36329 37381 36332
rect 37415 36329 37427 36363
rect 37369 36323 37427 36329
rect 38197 36363 38255 36369
rect 38197 36329 38209 36363
rect 38243 36360 38255 36363
rect 38286 36360 38292 36372
rect 38243 36332 38292 36360
rect 38243 36329 38255 36332
rect 38197 36323 38255 36329
rect 38286 36320 38292 36332
rect 38344 36320 38350 36372
rect 21634 36252 21640 36304
rect 21692 36292 21698 36304
rect 26789 36295 26847 36301
rect 26789 36292 26801 36295
rect 21692 36264 26801 36292
rect 21692 36252 21698 36264
rect 26789 36261 26801 36264
rect 26835 36261 26847 36295
rect 26789 36255 26847 36261
rect 22097 36227 22155 36233
rect 22097 36224 22109 36227
rect 19116 36196 19656 36224
rect 19996 36196 22109 36224
rect 19116 36184 19122 36196
rect 8570 36116 8576 36168
rect 8628 36156 8634 36168
rect 9122 36156 9128 36168
rect 8628 36128 9128 36156
rect 8628 36116 8634 36128
rect 9122 36116 9128 36128
rect 9180 36116 9186 36168
rect 11054 36116 11060 36168
rect 11112 36156 11118 36168
rect 11333 36159 11391 36165
rect 11333 36156 11345 36159
rect 11112 36128 11345 36156
rect 11112 36116 11118 36128
rect 11333 36125 11345 36128
rect 11379 36125 11391 36159
rect 11333 36119 11391 36125
rect 13725 36159 13783 36165
rect 13725 36125 13737 36159
rect 13771 36156 13783 36159
rect 16577 36159 16635 36165
rect 13771 36128 14504 36156
rect 13771 36125 13783 36128
rect 13725 36119 13783 36125
rect 9490 36088 9496 36100
rect 8404 36060 9496 36088
rect 9490 36048 9496 36060
rect 9548 36048 9554 36100
rect 11882 36088 11888 36100
rect 10626 36060 11888 36088
rect 11882 36048 11888 36060
rect 11940 36048 11946 36100
rect 13446 36088 13452 36100
rect 12834 36060 13452 36088
rect 13446 36048 13452 36060
rect 13504 36048 13510 36100
rect 10686 36020 10692 36032
rect 7024 35992 10692 36020
rect 10686 35980 10692 35992
rect 10744 35980 10750 36032
rect 10870 36020 10876 36032
rect 10831 35992 10876 36020
rect 10870 35980 10876 35992
rect 10928 35980 10934 36032
rect 10962 35980 10968 36032
rect 11020 36020 11026 36032
rect 13170 36020 13176 36032
rect 11020 35992 13176 36020
rect 11020 35980 11026 35992
rect 13170 35980 13176 35992
rect 13228 35980 13234 36032
rect 13262 35980 13268 36032
rect 13320 36020 13326 36032
rect 13541 36023 13599 36029
rect 13541 36020 13553 36023
rect 13320 35992 13553 36020
rect 13320 35980 13326 35992
rect 13541 35989 13553 35992
rect 13587 35989 13599 36023
rect 13541 35983 13599 35989
rect 13906 35980 13912 36032
rect 13964 36020 13970 36032
rect 14277 36023 14335 36029
rect 14277 36020 14289 36023
rect 13964 35992 14289 36020
rect 13964 35980 13970 35992
rect 14277 35989 14289 35992
rect 14323 35989 14335 36023
rect 14476 36020 14504 36128
rect 16577 36125 16589 36159
rect 16623 36156 16635 36159
rect 16758 36156 16764 36168
rect 16623 36128 16764 36156
rect 16623 36125 16635 36128
rect 16577 36119 16635 36125
rect 16758 36116 16764 36128
rect 16816 36116 16822 36168
rect 17218 36156 17224 36168
rect 17179 36128 17224 36156
rect 17218 36116 17224 36128
rect 17276 36116 17282 36168
rect 17862 36156 17868 36168
rect 17823 36128 17868 36156
rect 17862 36116 17868 36128
rect 17920 36116 17926 36168
rect 18877 36159 18935 36165
rect 18877 36125 18889 36159
rect 18923 36152 18935 36159
rect 18966 36152 18972 36168
rect 18923 36125 18972 36152
rect 18877 36124 18972 36125
rect 18877 36119 18935 36124
rect 18966 36116 18972 36124
rect 19024 36156 19030 36168
rect 19613 36159 19671 36165
rect 19613 36156 19625 36159
rect 19024 36128 19625 36156
rect 19024 36116 19030 36128
rect 19613 36125 19625 36128
rect 19659 36125 19671 36159
rect 19613 36119 19671 36125
rect 15102 36048 15108 36100
rect 15160 36048 15166 36100
rect 15746 36088 15752 36100
rect 15707 36060 15752 36088
rect 15746 36048 15752 36060
rect 15804 36048 15810 36100
rect 18782 36048 18788 36100
rect 18840 36088 18846 36100
rect 19996 36088 20024 36196
rect 22097 36193 22109 36196
rect 22143 36193 22155 36227
rect 22738 36224 22744 36236
rect 22699 36196 22744 36224
rect 22097 36187 22155 36193
rect 22738 36184 22744 36196
rect 22796 36184 22802 36236
rect 20073 36159 20131 36165
rect 20073 36125 20085 36159
rect 20119 36156 20131 36159
rect 20438 36156 20444 36168
rect 20119 36128 20444 36156
rect 20119 36125 20131 36128
rect 20073 36119 20131 36125
rect 20438 36116 20444 36128
rect 20496 36116 20502 36168
rect 20622 36116 20628 36168
rect 20680 36156 20686 36168
rect 21637 36159 21695 36165
rect 21637 36156 21649 36159
rect 20680 36128 21649 36156
rect 20680 36116 20686 36128
rect 21637 36125 21649 36128
rect 21683 36125 21695 36159
rect 21637 36119 21695 36125
rect 37553 36159 37611 36165
rect 37553 36125 37565 36159
rect 37599 36156 37611 36159
rect 37826 36156 37832 36168
rect 37599 36128 37832 36156
rect 37599 36125 37611 36128
rect 37553 36119 37611 36125
rect 37826 36116 37832 36128
rect 37884 36116 37890 36168
rect 37918 36116 37924 36168
rect 37976 36156 37982 36168
rect 38013 36159 38071 36165
rect 38013 36156 38025 36159
rect 37976 36128 38025 36156
rect 37976 36116 37982 36128
rect 38013 36125 38025 36128
rect 38059 36125 38071 36159
rect 38013 36119 38071 36125
rect 18840 36060 20024 36088
rect 20349 36091 20407 36097
rect 18840 36048 18846 36060
rect 20349 36057 20361 36091
rect 20395 36088 20407 36091
rect 20640 36088 20668 36116
rect 20395 36060 20668 36088
rect 20395 36057 20407 36060
rect 20349 36051 20407 36057
rect 20714 36048 20720 36100
rect 20772 36088 20778 36100
rect 22646 36088 22652 36100
rect 20772 36060 22094 36088
rect 22607 36060 22652 36088
rect 20772 36048 20778 36060
rect 16574 36020 16580 36032
rect 14476 35992 16580 36020
rect 14277 35983 14335 35989
rect 16574 35980 16580 35992
rect 16632 35980 16638 36032
rect 16669 36023 16727 36029
rect 16669 35989 16681 36023
rect 16715 36020 16727 36023
rect 17402 36020 17408 36032
rect 16715 35992 17408 36020
rect 16715 35989 16727 35992
rect 16669 35983 16727 35989
rect 17402 35980 17408 35992
rect 17460 35980 17466 36032
rect 17954 36020 17960 36032
rect 17915 35992 17960 36020
rect 17954 35980 17960 35992
rect 18012 35980 18018 36032
rect 18046 35980 18052 36032
rect 18104 36020 18110 36032
rect 21545 36023 21603 36029
rect 21545 36020 21557 36023
rect 18104 35992 21557 36020
rect 18104 35980 18110 35992
rect 21545 35989 21557 35992
rect 21591 35989 21603 36023
rect 22066 36020 22094 36060
rect 22646 36048 22652 36060
rect 22704 36048 22710 36100
rect 23293 36023 23351 36029
rect 23293 36020 23305 36023
rect 22066 35992 23305 36020
rect 21545 35983 21603 35989
rect 23293 35989 23305 35992
rect 23339 35989 23351 36023
rect 24670 36020 24676 36032
rect 24631 35992 24676 36020
rect 23293 35983 23351 35989
rect 24670 35980 24676 35992
rect 24728 36020 24734 36032
rect 25133 36023 25191 36029
rect 25133 36020 25145 36023
rect 24728 35992 25145 36020
rect 24728 35980 24734 35992
rect 25133 35989 25145 35992
rect 25179 36020 25191 36023
rect 25685 36023 25743 36029
rect 25685 36020 25697 36023
rect 25179 35992 25697 36020
rect 25179 35989 25191 35992
rect 25133 35983 25191 35989
rect 25685 35989 25697 35992
rect 25731 36020 25743 36023
rect 26237 36023 26295 36029
rect 26237 36020 26249 36023
rect 25731 35992 26249 36020
rect 25731 35989 25743 35992
rect 25685 35983 25743 35989
rect 26237 35989 26249 35992
rect 26283 35989 26295 36023
rect 27338 36020 27344 36032
rect 27299 35992 27344 36020
rect 26237 35983 26295 35989
rect 27338 35980 27344 35992
rect 27396 35980 27402 36032
rect 27890 36020 27896 36032
rect 27851 35992 27896 36020
rect 27890 35980 27896 35992
rect 27948 35980 27954 36032
rect 28442 36020 28448 36032
rect 28403 35992 28448 36020
rect 28442 35980 28448 35992
rect 28500 35980 28506 36032
rect 28994 36020 29000 36032
rect 28955 35992 29000 36020
rect 28994 35980 29000 35992
rect 29052 35980 29058 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 3878 35776 3884 35828
rect 3936 35816 3942 35828
rect 6917 35819 6975 35825
rect 3936 35788 6040 35816
rect 3936 35776 3942 35788
rect 1302 35708 1308 35760
rect 1360 35748 1366 35760
rect 1360 35720 2806 35748
rect 1360 35708 1366 35720
rect 5258 35708 5264 35760
rect 5316 35708 5322 35760
rect 5718 35748 5724 35760
rect 5679 35720 5724 35748
rect 5718 35708 5724 35720
rect 5776 35708 5782 35760
rect 1670 35640 1676 35692
rect 1728 35680 1734 35692
rect 6012 35689 6040 35788
rect 6917 35785 6929 35819
rect 6963 35816 6975 35819
rect 8386 35816 8392 35828
rect 6963 35788 8392 35816
rect 6963 35785 6975 35788
rect 6917 35779 6975 35785
rect 8386 35776 8392 35788
rect 8444 35776 8450 35828
rect 9122 35776 9128 35828
rect 9180 35776 9186 35828
rect 9214 35776 9220 35828
rect 9272 35816 9278 35828
rect 9766 35816 9772 35828
rect 9272 35788 9772 35816
rect 9272 35776 9278 35788
rect 9766 35776 9772 35788
rect 9824 35776 9830 35828
rect 10318 35776 10324 35828
rect 10376 35816 10382 35828
rect 10505 35819 10563 35825
rect 10505 35816 10517 35819
rect 10376 35788 10517 35816
rect 10376 35776 10382 35788
rect 10505 35785 10517 35788
rect 10551 35785 10563 35819
rect 10505 35779 10563 35785
rect 11606 35776 11612 35828
rect 11664 35816 11670 35828
rect 18785 35819 18843 35825
rect 11664 35788 18000 35816
rect 11664 35776 11670 35788
rect 8846 35708 8852 35760
rect 8904 35708 8910 35760
rect 9140 35748 9168 35776
rect 9140 35720 9628 35748
rect 2041 35683 2099 35689
rect 2041 35680 2053 35683
rect 1728 35652 2053 35680
rect 1728 35640 1734 35652
rect 2041 35649 2053 35652
rect 2087 35649 2099 35683
rect 2041 35643 2099 35649
rect 5997 35683 6055 35689
rect 5997 35649 6009 35683
rect 6043 35649 6055 35683
rect 7098 35680 7104 35692
rect 7059 35652 7104 35680
rect 5997 35643 6055 35649
rect 7098 35640 7104 35652
rect 7156 35640 7162 35692
rect 9600 35689 9628 35720
rect 10870 35708 10876 35760
rect 10928 35748 10934 35760
rect 11977 35751 12035 35757
rect 11977 35748 11989 35751
rect 10928 35720 11989 35748
rect 10928 35708 10934 35720
rect 11977 35717 11989 35720
rect 12023 35717 12035 35751
rect 11977 35711 12035 35717
rect 14918 35708 14924 35760
rect 14976 35708 14982 35760
rect 15102 35708 15108 35760
rect 15160 35748 15166 35760
rect 15381 35751 15439 35757
rect 15381 35748 15393 35751
rect 15160 35720 15393 35748
rect 15160 35708 15166 35720
rect 15381 35717 15393 35720
rect 15427 35717 15439 35751
rect 15381 35711 15439 35717
rect 15470 35708 15476 35760
rect 15528 35748 15534 35760
rect 16209 35751 16267 35757
rect 16209 35748 16221 35751
rect 15528 35720 16221 35748
rect 15528 35708 15534 35720
rect 16209 35717 16221 35720
rect 16255 35717 16267 35751
rect 16209 35711 16267 35717
rect 9585 35683 9643 35689
rect 9585 35649 9597 35683
rect 9631 35649 9643 35683
rect 9585 35643 9643 35649
rect 10689 35683 10747 35689
rect 10689 35649 10701 35683
rect 10735 35680 10747 35683
rect 10778 35680 10784 35692
rect 10735 35652 10784 35680
rect 10735 35649 10747 35652
rect 10689 35643 10747 35649
rect 10778 35640 10784 35652
rect 10836 35640 10842 35692
rect 14090 35680 14096 35692
rect 13110 35652 14096 35680
rect 14090 35640 14096 35652
rect 14148 35640 14154 35692
rect 16301 35683 16359 35689
rect 16301 35649 16313 35683
rect 16347 35680 16359 35683
rect 16390 35680 16396 35692
rect 16347 35652 16396 35680
rect 16347 35649 16359 35652
rect 16301 35643 16359 35649
rect 16390 35640 16396 35652
rect 16448 35640 16454 35692
rect 16666 35640 16672 35692
rect 16724 35680 16730 35692
rect 16942 35680 16948 35692
rect 16724 35652 16948 35680
rect 16724 35640 16730 35652
rect 16942 35640 16948 35652
rect 17000 35680 17006 35692
rect 17972 35689 18000 35788
rect 18785 35785 18797 35819
rect 18831 35816 18843 35819
rect 19978 35816 19984 35828
rect 18831 35788 19984 35816
rect 18831 35785 18843 35788
rect 18785 35779 18843 35785
rect 19978 35776 19984 35788
rect 20036 35776 20042 35828
rect 19426 35708 19432 35760
rect 19484 35748 19490 35760
rect 19613 35751 19671 35757
rect 19613 35748 19625 35751
rect 19484 35720 19625 35748
rect 19484 35708 19490 35720
rect 19613 35717 19625 35720
rect 19659 35717 19671 35751
rect 19613 35711 19671 35717
rect 19794 35708 19800 35760
rect 19852 35748 19858 35760
rect 20070 35748 20076 35760
rect 19852 35720 20076 35748
rect 19852 35708 19858 35720
rect 20070 35708 20076 35720
rect 20128 35748 20134 35760
rect 27154 35748 27160 35760
rect 20128 35720 22232 35748
rect 27115 35720 27160 35748
rect 20128 35708 20134 35720
rect 17037 35683 17095 35689
rect 17037 35680 17049 35683
rect 17000 35652 17049 35680
rect 17000 35640 17006 35652
rect 17037 35649 17049 35652
rect 17083 35649 17095 35683
rect 17037 35643 17095 35649
rect 17957 35683 18015 35689
rect 17957 35649 17969 35683
rect 18003 35649 18015 35683
rect 17957 35643 18015 35649
rect 18601 35683 18659 35689
rect 18601 35649 18613 35683
rect 18647 35649 18659 35683
rect 18601 35643 18659 35649
rect 19705 35683 19763 35689
rect 19705 35649 19717 35683
rect 19751 35680 19763 35683
rect 19978 35680 19984 35692
rect 19751 35652 19984 35680
rect 19751 35649 19763 35652
rect 19705 35643 19763 35649
rect 2317 35615 2375 35621
rect 2317 35581 2329 35615
rect 2363 35612 2375 35615
rect 2406 35612 2412 35624
rect 2363 35584 2412 35612
rect 2363 35581 2375 35584
rect 2317 35575 2375 35581
rect 2406 35572 2412 35584
rect 2464 35572 2470 35624
rect 4982 35572 4988 35624
rect 5040 35612 5046 35624
rect 7561 35615 7619 35621
rect 5040 35584 5948 35612
rect 5040 35572 5046 35584
rect 3789 35547 3847 35553
rect 3789 35513 3801 35547
rect 3835 35544 3847 35547
rect 4706 35544 4712 35556
rect 3835 35516 4712 35544
rect 3835 35513 3847 35516
rect 3789 35507 3847 35513
rect 4706 35504 4712 35516
rect 4764 35504 4770 35556
rect 5920 35544 5948 35584
rect 7561 35581 7573 35615
rect 7607 35612 7619 35615
rect 9214 35612 9220 35624
rect 7607 35584 9220 35612
rect 7607 35581 7619 35584
rect 7561 35575 7619 35581
rect 9214 35572 9220 35584
rect 9272 35572 9278 35624
rect 9309 35615 9367 35621
rect 9309 35581 9321 35615
rect 9355 35612 9367 35615
rect 9355 35584 9674 35612
rect 9355 35581 9367 35584
rect 9309 35575 9367 35581
rect 8294 35544 8300 35556
rect 5920 35516 8300 35544
rect 8294 35504 8300 35516
rect 8352 35504 8358 35556
rect 9646 35544 9674 35584
rect 11054 35572 11060 35624
rect 11112 35612 11118 35624
rect 11701 35615 11759 35621
rect 11701 35612 11713 35615
rect 11112 35584 11713 35612
rect 11112 35572 11118 35584
rect 11701 35581 11713 35584
rect 11747 35581 11759 35615
rect 12618 35612 12624 35624
rect 11701 35575 11759 35581
rect 11808 35584 12624 35612
rect 11808 35544 11836 35584
rect 12618 35572 12624 35584
rect 12676 35572 12682 35624
rect 13814 35572 13820 35624
rect 13872 35612 13878 35624
rect 13909 35615 13967 35621
rect 13909 35612 13921 35615
rect 13872 35584 13921 35612
rect 13872 35572 13878 35584
rect 13909 35581 13921 35584
rect 13955 35581 13967 35615
rect 13909 35575 13967 35581
rect 15657 35615 15715 35621
rect 15657 35581 15669 35615
rect 15703 35581 15715 35615
rect 15657 35575 15715 35581
rect 9646 35516 11836 35544
rect 13078 35504 13084 35556
rect 13136 35544 13142 35556
rect 14366 35544 14372 35556
rect 13136 35516 14372 35544
rect 13136 35504 13142 35516
rect 14366 35504 14372 35516
rect 14424 35504 14430 35556
rect 3694 35436 3700 35488
rect 3752 35476 3758 35488
rect 4249 35479 4307 35485
rect 4249 35476 4261 35479
rect 3752 35448 4261 35476
rect 3752 35436 3758 35448
rect 4249 35445 4261 35448
rect 4295 35476 4307 35479
rect 6454 35476 6460 35488
rect 4295 35448 6460 35476
rect 4295 35445 4307 35448
rect 4249 35439 4307 35445
rect 6454 35436 6460 35448
rect 6512 35436 6518 35488
rect 7190 35436 7196 35488
rect 7248 35476 7254 35488
rect 10594 35476 10600 35488
rect 7248 35448 10600 35476
rect 7248 35436 7254 35448
rect 10594 35436 10600 35448
rect 10652 35436 10658 35488
rect 13449 35479 13507 35485
rect 13449 35445 13461 35479
rect 13495 35476 13507 35479
rect 13630 35476 13636 35488
rect 13495 35448 13636 35476
rect 13495 35445 13507 35448
rect 13449 35439 13507 35445
rect 13630 35436 13636 35448
rect 13688 35436 13694 35488
rect 14274 35436 14280 35488
rect 14332 35476 14338 35488
rect 15672 35476 15700 35575
rect 16574 35572 16580 35624
rect 16632 35612 16638 35624
rect 18616 35612 18644 35643
rect 19978 35640 19984 35652
rect 20036 35680 20042 35692
rect 20162 35680 20168 35692
rect 20036 35652 20168 35680
rect 20036 35640 20042 35652
rect 20162 35640 20168 35652
rect 20220 35680 20226 35692
rect 20349 35683 20407 35689
rect 20349 35680 20361 35683
rect 20220 35652 20361 35680
rect 20220 35640 20226 35652
rect 20349 35649 20361 35652
rect 20395 35649 20407 35683
rect 20349 35643 20407 35649
rect 20806 35640 20812 35692
rect 20864 35680 20870 35692
rect 22204 35689 22232 35720
rect 27154 35708 27160 35720
rect 27212 35708 27218 35760
rect 20993 35683 21051 35689
rect 20993 35680 21005 35683
rect 20864 35652 21005 35680
rect 20864 35640 20870 35652
rect 20993 35649 21005 35652
rect 21039 35649 21051 35683
rect 20993 35643 21051 35649
rect 22189 35683 22247 35689
rect 22189 35649 22201 35683
rect 22235 35680 22247 35683
rect 22738 35680 22744 35692
rect 22235 35652 22744 35680
rect 22235 35649 22247 35652
rect 22189 35643 22247 35649
rect 22738 35640 22744 35652
rect 22796 35640 22802 35692
rect 22830 35640 22836 35692
rect 22888 35680 22894 35692
rect 30558 35680 30564 35692
rect 22888 35652 30564 35680
rect 22888 35640 22894 35652
rect 30558 35640 30564 35652
rect 30616 35640 30622 35692
rect 38013 35683 38071 35689
rect 38013 35680 38025 35683
rect 37476 35652 38025 35680
rect 16632 35584 18644 35612
rect 16632 35572 16638 35584
rect 18874 35572 18880 35624
rect 18932 35612 18938 35624
rect 20901 35615 20959 35621
rect 20901 35612 20913 35615
rect 18932 35584 20913 35612
rect 18932 35572 18938 35584
rect 20901 35581 20913 35584
rect 20947 35581 20959 35615
rect 23198 35612 23204 35624
rect 23159 35584 23204 35612
rect 20901 35575 20959 35581
rect 23198 35572 23204 35584
rect 23256 35572 23262 35624
rect 16758 35504 16764 35556
rect 16816 35544 16822 35556
rect 22370 35544 22376 35556
rect 16816 35516 22376 35544
rect 16816 35504 16822 35516
rect 22370 35504 22376 35516
rect 22428 35504 22434 35556
rect 27709 35547 27767 35553
rect 27709 35544 27721 35547
rect 26528 35516 27721 35544
rect 14332 35448 15700 35476
rect 16945 35479 17003 35485
rect 14332 35436 14338 35448
rect 16945 35445 16957 35479
rect 16991 35476 17003 35479
rect 17034 35476 17040 35488
rect 16991 35448 17040 35476
rect 16991 35445 17003 35448
rect 16945 35439 17003 35445
rect 17034 35436 17040 35448
rect 17092 35436 17098 35488
rect 18049 35479 18107 35485
rect 18049 35445 18061 35479
rect 18095 35476 18107 35479
rect 18230 35476 18236 35488
rect 18095 35448 18236 35476
rect 18095 35445 18107 35448
rect 18049 35439 18107 35445
rect 18230 35436 18236 35448
rect 18288 35436 18294 35488
rect 20254 35476 20260 35488
rect 20215 35448 20260 35476
rect 20254 35436 20260 35448
rect 20312 35436 20318 35488
rect 22094 35436 22100 35488
rect 22152 35476 22158 35488
rect 22738 35476 22744 35488
rect 22152 35448 22197 35476
rect 22699 35448 22744 35476
rect 22152 35436 22158 35448
rect 22738 35436 22744 35448
rect 22796 35436 22802 35488
rect 23750 35476 23756 35488
rect 23711 35448 23756 35476
rect 23750 35436 23756 35448
rect 23808 35436 23814 35488
rect 24026 35436 24032 35488
rect 24084 35476 24090 35488
rect 24305 35479 24363 35485
rect 24305 35476 24317 35479
rect 24084 35448 24317 35476
rect 24084 35436 24090 35448
rect 24305 35445 24317 35448
rect 24351 35476 24363 35479
rect 24670 35476 24676 35488
rect 24351 35448 24676 35476
rect 24351 35445 24363 35448
rect 24305 35439 24363 35445
rect 24670 35436 24676 35448
rect 24728 35476 24734 35488
rect 24857 35479 24915 35485
rect 24857 35476 24869 35479
rect 24728 35448 24869 35476
rect 24728 35436 24734 35448
rect 24857 35445 24869 35448
rect 24903 35476 24915 35479
rect 25409 35479 25467 35485
rect 25409 35476 25421 35479
rect 24903 35448 25421 35476
rect 24903 35445 24915 35448
rect 24857 35439 24915 35445
rect 25409 35445 25421 35448
rect 25455 35476 25467 35479
rect 25961 35479 26019 35485
rect 25961 35476 25973 35479
rect 25455 35448 25973 35476
rect 25455 35445 25467 35448
rect 25409 35439 25467 35445
rect 25961 35445 25973 35448
rect 26007 35476 26019 35479
rect 26234 35476 26240 35488
rect 26007 35448 26240 35476
rect 26007 35445 26019 35448
rect 25961 35439 26019 35445
rect 26234 35436 26240 35448
rect 26292 35476 26298 35488
rect 26528 35485 26556 35516
rect 27709 35513 27721 35516
rect 27755 35544 27767 35547
rect 28261 35547 28319 35553
rect 28261 35544 28273 35547
rect 27755 35516 28273 35544
rect 27755 35513 27767 35516
rect 27709 35507 27767 35513
rect 28261 35513 28273 35516
rect 28307 35544 28319 35547
rect 28442 35544 28448 35556
rect 28307 35516 28448 35544
rect 28307 35513 28319 35516
rect 28261 35507 28319 35513
rect 28442 35504 28448 35516
rect 28500 35544 28506 35556
rect 28813 35547 28871 35553
rect 28813 35544 28825 35547
rect 28500 35516 28825 35544
rect 28500 35504 28506 35516
rect 28813 35513 28825 35516
rect 28859 35513 28871 35547
rect 28813 35507 28871 35513
rect 26513 35479 26571 35485
rect 26513 35476 26525 35479
rect 26292 35448 26525 35476
rect 26292 35436 26298 35448
rect 26513 35445 26525 35448
rect 26559 35445 26571 35479
rect 26513 35439 26571 35445
rect 27982 35436 27988 35488
rect 28040 35476 28046 35488
rect 37476 35485 37504 35652
rect 38013 35649 38025 35652
rect 38059 35649 38071 35683
rect 38013 35643 38071 35649
rect 37461 35479 37519 35485
rect 37461 35476 37473 35479
rect 28040 35448 37473 35476
rect 28040 35436 28046 35448
rect 37461 35445 37473 35448
rect 37507 35445 37519 35479
rect 38194 35476 38200 35488
rect 38155 35448 38200 35476
rect 37461 35439 37519 35445
rect 38194 35436 38200 35448
rect 38252 35436 38258 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 3970 35232 3976 35284
rect 4028 35272 4034 35284
rect 6825 35275 6883 35281
rect 4028 35244 6776 35272
rect 4028 35232 4034 35244
rect 3786 35164 3792 35216
rect 3844 35204 3850 35216
rect 6748 35204 6776 35244
rect 6825 35241 6837 35275
rect 6871 35272 6883 35275
rect 7190 35272 7196 35284
rect 6871 35244 7196 35272
rect 6871 35241 6883 35244
rect 6825 35235 6883 35241
rect 7190 35232 7196 35244
rect 7248 35232 7254 35284
rect 7650 35272 7656 35284
rect 7300 35244 7656 35272
rect 7300 35204 7328 35244
rect 7650 35232 7656 35244
rect 7708 35232 7714 35284
rect 7834 35232 7840 35284
rect 7892 35272 7898 35284
rect 13078 35272 13084 35284
rect 7892 35244 13084 35272
rect 7892 35232 7898 35244
rect 13078 35232 13084 35244
rect 13136 35232 13142 35284
rect 14182 35232 14188 35284
rect 14240 35272 14246 35284
rect 19794 35272 19800 35284
rect 14240 35244 19800 35272
rect 14240 35232 14246 35244
rect 19794 35232 19800 35244
rect 19852 35232 19858 35284
rect 24581 35275 24639 35281
rect 24581 35272 24593 35275
rect 21284 35244 24593 35272
rect 9398 35204 9404 35216
rect 3844 35176 4752 35204
rect 6748 35176 7328 35204
rect 8496 35176 9404 35204
rect 3844 35164 3850 35176
rect 3418 35136 3424 35148
rect 3331 35108 3424 35136
rect 3418 35096 3424 35108
rect 3476 35136 3482 35148
rect 3878 35136 3884 35148
rect 3476 35108 3884 35136
rect 3476 35096 3482 35108
rect 3878 35096 3884 35108
rect 3936 35136 3942 35148
rect 4617 35139 4675 35145
rect 4617 35136 4629 35139
rect 3936 35108 4629 35136
rect 3936 35096 3942 35108
rect 4617 35105 4629 35108
rect 4663 35105 4675 35139
rect 4724 35136 4752 35176
rect 8496 35136 8524 35176
rect 9398 35164 9404 35176
rect 9456 35164 9462 35216
rect 14366 35164 14372 35216
rect 14424 35204 14430 35216
rect 18785 35207 18843 35213
rect 18785 35204 18797 35207
rect 14424 35176 18797 35204
rect 14424 35164 14430 35176
rect 18785 35173 18797 35176
rect 18831 35173 18843 35207
rect 18785 35167 18843 35173
rect 19058 35164 19064 35216
rect 19116 35204 19122 35216
rect 21284 35204 21312 35244
rect 24581 35241 24593 35244
rect 24627 35241 24639 35275
rect 25682 35272 25688 35284
rect 25643 35244 25688 35272
rect 24581 35235 24639 35241
rect 25682 35232 25688 35244
rect 25740 35232 25746 35284
rect 26234 35272 26240 35284
rect 26195 35244 26240 35272
rect 26234 35232 26240 35244
rect 26292 35272 26298 35284
rect 26789 35275 26847 35281
rect 26789 35272 26801 35275
rect 26292 35244 26801 35272
rect 26292 35232 26298 35244
rect 26789 35241 26801 35244
rect 26835 35272 26847 35275
rect 27341 35275 27399 35281
rect 27341 35272 27353 35275
rect 26835 35244 27353 35272
rect 26835 35241 26847 35244
rect 26789 35235 26847 35241
rect 27341 35241 27353 35244
rect 27387 35272 27399 35275
rect 27893 35275 27951 35281
rect 27893 35272 27905 35275
rect 27387 35244 27905 35272
rect 27387 35241 27399 35244
rect 27341 35235 27399 35241
rect 27893 35241 27905 35244
rect 27939 35241 27951 35275
rect 27893 35235 27951 35241
rect 19116 35176 21312 35204
rect 19116 35164 19122 35176
rect 21358 35164 21364 35216
rect 21416 35204 21422 35216
rect 22830 35204 22836 35216
rect 21416 35176 22836 35204
rect 21416 35164 21422 35176
rect 22830 35164 22836 35176
rect 22888 35164 22894 35216
rect 22925 35207 22983 35213
rect 22925 35173 22937 35207
rect 22971 35204 22983 35207
rect 25774 35204 25780 35216
rect 22971 35176 25780 35204
rect 22971 35173 22983 35176
rect 22925 35167 22983 35173
rect 10689 35139 10747 35145
rect 10689 35136 10701 35139
rect 4724 35108 8524 35136
rect 8588 35108 10701 35136
rect 4617 35099 4675 35105
rect 8588 35080 8616 35108
rect 10689 35105 10701 35108
rect 10735 35136 10747 35139
rect 11054 35136 11060 35148
rect 10735 35108 11060 35136
rect 10735 35105 10747 35108
rect 10689 35099 10747 35105
rect 11054 35096 11060 35108
rect 11112 35096 11118 35148
rect 15654 35136 15660 35148
rect 12084 35108 15660 35136
rect 2038 35028 2044 35080
rect 2096 35028 2102 35080
rect 3694 35028 3700 35080
rect 3752 35068 3758 35080
rect 3970 35068 3976 35080
rect 3752 35040 3976 35068
rect 3752 35028 3758 35040
rect 3970 35028 3976 35040
rect 4028 35028 4034 35080
rect 8570 35028 8576 35080
rect 8628 35068 8634 35080
rect 9122 35068 9128 35080
rect 8628 35040 8673 35068
rect 9083 35040 9128 35068
rect 8628 35028 8634 35040
rect 9122 35028 9128 35040
rect 9180 35028 9186 35080
rect 9401 35071 9459 35077
rect 9401 35037 9413 35071
rect 9447 35037 9459 35071
rect 12084 35054 12112 35108
rect 15654 35096 15660 35108
rect 15712 35096 15718 35148
rect 19426 35136 19432 35148
rect 15764 35108 19432 35136
rect 13262 35068 13268 35080
rect 13223 35040 13268 35068
rect 9401 35031 9459 35037
rect 3145 35003 3203 35009
rect 3145 34969 3157 35003
rect 3191 35000 3203 35003
rect 4893 35003 4951 35009
rect 3191 34972 4016 35000
rect 3191 34969 3203 34972
rect 3145 34963 3203 34969
rect 3988 34944 4016 34972
rect 4893 34969 4905 35003
rect 4939 35000 4951 35003
rect 5166 35000 5172 35012
rect 4939 34972 5172 35000
rect 4939 34969 4951 34972
rect 4893 34963 4951 34969
rect 5166 34960 5172 34972
rect 5224 34960 5230 35012
rect 6118 34972 7052 35000
rect 1673 34935 1731 34941
rect 1673 34901 1685 34935
rect 1719 34932 1731 34935
rect 2406 34932 2412 34944
rect 1719 34904 2412 34932
rect 1719 34901 1731 34904
rect 1673 34895 1731 34901
rect 2406 34892 2412 34904
rect 2464 34892 2470 34944
rect 3970 34892 3976 34944
rect 4028 34892 4034 34944
rect 4065 34935 4123 34941
rect 4065 34901 4077 34935
rect 4111 34932 4123 34935
rect 5626 34932 5632 34944
rect 4111 34904 5632 34932
rect 4111 34901 4123 34904
rect 4065 34895 4123 34901
rect 5626 34892 5632 34904
rect 5684 34892 5690 34944
rect 6365 34935 6423 34941
rect 6365 34901 6377 34935
rect 6411 34932 6423 34935
rect 6546 34932 6552 34944
rect 6411 34904 6552 34932
rect 6411 34901 6423 34904
rect 6365 34895 6423 34901
rect 6546 34892 6552 34904
rect 6604 34892 6610 34944
rect 7024 34932 7052 34972
rect 7834 34960 7840 35012
rect 7892 34960 7898 35012
rect 8297 35003 8355 35009
rect 8297 34969 8309 35003
rect 8343 34969 8355 35003
rect 8297 34963 8355 34969
rect 8202 34932 8208 34944
rect 7024 34904 8208 34932
rect 8202 34892 8208 34904
rect 8260 34892 8266 34944
rect 8312 34932 8340 34963
rect 8662 34960 8668 35012
rect 8720 35000 8726 35012
rect 9416 35000 9444 35031
rect 13262 35028 13268 35040
rect 13320 35028 13326 35080
rect 13814 35028 13820 35080
rect 13872 35068 13878 35080
rect 15010 35068 15016 35080
rect 13872 35040 15016 35068
rect 13872 35028 13878 35040
rect 15010 35028 15016 35040
rect 15068 35028 15074 35080
rect 15378 35028 15384 35080
rect 15436 35068 15442 35080
rect 15473 35071 15531 35077
rect 15473 35068 15485 35071
rect 15436 35040 15485 35068
rect 15436 35028 15442 35040
rect 15473 35037 15485 35040
rect 15519 35037 15531 35071
rect 15473 35031 15531 35037
rect 8720 34972 9444 35000
rect 8720 34960 8726 34972
rect 9490 34960 9496 35012
rect 9548 35000 9554 35012
rect 10965 35003 11023 35009
rect 10965 35000 10977 35003
rect 9548 34972 10977 35000
rect 9548 34960 9554 34972
rect 10965 34969 10977 34972
rect 11011 34969 11023 35003
rect 10965 34963 11023 34969
rect 12250 34960 12256 35012
rect 12308 35000 12314 35012
rect 12308 34972 12756 35000
rect 12308 34960 12314 34972
rect 8478 34932 8484 34944
rect 8312 34904 8484 34932
rect 8478 34892 8484 34904
rect 8536 34892 8542 34944
rect 8754 34892 8760 34944
rect 8812 34932 8818 34944
rect 12342 34932 12348 34944
rect 8812 34904 12348 34932
rect 8812 34892 8818 34904
rect 12342 34892 12348 34904
rect 12400 34892 12406 34944
rect 12437 34935 12495 34941
rect 12437 34901 12449 34935
rect 12483 34932 12495 34935
rect 12526 34932 12532 34944
rect 12483 34904 12532 34932
rect 12483 34901 12495 34904
rect 12437 34895 12495 34901
rect 12526 34892 12532 34904
rect 12584 34892 12590 34944
rect 12728 34932 12756 34972
rect 13722 34960 13728 35012
rect 13780 35000 13786 35012
rect 15764 35000 15792 35108
rect 19426 35096 19432 35108
rect 19484 35096 19490 35148
rect 20070 35096 20076 35148
rect 20128 35136 20134 35148
rect 20993 35139 21051 35145
rect 20128 35108 20173 35136
rect 20128 35096 20134 35108
rect 20993 35105 21005 35139
rect 21039 35105 21051 35139
rect 22940 35136 22968 35167
rect 25774 35164 25780 35176
rect 25832 35164 25838 35216
rect 25130 35136 25136 35148
rect 20993 35099 21051 35105
rect 22756 35108 22968 35136
rect 25091 35108 25136 35136
rect 16301 35071 16359 35077
rect 16301 35037 16313 35071
rect 16347 35068 16359 35071
rect 16390 35068 16396 35080
rect 16347 35040 16396 35068
rect 16347 35037 16359 35040
rect 16301 35031 16359 35037
rect 16390 35028 16396 35040
rect 16448 35028 16454 35080
rect 16850 35028 16856 35080
rect 16908 35068 16914 35080
rect 17221 35071 17279 35077
rect 17221 35068 17233 35071
rect 16908 35040 17233 35068
rect 16908 35028 16914 35040
rect 17221 35037 17233 35040
rect 17267 35037 17279 35071
rect 17221 35031 17279 35037
rect 17310 35028 17316 35080
rect 17368 35068 17374 35080
rect 17865 35071 17923 35077
rect 17368 35040 17413 35068
rect 17368 35028 17374 35040
rect 17865 35037 17877 35071
rect 17911 35037 17923 35071
rect 17865 35031 17923 35037
rect 17957 35071 18015 35077
rect 17957 35037 17969 35071
rect 18003 35070 18015 35071
rect 18003 35068 18092 35070
rect 18690 35068 18696 35080
rect 18003 35042 18696 35068
rect 18003 35037 18015 35042
rect 18064 35040 18696 35042
rect 17957 35031 18015 35037
rect 13780 34972 15792 35000
rect 13780 34960 13786 34972
rect 15838 34960 15844 35012
rect 15896 35000 15902 35012
rect 16209 35003 16267 35009
rect 16209 35000 16221 35003
rect 15896 34972 16221 35000
rect 15896 34960 15902 34972
rect 16209 34969 16221 34972
rect 16255 34969 16267 35003
rect 16209 34963 16267 34969
rect 16482 34960 16488 35012
rect 16540 35000 16546 35012
rect 17880 35000 17908 35031
rect 18690 35028 18696 35040
rect 18748 35028 18754 35080
rect 18877 35071 18935 35077
rect 18877 35037 18889 35071
rect 18923 35068 18935 35071
rect 19889 35071 19947 35077
rect 18923 35040 19334 35068
rect 18923 35037 18935 35040
rect 18877 35031 18935 35037
rect 16540 34972 17908 35000
rect 16540 34960 16546 34972
rect 18046 34960 18052 35012
rect 18104 35000 18110 35012
rect 19058 35000 19064 35012
rect 18104 34972 19064 35000
rect 18104 34960 18110 34972
rect 19058 34960 19064 34972
rect 19116 34960 19122 35012
rect 19306 35000 19334 35040
rect 19889 35037 19901 35071
rect 19935 35037 19947 35071
rect 19889 35031 19947 35037
rect 20809 35071 20867 35077
rect 20809 35037 20821 35071
rect 20855 35037 20867 35071
rect 20809 35031 20867 35037
rect 19904 35000 19932 35031
rect 19978 35000 19984 35012
rect 19306 34972 19984 35000
rect 19978 34960 19984 34972
rect 20036 35000 20042 35012
rect 20824 35000 20852 35031
rect 21008 35012 21036 35099
rect 21082 35028 21088 35080
rect 21140 35068 21146 35080
rect 22756 35068 22784 35108
rect 25130 35096 25136 35108
rect 25188 35096 25194 35148
rect 21140 35040 22784 35068
rect 21140 35028 21146 35040
rect 20036 34972 20852 35000
rect 20036 34960 20042 34972
rect 20990 34960 20996 35012
rect 21048 35000 21054 35012
rect 23198 35000 23204 35012
rect 21048 34972 23204 35000
rect 21048 34960 21054 34972
rect 23198 34960 23204 34972
rect 23256 34960 23262 35012
rect 13081 34935 13139 34941
rect 13081 34932 13093 34935
rect 12728 34904 13093 34932
rect 13081 34901 13093 34904
rect 13127 34901 13139 34935
rect 14274 34932 14280 34944
rect 14235 34904 14280 34932
rect 13081 34895 13139 34901
rect 14274 34892 14280 34904
rect 14332 34892 14338 34944
rect 14921 34935 14979 34941
rect 14921 34901 14933 34935
rect 14967 34932 14979 34935
rect 15010 34932 15016 34944
rect 14967 34904 15016 34932
rect 14967 34901 14979 34904
rect 14921 34895 14979 34901
rect 15010 34892 15016 34904
rect 15068 34892 15074 34944
rect 15565 34935 15623 34941
rect 15565 34901 15577 34935
rect 15611 34932 15623 34935
rect 16022 34932 16028 34944
rect 15611 34904 16028 34932
rect 15611 34901 15623 34904
rect 15565 34895 15623 34901
rect 16022 34892 16028 34904
rect 16080 34892 16086 34944
rect 16390 34892 16396 34944
rect 16448 34932 16454 34944
rect 21729 34935 21787 34941
rect 21729 34932 21741 34935
rect 16448 34904 21741 34932
rect 16448 34892 16454 34904
rect 21729 34901 21741 34904
rect 21775 34901 21787 34935
rect 22370 34932 22376 34944
rect 22331 34904 22376 34932
rect 21729 34895 21787 34901
rect 22370 34892 22376 34904
rect 22428 34892 22434 34944
rect 23477 34935 23535 34941
rect 23477 34901 23489 34935
rect 23523 34932 23535 34935
rect 24026 34932 24032 34944
rect 23523 34904 24032 34932
rect 23523 34901 23535 34904
rect 23477 34895 23535 34901
rect 24026 34892 24032 34904
rect 24084 34892 24090 34944
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 3786 34728 3792 34740
rect 2608 34700 3792 34728
rect 2608 34601 2636 34700
rect 3786 34688 3792 34700
rect 3844 34688 3850 34740
rect 3878 34688 3884 34740
rect 3936 34728 3942 34740
rect 8202 34728 8208 34740
rect 3936 34700 5488 34728
rect 3936 34688 3942 34700
rect 3142 34620 3148 34672
rect 3200 34660 3206 34672
rect 3694 34660 3700 34672
rect 3200 34632 3700 34660
rect 3200 34620 3206 34632
rect 3694 34620 3700 34632
rect 3752 34620 3758 34672
rect 4614 34620 4620 34672
rect 4672 34620 4678 34672
rect 5460 34660 5488 34700
rect 7668 34700 8208 34728
rect 7190 34660 7196 34672
rect 5460 34632 5580 34660
rect 5552 34604 5580 34632
rect 5736 34632 7196 34660
rect 2593 34595 2651 34601
rect 2593 34561 2605 34595
rect 2639 34561 2651 34595
rect 2593 34555 2651 34561
rect 5534 34552 5540 34604
rect 5592 34592 5598 34604
rect 5592 34564 5685 34592
rect 5592 34552 5598 34564
rect 1946 34484 1952 34536
rect 2004 34524 2010 34536
rect 2869 34527 2927 34533
rect 2869 34524 2881 34527
rect 2004 34496 2881 34524
rect 2004 34484 2010 34496
rect 2869 34493 2881 34496
rect 2915 34524 2927 34527
rect 3694 34524 3700 34536
rect 2915 34496 3700 34524
rect 2915 34493 2927 34496
rect 2869 34487 2927 34493
rect 3694 34484 3700 34496
rect 3752 34484 3758 34536
rect 3789 34527 3847 34533
rect 3789 34493 3801 34527
rect 3835 34524 3847 34527
rect 5736 34524 5764 34632
rect 7190 34620 7196 34632
rect 7248 34620 7254 34672
rect 5810 34552 5816 34604
rect 5868 34592 5874 34604
rect 6549 34595 6607 34601
rect 6549 34592 6561 34595
rect 5868 34564 6561 34592
rect 5868 34552 5874 34564
rect 6549 34561 6561 34564
rect 6595 34592 6607 34595
rect 7668 34592 7696 34700
rect 8202 34688 8208 34700
rect 8260 34688 8266 34740
rect 8846 34688 8852 34740
rect 8904 34728 8910 34740
rect 10413 34731 10471 34737
rect 10413 34728 10425 34731
rect 8904 34700 10425 34728
rect 8904 34688 8910 34700
rect 10413 34697 10425 34700
rect 10459 34697 10471 34731
rect 10413 34691 10471 34697
rect 10686 34688 10692 34740
rect 10744 34728 10750 34740
rect 11057 34731 11115 34737
rect 11057 34728 11069 34731
rect 10744 34700 11069 34728
rect 10744 34688 10750 34700
rect 11057 34697 11069 34700
rect 11103 34697 11115 34731
rect 11057 34691 11115 34697
rect 12158 34688 12164 34740
rect 12216 34728 12222 34740
rect 14274 34728 14280 34740
rect 12216 34700 14280 34728
rect 12216 34688 12222 34700
rect 8510 34632 9352 34660
rect 6595 34564 7696 34592
rect 6595 34561 6607 34564
rect 6549 34555 6607 34561
rect 3835 34496 5764 34524
rect 6641 34527 6699 34533
rect 3835 34493 3847 34496
rect 3789 34487 3847 34493
rect 6641 34493 6653 34527
rect 6687 34524 6699 34527
rect 6914 34524 6920 34536
rect 6687 34496 6920 34524
rect 6687 34493 6699 34496
rect 6641 34487 6699 34493
rect 6914 34484 6920 34496
rect 6972 34484 6978 34536
rect 7193 34527 7251 34533
rect 7193 34493 7205 34527
rect 7239 34524 7251 34527
rect 7282 34524 7288 34536
rect 7239 34496 7288 34524
rect 7239 34493 7251 34496
rect 7193 34487 7251 34493
rect 7282 34484 7288 34496
rect 7340 34524 7346 34536
rect 8202 34524 8208 34536
rect 7340 34496 8208 34524
rect 7340 34484 7346 34496
rect 8202 34484 8208 34496
rect 8260 34484 8266 34536
rect 8938 34524 8944 34536
rect 8899 34496 8944 34524
rect 8938 34484 8944 34496
rect 8996 34484 9002 34536
rect 9217 34527 9275 34533
rect 9217 34493 9229 34527
rect 9263 34493 9275 34527
rect 9217 34487 9275 34493
rect 7926 34456 7932 34468
rect 5460 34428 7932 34456
rect 5460 34400 5488 34428
rect 7926 34416 7932 34428
rect 7984 34416 7990 34468
rect 5258 34348 5264 34400
rect 5316 34397 5322 34400
rect 5316 34391 5331 34397
rect 5319 34357 5331 34391
rect 5316 34351 5331 34357
rect 5316 34348 5322 34351
rect 5442 34348 5448 34400
rect 5500 34348 5506 34400
rect 7006 34348 7012 34400
rect 7064 34388 7070 34400
rect 7558 34388 7564 34400
rect 7064 34360 7564 34388
rect 7064 34348 7070 34360
rect 7558 34348 7564 34360
rect 7616 34348 7622 34400
rect 7834 34348 7840 34400
rect 7892 34388 7898 34400
rect 8570 34388 8576 34400
rect 7892 34360 8576 34388
rect 7892 34348 7898 34360
rect 8570 34348 8576 34360
rect 8628 34388 8634 34400
rect 9232 34388 9260 34487
rect 9324 34456 9352 34632
rect 9674 34620 9680 34672
rect 9732 34660 9738 34672
rect 9769 34663 9827 34669
rect 9769 34660 9781 34663
rect 9732 34632 9781 34660
rect 9732 34620 9738 34632
rect 9769 34629 9781 34632
rect 9815 34629 9827 34663
rect 13262 34660 13268 34672
rect 12742 34632 13268 34660
rect 9769 34623 9827 34629
rect 13262 34620 13268 34632
rect 13320 34620 13326 34672
rect 9858 34552 9864 34604
rect 9916 34592 9922 34604
rect 10502 34592 10508 34604
rect 9916 34564 9961 34592
rect 10415 34564 10508 34592
rect 9916 34552 9922 34564
rect 10502 34552 10508 34564
rect 10560 34592 10566 34604
rect 11146 34592 11152 34604
rect 10560 34564 11152 34592
rect 10560 34552 10566 34564
rect 11146 34552 11152 34564
rect 11204 34552 11210 34604
rect 13464 34601 13492 34700
rect 14274 34688 14280 34700
rect 14332 34688 14338 34740
rect 14366 34688 14372 34740
rect 14424 34728 14430 34740
rect 15102 34728 15108 34740
rect 14424 34700 15108 34728
rect 14424 34688 14430 34700
rect 15102 34688 15108 34700
rect 15160 34688 15166 34740
rect 15654 34688 15660 34740
rect 15712 34728 15718 34740
rect 18233 34731 18291 34737
rect 18233 34728 18245 34731
rect 15712 34700 18245 34728
rect 15712 34688 15718 34700
rect 18233 34697 18245 34700
rect 18279 34697 18291 34731
rect 18233 34691 18291 34697
rect 19242 34688 19248 34740
rect 19300 34728 19306 34740
rect 21358 34728 21364 34740
rect 19300 34700 21364 34728
rect 19300 34688 19306 34700
rect 21358 34688 21364 34700
rect 21416 34688 21422 34740
rect 22738 34688 22744 34740
rect 22796 34728 22802 34740
rect 25317 34731 25375 34737
rect 25317 34728 25329 34731
rect 22796 34700 25329 34728
rect 22796 34688 22802 34700
rect 25317 34697 25329 34700
rect 25363 34697 25375 34731
rect 25317 34691 25375 34697
rect 26513 34731 26571 34737
rect 26513 34697 26525 34731
rect 26559 34728 26571 34731
rect 28994 34728 29000 34740
rect 26559 34700 29000 34728
rect 26559 34697 26571 34700
rect 26513 34691 26571 34697
rect 14090 34620 14096 34672
rect 14148 34660 14154 34672
rect 17402 34660 17408 34672
rect 14148 34632 16252 34660
rect 17363 34632 17408 34660
rect 14148 34620 14154 34632
rect 13449 34595 13507 34601
rect 13449 34561 13461 34595
rect 13495 34561 13507 34595
rect 13449 34555 13507 34561
rect 13538 34552 13544 34604
rect 13596 34592 13602 34604
rect 13909 34595 13967 34601
rect 13909 34592 13921 34595
rect 13596 34564 13921 34592
rect 13596 34552 13602 34564
rect 13909 34561 13921 34564
rect 13955 34592 13967 34595
rect 14642 34592 14648 34604
rect 13955 34564 14648 34592
rect 13955 34561 13967 34564
rect 13909 34555 13967 34561
rect 14642 34552 14648 34564
rect 14700 34552 14706 34604
rect 14826 34592 14832 34604
rect 14787 34564 14832 34592
rect 14826 34552 14832 34564
rect 14884 34552 14890 34604
rect 15286 34552 15292 34604
rect 15344 34592 15350 34604
rect 15565 34595 15623 34601
rect 15565 34592 15577 34595
rect 15344 34564 15577 34592
rect 15344 34552 15350 34564
rect 15565 34561 15577 34564
rect 15611 34561 15623 34595
rect 15565 34555 15623 34561
rect 9398 34484 9404 34536
rect 9456 34524 9462 34536
rect 13078 34524 13084 34536
rect 9456 34496 13084 34524
rect 9456 34484 9462 34496
rect 13078 34484 13084 34496
rect 13136 34484 13142 34536
rect 13173 34527 13231 34533
rect 13173 34493 13185 34527
rect 13219 34524 13231 34527
rect 13630 34524 13636 34536
rect 13219 34496 13636 34524
rect 13219 34493 13231 34496
rect 13173 34487 13231 34493
rect 13630 34484 13636 34496
rect 13688 34484 13694 34536
rect 14550 34484 14556 34536
rect 14608 34524 14614 34536
rect 14737 34527 14795 34533
rect 14737 34524 14749 34527
rect 14608 34496 14749 34524
rect 14608 34484 14614 34496
rect 14737 34493 14749 34496
rect 14783 34493 14795 34527
rect 14737 34487 14795 34493
rect 15473 34527 15531 34533
rect 15473 34493 15485 34527
rect 15519 34524 15531 34527
rect 15654 34524 15660 34536
rect 15519 34496 15660 34524
rect 15519 34493 15531 34496
rect 15473 34487 15531 34493
rect 15654 34484 15660 34496
rect 15712 34484 15718 34536
rect 15746 34484 15752 34536
rect 15804 34524 15810 34536
rect 16025 34527 16083 34533
rect 16025 34524 16037 34527
rect 15804 34496 16037 34524
rect 15804 34484 15810 34496
rect 16025 34493 16037 34496
rect 16071 34493 16083 34527
rect 16224 34524 16252 34632
rect 17402 34620 17408 34632
rect 17460 34620 17466 34672
rect 17497 34663 17555 34669
rect 17497 34629 17509 34663
rect 17543 34660 17555 34663
rect 17678 34660 17684 34672
rect 17543 34632 17684 34660
rect 17543 34629 17555 34632
rect 17497 34623 17555 34629
rect 17678 34620 17684 34632
rect 17736 34620 17742 34672
rect 17862 34620 17868 34672
rect 17920 34660 17926 34672
rect 17920 34632 20116 34660
rect 17920 34620 17926 34632
rect 16850 34592 16856 34604
rect 16811 34564 16856 34592
rect 16850 34552 16856 34564
rect 16908 34552 16914 34604
rect 18325 34595 18383 34601
rect 18325 34561 18337 34595
rect 18371 34592 18383 34595
rect 18966 34592 18972 34604
rect 18371 34564 18972 34592
rect 18371 34561 18383 34564
rect 18325 34555 18383 34561
rect 18966 34552 18972 34564
rect 19024 34552 19030 34604
rect 19889 34595 19947 34601
rect 19889 34561 19901 34595
rect 19935 34592 19947 34595
rect 19978 34592 19984 34604
rect 19935 34564 19984 34592
rect 19935 34561 19947 34564
rect 19889 34555 19947 34561
rect 19978 34552 19984 34564
rect 20036 34552 20042 34604
rect 20088 34592 20116 34632
rect 21818 34620 21824 34672
rect 21876 34660 21882 34672
rect 22557 34663 22615 34669
rect 22557 34660 22569 34663
rect 21876 34632 22569 34660
rect 21876 34620 21882 34632
rect 22557 34629 22569 34632
rect 22603 34629 22615 34663
rect 23198 34660 23204 34672
rect 23111 34632 23204 34660
rect 22557 34623 22615 34629
rect 23198 34620 23204 34632
rect 23256 34660 23262 34672
rect 26528 34660 26556 34691
rect 28994 34688 29000 34700
rect 29052 34688 29058 34740
rect 37734 34660 37740 34672
rect 23256 34632 26556 34660
rect 35866 34632 37740 34660
rect 23256 34620 23262 34632
rect 22005 34595 22063 34601
rect 22005 34592 22017 34595
rect 20088 34564 22017 34592
rect 22005 34561 22017 34564
rect 22051 34561 22063 34595
rect 22005 34555 22063 34561
rect 18877 34527 18935 34533
rect 18877 34524 18889 34527
rect 16224 34496 18889 34524
rect 16025 34487 16083 34493
rect 18877 34493 18889 34496
rect 18923 34493 18935 34527
rect 18877 34487 18935 34493
rect 20165 34527 20223 34533
rect 20165 34493 20177 34527
rect 20211 34524 20223 34527
rect 24302 34524 24308 34536
rect 20211 34496 20852 34524
rect 24215 34496 24308 34524
rect 20211 34493 20223 34496
rect 20165 34487 20223 34493
rect 19426 34456 19432 34468
rect 9324 34428 12112 34456
rect 9306 34388 9312 34400
rect 8628 34360 9312 34388
rect 8628 34348 8634 34360
rect 9306 34348 9312 34360
rect 9364 34348 9370 34400
rect 9674 34348 9680 34400
rect 9732 34388 9738 34400
rect 11606 34388 11612 34400
rect 9732 34360 11612 34388
rect 9732 34348 9738 34360
rect 11606 34348 11612 34360
rect 11664 34348 11670 34400
rect 11701 34391 11759 34397
rect 11701 34357 11713 34391
rect 11747 34388 11759 34391
rect 11974 34388 11980 34400
rect 11747 34360 11980 34388
rect 11747 34357 11759 34360
rect 11701 34351 11759 34357
rect 11974 34348 11980 34360
rect 12032 34348 12038 34400
rect 12084 34388 12112 34428
rect 14016 34428 19432 34456
rect 14016 34388 14044 34428
rect 19426 34416 19432 34428
rect 19484 34416 19490 34468
rect 20824 34400 20852 34496
rect 24302 34484 24308 34496
rect 24360 34524 24366 34536
rect 35866 34524 35894 34632
rect 37734 34620 37740 34632
rect 37792 34620 37798 34672
rect 24360 34496 35894 34524
rect 24360 34484 24366 34496
rect 24026 34416 24032 34468
rect 24084 34456 24090 34468
rect 24765 34459 24823 34465
rect 24765 34456 24777 34459
rect 24084 34428 24777 34456
rect 24084 34416 24090 34428
rect 24765 34425 24777 34428
rect 24811 34456 24823 34459
rect 25682 34456 25688 34468
rect 24811 34428 25688 34456
rect 24811 34425 24823 34428
rect 24765 34419 24823 34425
rect 25682 34416 25688 34428
rect 25740 34456 25746 34468
rect 25869 34459 25927 34465
rect 25869 34456 25881 34459
rect 25740 34428 25881 34456
rect 25740 34416 25746 34428
rect 25869 34425 25881 34428
rect 25915 34456 25927 34459
rect 27157 34459 27215 34465
rect 27157 34456 27169 34459
rect 25915 34428 27169 34456
rect 25915 34425 25927 34428
rect 25869 34419 25927 34425
rect 27157 34425 27169 34428
rect 27203 34425 27215 34459
rect 27157 34419 27215 34425
rect 12084 34360 14044 34388
rect 14093 34391 14151 34397
rect 14093 34357 14105 34391
rect 14139 34388 14151 34391
rect 15194 34388 15200 34400
rect 14139 34360 15200 34388
rect 14139 34357 14151 34360
rect 14093 34351 14151 34357
rect 15194 34348 15200 34360
rect 15252 34348 15258 34400
rect 15378 34348 15384 34400
rect 15436 34388 15442 34400
rect 20714 34388 20720 34400
rect 15436 34360 20720 34388
rect 15436 34348 15442 34360
rect 20714 34348 20720 34360
rect 20772 34348 20778 34400
rect 20806 34348 20812 34400
rect 20864 34388 20870 34400
rect 23658 34388 23664 34400
rect 20864 34360 20909 34388
rect 23619 34360 23664 34388
rect 20864 34348 20870 34360
rect 23658 34348 23664 34360
rect 23716 34348 23722 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 1936 34187 1994 34193
rect 1936 34153 1948 34187
rect 1982 34184 1994 34187
rect 2498 34184 2504 34196
rect 1982 34156 2504 34184
rect 1982 34153 1994 34156
rect 1936 34147 1994 34153
rect 2498 34144 2504 34156
rect 2556 34184 2562 34196
rect 4801 34187 4859 34193
rect 2556 34156 3832 34184
rect 2556 34144 2562 34156
rect 1673 34051 1731 34057
rect 1673 34017 1685 34051
rect 1719 34048 1731 34051
rect 2958 34048 2964 34060
rect 1719 34020 2964 34048
rect 1719 34017 1731 34020
rect 1673 34011 1731 34017
rect 2958 34008 2964 34020
rect 3016 34048 3022 34060
rect 3418 34048 3424 34060
rect 3016 34020 3424 34048
rect 3016 34008 3022 34020
rect 3418 34008 3424 34020
rect 3476 34008 3482 34060
rect 2056 33884 2438 33912
rect 1118 33804 1124 33856
rect 1176 33844 1182 33856
rect 2056 33844 2084 33884
rect 3418 33844 3424 33856
rect 1176 33816 2084 33844
rect 3379 33816 3424 33844
rect 1176 33804 1182 33816
rect 3418 33804 3424 33816
rect 3476 33804 3482 33856
rect 3804 33844 3832 34156
rect 4801 34153 4813 34187
rect 4847 34184 4859 34187
rect 5074 34184 5080 34196
rect 4847 34156 5080 34184
rect 4847 34153 4859 34156
rect 4801 34147 4859 34153
rect 5074 34144 5080 34156
rect 5132 34144 5138 34196
rect 5258 34144 5264 34196
rect 5316 34184 5322 34196
rect 7650 34184 7656 34196
rect 5316 34156 7656 34184
rect 5316 34144 5322 34156
rect 5368 34057 5396 34156
rect 7650 34144 7656 34156
rect 7708 34144 7714 34196
rect 7834 34184 7840 34196
rect 7760 34156 7840 34184
rect 7760 34116 7788 34156
rect 7834 34144 7840 34156
rect 7892 34144 7898 34196
rect 8294 34144 8300 34196
rect 8352 34184 8358 34196
rect 9217 34187 9275 34193
rect 9217 34184 9229 34187
rect 8352 34156 9229 34184
rect 8352 34144 8358 34156
rect 9217 34153 9229 34156
rect 9263 34153 9275 34187
rect 9766 34184 9772 34196
rect 9727 34156 9772 34184
rect 9217 34147 9275 34153
rect 9766 34144 9772 34156
rect 9824 34144 9830 34196
rect 10704 34156 12112 34184
rect 7392 34088 7788 34116
rect 5353 34051 5411 34057
rect 3988 34020 4936 34048
rect 3988 33989 4016 34020
rect 3973 33983 4031 33989
rect 3973 33949 3985 33983
rect 4019 33949 4031 33983
rect 3973 33943 4031 33949
rect 4617 33983 4675 33989
rect 4617 33949 4629 33983
rect 4663 33980 4675 33983
rect 4798 33980 4804 33992
rect 4663 33952 4804 33980
rect 4663 33949 4675 33952
rect 4617 33943 4675 33949
rect 4798 33940 4804 33952
rect 4856 33940 4862 33992
rect 4908 33980 4936 34020
rect 5353 34017 5365 34051
rect 5399 34017 5411 34051
rect 5353 34011 5411 34017
rect 5534 34008 5540 34060
rect 5592 34048 5598 34060
rect 7392 34057 7420 34088
rect 9582 34076 9588 34128
rect 9640 34116 9646 34128
rect 10704 34116 10732 34156
rect 9640 34088 10732 34116
rect 9640 34076 9646 34088
rect 10778 34076 10784 34128
rect 10836 34076 10842 34128
rect 12084 34116 12112 34156
rect 12342 34144 12348 34196
rect 12400 34184 12406 34196
rect 14274 34184 14280 34196
rect 12400 34156 14280 34184
rect 12400 34144 12406 34156
rect 14274 34144 14280 34156
rect 14332 34144 14338 34196
rect 14366 34144 14372 34196
rect 14424 34184 14430 34196
rect 21726 34184 21732 34196
rect 14424 34156 21732 34184
rect 14424 34144 14430 34156
rect 21726 34144 21732 34156
rect 21784 34144 21790 34196
rect 22830 34184 22836 34196
rect 21836 34156 22836 34184
rect 12084 34088 12388 34116
rect 7377 34051 7435 34057
rect 7377 34048 7389 34051
rect 5592 34020 7389 34048
rect 5592 34008 5598 34020
rect 7377 34017 7389 34020
rect 7423 34017 7435 34051
rect 10796 34048 10824 34076
rect 7377 34011 7435 34017
rect 8036 34020 10824 34048
rect 4982 33980 4988 33992
rect 4908 33952 4988 33980
rect 4982 33940 4988 33952
rect 5040 33980 5046 33992
rect 5442 33980 5448 33992
rect 5040 33952 5448 33980
rect 5040 33940 5046 33952
rect 5442 33940 5448 33952
rect 5500 33940 5506 33992
rect 5626 33940 5632 33992
rect 5684 33980 5690 33992
rect 5684 33952 6026 33980
rect 5684 33940 5690 33952
rect 7466 33940 7472 33992
rect 7524 33980 7530 33992
rect 7742 33980 7748 33992
rect 7524 33952 7748 33980
rect 7524 33940 7530 33952
rect 7742 33940 7748 33952
rect 7800 33940 7806 33992
rect 7837 33983 7895 33989
rect 7837 33949 7849 33983
rect 7883 33980 7895 33983
rect 7926 33980 7932 33992
rect 7883 33952 7932 33980
rect 7883 33949 7895 33952
rect 7837 33943 7895 33949
rect 7926 33940 7932 33952
rect 7984 33980 7990 33992
rect 8036 33980 8064 34020
rect 11146 34008 11152 34060
rect 11204 34048 11210 34060
rect 12158 34048 12164 34060
rect 11204 34020 12164 34048
rect 11204 34008 11210 34020
rect 12158 34008 12164 34020
rect 12216 34008 12222 34060
rect 12360 34048 12388 34088
rect 12434 34076 12440 34128
rect 12492 34116 12498 34128
rect 20530 34116 20536 34128
rect 12492 34088 20536 34116
rect 12492 34076 12498 34088
rect 12360 34020 16068 34048
rect 7984 33952 8077 33980
rect 7984 33940 7990 33952
rect 8294 33940 8300 33992
rect 8352 33980 8358 33992
rect 9309 33983 9367 33989
rect 9309 33980 9321 33983
rect 8352 33952 9321 33980
rect 8352 33940 8358 33952
rect 9309 33949 9321 33952
rect 9355 33980 9367 33983
rect 9950 33980 9956 33992
rect 9355 33952 9956 33980
rect 9355 33949 9367 33952
rect 9309 33943 9367 33949
rect 9950 33940 9956 33952
rect 10008 33980 10014 33992
rect 10594 33980 10600 33992
rect 10008 33952 10600 33980
rect 10008 33940 10014 33952
rect 10594 33940 10600 33952
rect 10652 33940 10658 33992
rect 13081 33983 13139 33989
rect 13081 33980 13093 33983
rect 12176 33952 13093 33980
rect 3988 33884 5764 33912
rect 3988 33844 4016 33884
rect 3804 33816 4016 33844
rect 4065 33847 4123 33853
rect 4065 33813 4077 33847
rect 4111 33844 4123 33847
rect 5626 33844 5632 33856
rect 4111 33816 5632 33844
rect 4111 33813 4123 33816
rect 4065 33807 4123 33813
rect 5626 33804 5632 33816
rect 5684 33804 5690 33856
rect 5736 33844 5764 33884
rect 7006 33872 7012 33924
rect 7064 33912 7070 33924
rect 7101 33915 7159 33921
rect 7101 33912 7113 33915
rect 7064 33884 7113 33912
rect 7064 33872 7070 33884
rect 7101 33881 7113 33884
rect 7147 33881 7159 33915
rect 8754 33912 8760 33924
rect 7101 33875 7159 33881
rect 7208 33884 8760 33912
rect 7208 33844 7236 33884
rect 8754 33872 8760 33884
rect 8812 33872 8818 33924
rect 11422 33872 11428 33924
rect 11480 33872 11486 33924
rect 11790 33872 11796 33924
rect 11848 33912 11854 33924
rect 11885 33915 11943 33921
rect 11885 33912 11897 33915
rect 11848 33884 11897 33912
rect 11848 33872 11854 33884
rect 11885 33881 11897 33884
rect 11931 33881 11943 33915
rect 11885 33875 11943 33881
rect 7926 33844 7932 33856
rect 5736 33816 7236 33844
rect 7887 33816 7932 33844
rect 7926 33804 7932 33816
rect 7984 33804 7990 33856
rect 8573 33847 8631 33853
rect 8573 33813 8585 33847
rect 8619 33844 8631 33847
rect 10413 33847 10471 33853
rect 10413 33844 10425 33847
rect 8619 33816 10425 33844
rect 8619 33813 8631 33816
rect 8573 33807 8631 33813
rect 10413 33813 10425 33816
rect 10459 33844 10471 33847
rect 11514 33844 11520 33856
rect 10459 33816 11520 33844
rect 10459 33813 10471 33816
rect 10413 33807 10471 33813
rect 11514 33804 11520 33816
rect 11572 33804 11578 33856
rect 11606 33804 11612 33856
rect 11664 33844 11670 33856
rect 12176 33844 12204 33952
rect 13081 33949 13093 33952
rect 13127 33949 13139 33983
rect 13081 33943 13139 33949
rect 13262 33940 13268 33992
rect 13320 33980 13326 33992
rect 13538 33980 13544 33992
rect 13320 33952 13544 33980
rect 13320 33940 13326 33952
rect 13538 33940 13544 33952
rect 13596 33940 13602 33992
rect 14829 33983 14887 33989
rect 14660 33980 14780 33982
rect 14829 33980 14841 33983
rect 14292 33954 14841 33980
rect 14292 33952 14688 33954
rect 14752 33952 14841 33954
rect 12434 33872 12440 33924
rect 12492 33912 12498 33924
rect 14292 33912 14320 33952
rect 14829 33949 14841 33952
rect 14875 33980 14887 33983
rect 15194 33980 15200 33992
rect 14875 33952 15200 33980
rect 14875 33949 14887 33952
rect 14829 33943 14887 33949
rect 15194 33940 15200 33952
rect 15252 33940 15258 33992
rect 16040 33980 16068 34020
rect 16482 34008 16488 34060
rect 16540 34048 16546 34060
rect 19518 34048 19524 34060
rect 16540 34020 19334 34048
rect 19479 34020 19524 34048
rect 16540 34008 16546 34020
rect 17037 33983 17095 33989
rect 17037 33980 17049 33983
rect 16040 33952 17049 33980
rect 17037 33949 17049 33952
rect 17083 33949 17095 33983
rect 17037 33943 17095 33949
rect 17218 33940 17224 33992
rect 17276 33980 17282 33992
rect 17862 33980 17868 33992
rect 17276 33952 17868 33980
rect 17276 33940 17282 33952
rect 17862 33940 17868 33952
rect 17920 33940 17926 33992
rect 12492 33884 14320 33912
rect 14737 33915 14795 33921
rect 12492 33872 12498 33884
rect 14737 33881 14749 33915
rect 14783 33912 14795 33915
rect 14918 33912 14924 33924
rect 14783 33884 14924 33912
rect 14783 33881 14795 33884
rect 14737 33875 14795 33881
rect 14918 33872 14924 33884
rect 14976 33872 14982 33924
rect 15010 33872 15016 33924
rect 15068 33912 15074 33924
rect 15381 33915 15439 33921
rect 15381 33912 15393 33915
rect 15068 33884 15393 33912
rect 15068 33872 15074 33884
rect 15381 33881 15393 33884
rect 15427 33881 15439 33915
rect 15381 33875 15439 33881
rect 15473 33915 15531 33921
rect 15473 33881 15485 33915
rect 15519 33912 15531 33915
rect 15838 33912 15844 33924
rect 15519 33884 15844 33912
rect 15519 33881 15531 33884
rect 15473 33875 15531 33881
rect 15838 33872 15844 33884
rect 15896 33872 15902 33924
rect 16025 33915 16083 33921
rect 16025 33881 16037 33915
rect 16071 33912 16083 33915
rect 16114 33912 16120 33924
rect 16071 33884 16120 33912
rect 16071 33881 16083 33884
rect 16025 33875 16083 33881
rect 16114 33872 16120 33884
rect 16172 33872 16178 33924
rect 16482 33912 16488 33924
rect 16443 33884 16488 33912
rect 16482 33872 16488 33884
rect 16540 33872 16546 33924
rect 17129 33915 17187 33921
rect 17129 33881 17141 33915
rect 17175 33912 17187 33915
rect 17175 33884 17356 33912
rect 17175 33881 17187 33884
rect 17129 33875 17187 33881
rect 11664 33816 12204 33844
rect 13173 33847 13231 33853
rect 11664 33804 11670 33816
rect 13173 33813 13185 33847
rect 13219 33844 13231 33847
rect 13722 33844 13728 33856
rect 13219 33816 13728 33844
rect 13219 33813 13231 33816
rect 13173 33807 13231 33813
rect 13722 33804 13728 33816
rect 13780 33804 13786 33856
rect 14274 33804 14280 33856
rect 14332 33844 14338 33856
rect 17218 33844 17224 33856
rect 14332 33816 17224 33844
rect 14332 33804 14338 33816
rect 17218 33804 17224 33816
rect 17276 33804 17282 33856
rect 17328 33844 17356 33884
rect 17494 33872 17500 33924
rect 17552 33912 17558 33924
rect 17954 33912 17960 33924
rect 17552 33884 17960 33912
rect 17552 33872 17558 33884
rect 17954 33872 17960 33884
rect 18012 33872 18018 33924
rect 18138 33912 18144 33924
rect 18099 33884 18144 33912
rect 18138 33872 18144 33884
rect 18196 33872 18202 33924
rect 18230 33872 18236 33924
rect 18288 33912 18294 33924
rect 18782 33912 18788 33924
rect 18288 33884 18333 33912
rect 18743 33884 18788 33912
rect 18288 33872 18294 33884
rect 18782 33872 18788 33884
rect 18840 33872 18846 33924
rect 17678 33844 17684 33856
rect 17328 33816 17684 33844
rect 17678 33804 17684 33816
rect 17736 33804 17742 33856
rect 19306 33844 19334 34020
rect 19518 34008 19524 34020
rect 19576 34008 19582 34060
rect 20180 34057 20208 34088
rect 20530 34076 20536 34088
rect 20588 34076 20594 34128
rect 20714 34076 20720 34128
rect 20772 34116 20778 34128
rect 21453 34119 21511 34125
rect 21453 34116 21465 34119
rect 20772 34088 21465 34116
rect 20772 34076 20778 34088
rect 21453 34085 21465 34088
rect 21499 34116 21511 34119
rect 21836 34116 21864 34156
rect 22830 34144 22836 34156
rect 22888 34144 22894 34196
rect 23198 34184 23204 34196
rect 23159 34156 23204 34184
rect 23198 34144 23204 34156
rect 23256 34144 23262 34196
rect 25682 34184 25688 34196
rect 25643 34156 25688 34184
rect 25682 34144 25688 34156
rect 25740 34184 25746 34196
rect 26237 34187 26295 34193
rect 26237 34184 26249 34187
rect 25740 34156 26249 34184
rect 25740 34144 25746 34156
rect 26237 34153 26249 34156
rect 26283 34153 26295 34187
rect 26237 34147 26295 34153
rect 26326 34144 26332 34196
rect 26384 34184 26390 34196
rect 37458 34184 37464 34196
rect 26384 34156 37464 34184
rect 26384 34144 26390 34156
rect 37458 34144 37464 34156
rect 37516 34144 37522 34196
rect 25406 34116 25412 34128
rect 21499 34088 21864 34116
rect 21928 34088 25412 34116
rect 21499 34085 21511 34088
rect 21453 34079 21511 34085
rect 20165 34051 20223 34057
rect 20165 34017 20177 34051
rect 20211 34017 20223 34051
rect 21928 34048 21956 34088
rect 25406 34076 25412 34088
rect 25464 34076 25470 34128
rect 38010 34116 38016 34128
rect 35866 34088 38016 34116
rect 20165 34011 20223 34017
rect 20456 34020 21956 34048
rect 19978 33980 19984 33992
rect 19939 33952 19984 33980
rect 19978 33940 19984 33952
rect 20036 33940 20042 33992
rect 20456 33844 20484 34020
rect 20806 33940 20812 33992
rect 20864 33980 20870 33992
rect 24581 33983 24639 33989
rect 24581 33980 24593 33983
rect 20864 33952 24593 33980
rect 20864 33940 20870 33952
rect 24581 33949 24593 33952
rect 24627 33980 24639 33983
rect 25222 33980 25228 33992
rect 24627 33952 25228 33980
rect 24627 33949 24639 33952
rect 24581 33943 24639 33949
rect 25222 33940 25228 33952
rect 25280 33940 25286 33992
rect 25406 33940 25412 33992
rect 25464 33980 25470 33992
rect 35866 33980 35894 34088
rect 38010 34076 38016 34088
rect 38068 34076 38074 34128
rect 25464 33952 35894 33980
rect 25464 33940 25470 33952
rect 20530 33872 20536 33924
rect 20588 33912 20594 33924
rect 20588 33884 22692 33912
rect 20588 33872 20594 33884
rect 20898 33844 20904 33856
rect 19306 33816 20484 33844
rect 20859 33816 20904 33844
rect 20898 33804 20904 33816
rect 20956 33804 20962 33856
rect 22094 33804 22100 33856
rect 22152 33844 22158 33856
rect 22557 33847 22615 33853
rect 22557 33844 22569 33847
rect 22152 33816 22569 33844
rect 22152 33804 22158 33816
rect 22557 33813 22569 33816
rect 22603 33813 22615 33847
rect 22664 33844 22692 33884
rect 22738 33872 22744 33924
rect 22796 33912 22802 33924
rect 25133 33915 25191 33921
rect 25133 33912 25145 33915
rect 22796 33884 25145 33912
rect 22796 33872 22802 33884
rect 25133 33881 25145 33884
rect 25179 33881 25191 33915
rect 25133 33875 25191 33881
rect 23658 33844 23664 33856
rect 22664 33816 23664 33844
rect 22557 33807 22615 33813
rect 23658 33804 23664 33816
rect 23716 33804 23722 33856
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 3053 33643 3111 33649
rect 3053 33609 3065 33643
rect 3099 33640 3111 33643
rect 3099 33612 11376 33640
rect 3099 33609 3111 33612
rect 3053 33603 3111 33609
rect 2774 33572 2780 33584
rect 2424 33544 2780 33572
rect 1026 33464 1032 33516
rect 1084 33504 1090 33516
rect 2424 33513 2452 33544
rect 2774 33532 2780 33544
rect 2832 33532 2838 33584
rect 4614 33532 4620 33584
rect 4672 33532 4678 33584
rect 5261 33575 5319 33581
rect 5261 33541 5273 33575
rect 5307 33572 5319 33575
rect 5902 33572 5908 33584
rect 5307 33544 5908 33572
rect 5307 33541 5319 33544
rect 5261 33535 5319 33541
rect 5902 33532 5908 33544
rect 5960 33532 5966 33584
rect 7282 33532 7288 33584
rect 7340 33572 7346 33584
rect 7340 33544 7385 33572
rect 7340 33532 7346 33544
rect 7926 33532 7932 33584
rect 7984 33532 7990 33584
rect 11348 33572 11376 33612
rect 11422 33600 11428 33652
rect 11480 33640 11486 33652
rect 14366 33640 14372 33652
rect 11480 33612 14372 33640
rect 11480 33600 11486 33612
rect 14366 33600 14372 33612
rect 14424 33600 14430 33652
rect 14458 33600 14464 33652
rect 14516 33640 14522 33652
rect 19242 33640 19248 33652
rect 14516 33612 19248 33640
rect 14516 33600 14522 33612
rect 19242 33600 19248 33612
rect 19300 33600 19306 33652
rect 19426 33600 19432 33652
rect 19484 33640 19490 33652
rect 19521 33643 19579 33649
rect 19521 33640 19533 33643
rect 19484 33612 19533 33640
rect 19484 33600 19490 33612
rect 19521 33609 19533 33612
rect 19567 33609 19579 33643
rect 19521 33603 19579 33609
rect 22649 33643 22707 33649
rect 22649 33609 22661 33643
rect 22695 33640 22707 33643
rect 23198 33640 23204 33652
rect 22695 33612 23204 33640
rect 22695 33609 22707 33612
rect 22649 33603 22707 33609
rect 23198 33600 23204 33612
rect 23256 33600 23262 33652
rect 25222 33600 25228 33652
rect 25280 33640 25286 33652
rect 25317 33643 25375 33649
rect 25317 33640 25329 33643
rect 25280 33612 25329 33640
rect 25280 33600 25286 33612
rect 25317 33609 25329 33612
rect 25363 33609 25375 33643
rect 25317 33603 25375 33609
rect 12250 33572 12256 33584
rect 11348 33544 12256 33572
rect 12250 33532 12256 33544
rect 12308 33532 12314 33584
rect 13446 33572 13452 33584
rect 13202 33544 13452 33572
rect 13446 33532 13452 33544
rect 13504 33532 13510 33584
rect 13538 33532 13544 33584
rect 13596 33572 13602 33584
rect 15838 33572 15844 33584
rect 13596 33544 15844 33572
rect 13596 33532 13602 33544
rect 15838 33532 15844 33544
rect 15896 33532 15902 33584
rect 16022 33572 16028 33584
rect 15983 33544 16028 33572
rect 16022 33532 16028 33544
rect 16080 33532 16086 33584
rect 16117 33575 16175 33581
rect 16117 33541 16129 33575
rect 16163 33572 16175 33575
rect 17494 33572 17500 33584
rect 16163 33544 17500 33572
rect 16163 33541 16175 33544
rect 16117 33535 16175 33541
rect 17494 33532 17500 33544
rect 17552 33532 17558 33584
rect 17862 33532 17868 33584
rect 17920 33572 17926 33584
rect 20806 33572 20812 33584
rect 17920 33544 20812 33572
rect 17920 33532 17926 33544
rect 2409 33507 2467 33513
rect 2409 33504 2421 33507
rect 1084 33476 2421 33504
rect 1084 33464 1090 33476
rect 2409 33473 2421 33476
rect 2455 33473 2467 33507
rect 2409 33467 2467 33473
rect 2866 33464 2872 33516
rect 2924 33504 2930 33516
rect 2961 33507 3019 33513
rect 2961 33504 2973 33507
rect 2924 33476 2973 33504
rect 2924 33464 2930 33476
rect 2961 33473 2973 33476
rect 3007 33473 3019 33507
rect 2961 33467 3019 33473
rect 3418 33464 3424 33516
rect 3476 33504 3482 33516
rect 3476 33476 4108 33504
rect 3476 33464 3482 33476
rect 2133 33439 2191 33445
rect 2133 33405 2145 33439
rect 2179 33405 2191 33439
rect 4080 33436 4108 33476
rect 5534 33464 5540 33516
rect 5592 33504 5598 33516
rect 7009 33507 7067 33513
rect 7009 33504 7021 33507
rect 5592 33476 7021 33504
rect 5592 33464 5598 33476
rect 7009 33473 7021 33476
rect 7055 33473 7067 33507
rect 9306 33504 9312 33516
rect 9267 33476 9312 33504
rect 7009 33467 7067 33473
rect 9306 33464 9312 33476
rect 9364 33464 9370 33516
rect 10718 33476 11008 33504
rect 9585 33439 9643 33445
rect 9585 33436 9597 33439
rect 4080 33408 9597 33436
rect 2133 33399 2191 33405
rect 9585 33405 9597 33408
rect 9631 33405 9643 33439
rect 9585 33399 9643 33405
rect 2148 33368 2176 33399
rect 9674 33396 9680 33448
rect 9732 33436 9738 33448
rect 9950 33436 9956 33448
rect 9732 33408 9956 33436
rect 9732 33396 9738 33408
rect 9950 33396 9956 33408
rect 10008 33396 10014 33448
rect 10980 33368 11008 33476
rect 11054 33464 11060 33516
rect 11112 33504 11118 33516
rect 11701 33507 11759 33513
rect 11701 33504 11713 33507
rect 11112 33476 11713 33504
rect 11112 33464 11118 33476
rect 11701 33473 11713 33476
rect 11747 33473 11759 33507
rect 11701 33467 11759 33473
rect 14366 33464 14372 33516
rect 14424 33504 14430 33516
rect 14645 33507 14703 33513
rect 14645 33504 14657 33507
rect 14424 33476 14657 33504
rect 14424 33464 14430 33476
rect 14645 33473 14657 33476
rect 14691 33473 14703 33507
rect 14645 33467 14703 33473
rect 11974 33436 11980 33448
rect 11935 33408 11980 33436
rect 11974 33396 11980 33408
rect 12032 33396 12038 33448
rect 13170 33396 13176 33448
rect 13228 33436 13234 33448
rect 13725 33439 13783 33445
rect 13725 33436 13737 33439
rect 13228 33408 13737 33436
rect 13228 33396 13234 33408
rect 13725 33405 13737 33408
rect 13771 33405 13783 33439
rect 13725 33399 13783 33405
rect 14660 33368 14688 33467
rect 16666 33464 16672 33516
rect 16724 33504 16730 33516
rect 16853 33507 16911 33513
rect 16853 33504 16865 33507
rect 16724 33476 16865 33504
rect 16724 33464 16730 33476
rect 16853 33473 16865 33476
rect 16899 33473 16911 33507
rect 17954 33504 17960 33516
rect 17915 33476 17960 33504
rect 16853 33467 16911 33473
rect 17954 33464 17960 33476
rect 18012 33464 18018 33516
rect 18966 33504 18972 33516
rect 18879 33476 18972 33504
rect 18966 33464 18972 33476
rect 19024 33504 19030 33516
rect 19334 33504 19340 33516
rect 19024 33476 19340 33504
rect 19024 33464 19030 33476
rect 19334 33464 19340 33476
rect 19392 33464 19398 33516
rect 19628 33513 19656 33544
rect 20806 33532 20812 33544
rect 20864 33572 20870 33584
rect 21085 33575 21143 33581
rect 21085 33572 21097 33575
rect 20864 33544 21097 33572
rect 20864 33532 20870 33544
rect 21085 33541 21097 33544
rect 21131 33541 21143 33575
rect 21085 33535 21143 33541
rect 19613 33507 19671 33513
rect 19613 33473 19625 33507
rect 19659 33473 19671 33507
rect 20622 33504 20628 33516
rect 20583 33476 20628 33504
rect 19613 33467 19671 33473
rect 20622 33464 20628 33476
rect 20680 33464 20686 33516
rect 22830 33464 22836 33516
rect 22888 33504 22894 33516
rect 24857 33507 24915 33513
rect 24857 33504 24869 33507
rect 22888 33476 24869 33504
rect 22888 33464 22894 33476
rect 24857 33473 24869 33476
rect 24903 33473 24915 33507
rect 26418 33504 26424 33516
rect 26379 33476 26424 33504
rect 24857 33467 24915 33473
rect 26418 33464 26424 33476
rect 26476 33464 26482 33516
rect 37553 33507 37611 33513
rect 37553 33473 37565 33507
rect 37599 33504 37611 33507
rect 38194 33504 38200 33516
rect 37599 33476 38200 33504
rect 37599 33473 37611 33476
rect 37553 33467 37611 33473
rect 38194 33464 38200 33476
rect 38252 33464 38258 33516
rect 15838 33436 15844 33448
rect 15799 33408 15844 33436
rect 15838 33396 15844 33408
rect 15896 33396 15902 33448
rect 15930 33396 15936 33448
rect 15988 33436 15994 33448
rect 18877 33439 18935 33445
rect 18877 33436 18889 33439
rect 15988 33424 16804 33436
rect 17052 33424 18889 33436
rect 15988 33408 18889 33424
rect 15988 33396 15994 33408
rect 16776 33396 17080 33408
rect 18877 33405 18889 33408
rect 18923 33405 18935 33439
rect 18877 33399 18935 33405
rect 20714 33396 20720 33448
rect 20772 33436 20778 33448
rect 23661 33439 23719 33445
rect 23661 33436 23673 33439
rect 20772 33408 23673 33436
rect 20772 33396 20778 33408
rect 23661 33405 23673 33408
rect 23707 33405 23719 33439
rect 23661 33399 23719 33405
rect 2148 33340 4016 33368
rect 3786 33300 3792 33312
rect 3747 33272 3792 33300
rect 3786 33260 3792 33272
rect 3844 33260 3850 33312
rect 3988 33300 4016 33340
rect 8680 33340 9444 33368
rect 10980 33340 11560 33368
rect 14660 33340 15516 33368
rect 7834 33300 7840 33312
rect 3988 33272 7840 33300
rect 7834 33260 7840 33272
rect 7892 33260 7898 33312
rect 7926 33260 7932 33312
rect 7984 33300 7990 33312
rect 8680 33300 8708 33340
rect 7984 33272 8708 33300
rect 8757 33303 8815 33309
rect 7984 33260 7990 33272
rect 8757 33269 8769 33303
rect 8803 33300 8815 33303
rect 9306 33300 9312 33312
rect 8803 33272 9312 33300
rect 8803 33269 8815 33272
rect 8757 33263 8815 33269
rect 9306 33260 9312 33272
rect 9364 33260 9370 33312
rect 9416 33300 9444 33340
rect 11057 33303 11115 33309
rect 11057 33300 11069 33303
rect 9416 33272 11069 33300
rect 11057 33269 11069 33272
rect 11103 33300 11115 33303
rect 11330 33300 11336 33312
rect 11103 33272 11336 33300
rect 11103 33269 11115 33272
rect 11057 33263 11115 33269
rect 11330 33260 11336 33272
rect 11388 33260 11394 33312
rect 11532 33300 11560 33340
rect 14458 33300 14464 33312
rect 11532 33272 14464 33300
rect 14458 33260 14464 33272
rect 14516 33260 14522 33312
rect 14553 33303 14611 33309
rect 14553 33269 14565 33303
rect 14599 33300 14611 33303
rect 14734 33300 14740 33312
rect 14599 33272 14740 33300
rect 14599 33269 14611 33272
rect 14553 33263 14611 33269
rect 14734 33260 14740 33272
rect 14792 33260 14798 33312
rect 15488 33300 15516 33340
rect 15562 33328 15568 33380
rect 15620 33368 15626 33380
rect 20533 33371 20591 33377
rect 20533 33368 20545 33371
rect 15620 33340 20545 33368
rect 15620 33328 15626 33340
rect 20533 33337 20545 33340
rect 20579 33337 20591 33371
rect 23109 33371 23167 33377
rect 23109 33368 23121 33371
rect 20533 33331 20591 33337
rect 22112 33340 23121 33368
rect 22112 33312 22140 33340
rect 23109 33337 23121 33340
rect 23155 33337 23167 33371
rect 25866 33368 25872 33380
rect 25827 33340 25872 33368
rect 23109 33331 23167 33337
rect 25866 33328 25872 33340
rect 25924 33328 25930 33380
rect 37366 33328 37372 33380
rect 37424 33368 37430 33380
rect 38013 33371 38071 33377
rect 38013 33368 38025 33371
rect 37424 33340 38025 33368
rect 37424 33328 37430 33340
rect 38013 33337 38025 33340
rect 38059 33337 38071 33371
rect 38013 33331 38071 33337
rect 16482 33300 16488 33312
rect 15488 33272 16488 33300
rect 16482 33260 16488 33272
rect 16540 33260 16546 33312
rect 16945 33303 17003 33309
rect 16945 33269 16957 33303
rect 16991 33300 17003 33303
rect 17862 33300 17868 33312
rect 16991 33272 17868 33300
rect 16991 33269 17003 33272
rect 16945 33263 17003 33269
rect 17862 33260 17868 33272
rect 17920 33260 17926 33312
rect 18049 33303 18107 33309
rect 18049 33269 18061 33303
rect 18095 33300 18107 33303
rect 18598 33300 18604 33312
rect 18095 33272 18604 33300
rect 18095 33269 18107 33272
rect 18049 33263 18107 33269
rect 18598 33260 18604 33272
rect 18656 33260 18662 33312
rect 22094 33260 22100 33312
rect 22152 33300 22158 33312
rect 22152 33272 22197 33300
rect 22152 33260 22158 33272
rect 24026 33260 24032 33312
rect 24084 33300 24090 33312
rect 24213 33303 24271 33309
rect 24213 33300 24225 33303
rect 24084 33272 24225 33300
rect 24084 33260 24090 33272
rect 24213 33269 24225 33272
rect 24259 33269 24271 33303
rect 24213 33263 24271 33269
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 1936 33099 1994 33105
rect 1936 33065 1948 33099
rect 1982 33096 1994 33099
rect 3326 33096 3332 33108
rect 1982 33068 3332 33096
rect 1982 33065 1994 33068
rect 1936 33059 1994 33065
rect 3326 33056 3332 33068
rect 3384 33056 3390 33108
rect 3421 33099 3479 33105
rect 3421 33065 3433 33099
rect 3467 33096 3479 33099
rect 7006 33096 7012 33108
rect 3467 33068 7012 33096
rect 3467 33065 3479 33068
rect 3421 33059 3479 33065
rect 7006 33056 7012 33068
rect 7064 33056 7070 33108
rect 7282 33056 7288 33108
rect 7340 33096 7346 33108
rect 11146 33096 11152 33108
rect 7340 33068 11152 33096
rect 7340 33056 7346 33068
rect 11146 33056 11152 33068
rect 11204 33056 11210 33108
rect 16390 33096 16396 33108
rect 11348 33068 16396 33096
rect 5534 32988 5540 33040
rect 5592 32988 5598 33040
rect 7098 32988 7104 33040
rect 7156 33028 7162 33040
rect 11348 33028 11376 33068
rect 16390 33056 16396 33068
rect 16448 33056 16454 33108
rect 16574 33056 16580 33108
rect 16632 33096 16638 33108
rect 17402 33096 17408 33108
rect 16632 33068 17408 33096
rect 16632 33056 16638 33068
rect 17402 33056 17408 33068
rect 17460 33056 17466 33108
rect 19242 33056 19248 33108
rect 19300 33096 19306 33108
rect 19521 33099 19579 33105
rect 19521 33096 19533 33099
rect 19300 33068 19533 33096
rect 19300 33056 19306 33068
rect 19521 33065 19533 33068
rect 19567 33065 19579 33099
rect 19521 33059 19579 33065
rect 20717 33099 20775 33105
rect 20717 33065 20729 33099
rect 20763 33096 20775 33099
rect 20898 33096 20904 33108
rect 20763 33068 20904 33096
rect 20763 33065 20775 33068
rect 20717 33059 20775 33065
rect 20898 33056 20904 33068
rect 20956 33056 20962 33108
rect 21726 33096 21732 33108
rect 21687 33068 21732 33096
rect 21726 33056 21732 33068
rect 21784 33056 21790 33108
rect 22925 33099 22983 33105
rect 22925 33065 22937 33099
rect 22971 33096 22983 33099
rect 23198 33096 23204 33108
rect 22971 33068 23204 33096
rect 22971 33065 22983 33068
rect 22925 33059 22983 33065
rect 23198 33056 23204 33068
rect 23256 33056 23262 33108
rect 23477 33099 23535 33105
rect 23477 33065 23489 33099
rect 23523 33096 23535 33099
rect 23658 33096 23664 33108
rect 23523 33068 23664 33096
rect 23523 33065 23535 33068
rect 23477 33059 23535 33065
rect 23658 33056 23664 33068
rect 23716 33056 23722 33108
rect 25222 33096 25228 33108
rect 25183 33068 25228 33096
rect 25222 33056 25228 33068
rect 25280 33056 25286 33108
rect 7156 33000 11376 33028
rect 7156 32988 7162 33000
rect 12618 32988 12624 33040
rect 12676 33028 12682 33040
rect 22186 33028 22192 33040
rect 12676 33000 22192 33028
rect 12676 32988 12682 33000
rect 22186 32988 22192 33000
rect 22244 32988 22250 33040
rect 1673 32963 1731 32969
rect 1673 32929 1685 32963
rect 1719 32960 1731 32963
rect 2958 32960 2964 32972
rect 1719 32932 2964 32960
rect 1719 32929 1731 32932
rect 1673 32923 1731 32929
rect 2958 32920 2964 32932
rect 3016 32920 3022 32972
rect 4893 32963 4951 32969
rect 4893 32929 4905 32963
rect 4939 32960 4951 32963
rect 5442 32960 5448 32972
rect 4939 32932 5448 32960
rect 4939 32929 4951 32932
rect 4893 32923 4951 32929
rect 5442 32920 5448 32932
rect 5500 32920 5506 32972
rect 5552 32960 5580 32988
rect 6917 32963 6975 32969
rect 6917 32960 6929 32963
rect 5552 32932 6929 32960
rect 6917 32929 6929 32932
rect 6963 32929 6975 32963
rect 6917 32923 6975 32929
rect 7282 32920 7288 32972
rect 7340 32960 7346 32972
rect 7340 32932 10640 32960
rect 7340 32920 7346 32932
rect 4249 32895 4307 32901
rect 4249 32861 4261 32895
rect 4295 32892 4307 32895
rect 4982 32892 4988 32904
rect 4295 32864 4988 32892
rect 4295 32861 4307 32864
rect 4249 32855 4307 32861
rect 4982 32852 4988 32864
rect 5040 32852 5046 32904
rect 7466 32852 7472 32904
rect 7524 32892 7530 32904
rect 7745 32895 7803 32901
rect 7745 32892 7757 32895
rect 7524 32864 7757 32892
rect 7524 32852 7530 32864
rect 7745 32861 7757 32864
rect 7791 32892 7803 32895
rect 8294 32892 8300 32904
rect 7791 32864 8300 32892
rect 7791 32861 7803 32864
rect 7745 32855 7803 32861
rect 8294 32852 8300 32864
rect 8352 32852 8358 32904
rect 8573 32895 8631 32901
rect 8573 32861 8585 32895
rect 8619 32892 8631 32895
rect 8846 32892 8852 32904
rect 8619 32864 8852 32892
rect 8619 32861 8631 32864
rect 8573 32855 8631 32861
rect 8846 32852 8852 32864
rect 8904 32892 8910 32904
rect 9125 32895 9183 32901
rect 9125 32892 9137 32895
rect 8904 32864 9137 32892
rect 8904 32852 8910 32864
rect 9125 32861 9137 32864
rect 9171 32861 9183 32895
rect 9125 32855 9183 32861
rect 9306 32852 9312 32904
rect 9364 32892 9370 32904
rect 10612 32901 10640 32932
rect 11054 32920 11060 32972
rect 11112 32960 11118 32972
rect 11241 32963 11299 32969
rect 11241 32960 11253 32963
rect 11112 32932 11253 32960
rect 11112 32920 11118 32932
rect 11241 32929 11253 32932
rect 11287 32929 11299 32963
rect 11514 32960 11520 32972
rect 11475 32932 11520 32960
rect 11241 32923 11299 32929
rect 11514 32920 11520 32932
rect 11572 32960 11578 32972
rect 12158 32960 12164 32972
rect 11572 32932 12164 32960
rect 11572 32920 11578 32932
rect 12158 32920 12164 32932
rect 12216 32920 12222 32972
rect 13446 32920 13452 32972
rect 13504 32960 13510 32972
rect 14274 32960 14280 32972
rect 13504 32932 14280 32960
rect 13504 32920 13510 32932
rect 14274 32920 14280 32932
rect 14332 32920 14338 32972
rect 15565 32963 15623 32969
rect 15565 32929 15577 32963
rect 15611 32960 15623 32963
rect 16114 32960 16120 32972
rect 15611 32932 16120 32960
rect 15611 32929 15623 32932
rect 15565 32923 15623 32929
rect 16114 32920 16120 32932
rect 16172 32960 16178 32972
rect 16574 32960 16580 32972
rect 16172 32932 16580 32960
rect 16172 32920 16178 32932
rect 16574 32920 16580 32932
rect 16632 32920 16638 32972
rect 16942 32960 16948 32972
rect 16903 32932 16948 32960
rect 16942 32920 16948 32932
rect 17000 32920 17006 32972
rect 17218 32920 17224 32972
rect 17276 32960 17282 32972
rect 20714 32960 20720 32972
rect 17276 32932 20720 32960
rect 17276 32920 17282 32932
rect 20714 32920 20720 32932
rect 20772 32920 20778 32972
rect 9861 32895 9919 32901
rect 9861 32892 9873 32895
rect 9364 32864 9873 32892
rect 9364 32852 9370 32864
rect 9861 32861 9873 32864
rect 9907 32861 9919 32895
rect 9861 32855 9919 32861
rect 10597 32895 10655 32901
rect 10597 32861 10609 32895
rect 10643 32861 10655 32895
rect 10597 32855 10655 32861
rect 12618 32852 12624 32904
rect 12676 32852 12682 32904
rect 13354 32852 13360 32904
rect 13412 32892 13418 32904
rect 14369 32895 14427 32901
rect 14369 32892 14381 32895
rect 13412 32864 14381 32892
rect 13412 32852 13418 32864
rect 14369 32861 14381 32864
rect 14415 32892 14427 32895
rect 14642 32892 14648 32904
rect 14415 32864 14648 32892
rect 14415 32861 14427 32864
rect 14369 32855 14427 32861
rect 14642 32852 14648 32864
rect 14700 32852 14706 32904
rect 18322 32892 18328 32904
rect 18283 32864 18328 32892
rect 18322 32852 18328 32864
rect 18380 32852 18386 32904
rect 19334 32852 19340 32904
rect 19392 32892 19398 32904
rect 19613 32895 19671 32901
rect 19613 32892 19625 32895
rect 19392 32864 19625 32892
rect 19392 32852 19398 32864
rect 19613 32861 19625 32864
rect 19659 32861 19671 32895
rect 19613 32855 19671 32861
rect 20622 32852 20628 32904
rect 20680 32892 20686 32904
rect 21821 32895 21879 32901
rect 21821 32892 21833 32895
rect 20680 32864 21833 32892
rect 20680 32852 20686 32864
rect 21821 32861 21833 32864
rect 21867 32892 21879 32895
rect 22278 32892 22284 32904
rect 21867 32864 22284 32892
rect 21867 32861 21879 32864
rect 21821 32855 21879 32861
rect 22278 32852 22284 32864
rect 22336 32852 22342 32904
rect 25682 32892 25688 32904
rect 25643 32864 25688 32892
rect 25682 32852 25688 32864
rect 25740 32852 25746 32904
rect 2056 32796 2438 32824
rect 1210 32716 1216 32768
rect 1268 32756 1274 32768
rect 2056 32756 2084 32796
rect 5626 32784 5632 32836
rect 5684 32784 5690 32836
rect 6638 32824 6644 32836
rect 6599 32796 6644 32824
rect 6638 32784 6644 32796
rect 6696 32784 6702 32836
rect 9953 32827 10011 32833
rect 9953 32793 9965 32827
rect 9999 32824 10011 32827
rect 11422 32824 11428 32836
rect 9999 32796 11428 32824
rect 9999 32793 10011 32796
rect 9953 32787 10011 32793
rect 11422 32784 11428 32796
rect 11480 32784 11486 32836
rect 13262 32824 13268 32836
rect 13223 32796 13268 32824
rect 13262 32784 13268 32796
rect 13320 32784 13326 32836
rect 14200 32796 14504 32824
rect 1268 32728 2084 32756
rect 4341 32759 4399 32765
rect 1268 32716 1274 32728
rect 4341 32725 4353 32759
rect 4387 32756 4399 32759
rect 5994 32756 6000 32768
rect 4387 32728 6000 32756
rect 4387 32725 4399 32728
rect 4341 32719 4399 32725
rect 5994 32716 6000 32728
rect 6052 32716 6058 32768
rect 7653 32759 7711 32765
rect 7653 32725 7665 32759
rect 7699 32756 7711 32759
rect 7742 32756 7748 32768
rect 7699 32728 7748 32756
rect 7699 32725 7711 32728
rect 7653 32719 7711 32725
rect 7742 32716 7748 32728
rect 7800 32716 7806 32768
rect 8478 32756 8484 32768
rect 8439 32728 8484 32756
rect 8478 32716 8484 32728
rect 8536 32716 8542 32768
rect 9214 32756 9220 32768
rect 9175 32728 9220 32756
rect 9214 32716 9220 32728
rect 9272 32716 9278 32768
rect 9490 32716 9496 32768
rect 9548 32756 9554 32768
rect 10502 32756 10508 32768
rect 9548 32728 10508 32756
rect 9548 32716 9554 32728
rect 10502 32716 10508 32728
rect 10560 32716 10566 32768
rect 10686 32756 10692 32768
rect 10647 32728 10692 32756
rect 10686 32716 10692 32728
rect 10744 32716 10750 32768
rect 12250 32716 12256 32768
rect 12308 32756 12314 32768
rect 14200 32756 14228 32796
rect 12308 32728 14228 32756
rect 14476 32756 14504 32796
rect 14734 32784 14740 32836
rect 14792 32824 14798 32836
rect 14921 32827 14979 32833
rect 14921 32824 14933 32827
rect 14792 32796 14933 32824
rect 14792 32784 14798 32796
rect 14921 32793 14933 32796
rect 14967 32793 14979 32827
rect 14921 32787 14979 32793
rect 15013 32827 15071 32833
rect 15013 32793 15025 32827
rect 15059 32824 15071 32827
rect 16390 32824 16396 32836
rect 15059 32796 16396 32824
rect 15059 32793 15071 32796
rect 15013 32787 15071 32793
rect 16390 32784 16396 32796
rect 16448 32784 16454 32836
rect 16669 32827 16727 32833
rect 16669 32793 16681 32827
rect 16715 32793 16727 32827
rect 16669 32787 16727 32793
rect 16574 32756 16580 32768
rect 14476 32728 16580 32756
rect 12308 32716 12314 32728
rect 16574 32716 16580 32728
rect 16632 32716 16638 32768
rect 16684 32756 16712 32787
rect 16758 32784 16764 32836
rect 16816 32824 16822 32836
rect 20070 32824 20076 32836
rect 16816 32796 20076 32824
rect 16816 32784 16822 32796
rect 20070 32784 20076 32796
rect 20128 32784 20134 32836
rect 17034 32756 17040 32768
rect 16684 32728 17040 32756
rect 17034 32716 17040 32728
rect 17092 32716 17098 32768
rect 18417 32759 18475 32765
rect 18417 32725 18429 32759
rect 18463 32756 18475 32759
rect 18506 32756 18512 32768
rect 18463 32728 18512 32756
rect 18463 32725 18475 32728
rect 18417 32719 18475 32725
rect 18506 32716 18512 32728
rect 18564 32716 18570 32768
rect 20165 32759 20223 32765
rect 20165 32725 20177 32759
rect 20211 32756 20223 32759
rect 20346 32756 20352 32768
rect 20211 32728 20352 32756
rect 20211 32725 20223 32728
rect 20165 32719 20223 32725
rect 20346 32716 20352 32728
rect 20404 32716 20410 32768
rect 22094 32716 22100 32768
rect 22152 32756 22158 32768
rect 22281 32759 22339 32765
rect 22281 32756 22293 32759
rect 22152 32728 22293 32756
rect 22152 32716 22158 32728
rect 22281 32725 22293 32728
rect 22327 32725 22339 32759
rect 24026 32756 24032 32768
rect 23987 32728 24032 32756
rect 22281 32719 22339 32725
rect 24026 32716 24032 32728
rect 24084 32756 24090 32768
rect 24581 32759 24639 32765
rect 24581 32756 24593 32759
rect 24084 32728 24593 32756
rect 24084 32716 24090 32728
rect 24581 32725 24593 32728
rect 24627 32725 24639 32759
rect 24581 32719 24639 32725
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 1765 32555 1823 32561
rect 1765 32521 1777 32555
rect 1811 32552 1823 32555
rect 1811 32524 2774 32552
rect 1811 32521 1823 32524
rect 1765 32515 1823 32521
rect 1670 32416 1676 32428
rect 1631 32388 1676 32416
rect 1670 32376 1676 32388
rect 1728 32376 1734 32428
rect 2590 32416 2596 32428
rect 2551 32388 2596 32416
rect 2590 32376 2596 32388
rect 2648 32376 2654 32428
rect 2746 32348 2774 32524
rect 2958 32512 2964 32564
rect 3016 32552 3022 32564
rect 3053 32555 3111 32561
rect 3053 32552 3065 32555
rect 3016 32524 3065 32552
rect 3016 32512 3022 32524
rect 3053 32521 3065 32524
rect 3099 32521 3111 32555
rect 5074 32552 5080 32564
rect 3053 32515 3111 32521
rect 3160 32524 5080 32552
rect 2866 32444 2872 32496
rect 2924 32484 2930 32496
rect 3160 32484 3188 32524
rect 5074 32512 5080 32524
rect 5132 32512 5138 32564
rect 5534 32512 5540 32564
rect 5592 32552 5598 32564
rect 5905 32555 5963 32561
rect 5905 32552 5917 32555
rect 5592 32524 5917 32552
rect 5592 32512 5598 32524
rect 5905 32521 5917 32524
rect 5951 32521 5963 32555
rect 5905 32515 5963 32521
rect 7006 32512 7012 32564
rect 7064 32552 7070 32564
rect 11793 32555 11851 32561
rect 7064 32524 9720 32552
rect 7064 32512 7070 32524
rect 2924 32456 3188 32484
rect 2924 32444 2930 32456
rect 3510 32444 3516 32496
rect 3568 32484 3574 32496
rect 3568 32456 4002 32484
rect 3568 32444 3574 32456
rect 5445 32419 5503 32425
rect 5445 32385 5457 32419
rect 5491 32416 5503 32419
rect 5552 32416 5580 32512
rect 7742 32444 7748 32496
rect 7800 32444 7806 32496
rect 8481 32487 8539 32493
rect 8481 32453 8493 32487
rect 8527 32484 8539 32487
rect 9030 32484 9036 32496
rect 8527 32456 9036 32484
rect 8527 32453 8539 32456
rect 8481 32447 8539 32453
rect 9030 32444 9036 32456
rect 9088 32444 9094 32496
rect 9692 32493 9720 32524
rect 11793 32521 11805 32555
rect 11839 32552 11851 32555
rect 12894 32552 12900 32564
rect 11839 32524 12900 32552
rect 11839 32521 11851 32524
rect 11793 32515 11851 32521
rect 9677 32487 9735 32493
rect 9677 32453 9689 32487
rect 9723 32453 9735 32487
rect 11606 32484 11612 32496
rect 10902 32456 11612 32484
rect 9677 32447 9735 32453
rect 11606 32444 11612 32456
rect 11664 32444 11670 32496
rect 5491 32388 5580 32416
rect 5491 32385 5503 32388
rect 5445 32379 5503 32385
rect 11146 32376 11152 32428
rect 11204 32416 11210 32428
rect 11808 32416 11836 32515
rect 12894 32512 12900 32524
rect 12952 32512 12958 32564
rect 15378 32512 15384 32564
rect 15436 32552 15442 32564
rect 16850 32552 16856 32564
rect 15436 32524 16856 32552
rect 15436 32512 15442 32524
rect 16850 32512 16856 32524
rect 16908 32512 16914 32564
rect 20165 32555 20223 32561
rect 20165 32552 20177 32555
rect 17604 32524 20177 32552
rect 12986 32444 12992 32496
rect 13044 32484 13050 32496
rect 13044 32456 13584 32484
rect 13044 32444 13050 32456
rect 11204 32388 11836 32416
rect 11204 32376 11210 32388
rect 2746 32320 3832 32348
rect 2314 32240 2320 32292
rect 2372 32280 2378 32292
rect 2409 32283 2467 32289
rect 2409 32280 2421 32283
rect 2372 32252 2421 32280
rect 2372 32240 2378 32252
rect 2409 32249 2421 32252
rect 2455 32249 2467 32283
rect 3694 32280 3700 32292
rect 3655 32252 3700 32280
rect 2409 32243 2467 32249
rect 3694 32240 3700 32252
rect 3752 32240 3758 32292
rect 3804 32212 3832 32320
rect 3878 32308 3884 32360
rect 3936 32348 3942 32360
rect 5169 32351 5227 32357
rect 5169 32348 5181 32351
rect 3936 32320 5181 32348
rect 3936 32308 3942 32320
rect 5169 32317 5181 32320
rect 5215 32317 5227 32351
rect 5169 32311 5227 32317
rect 6733 32351 6791 32357
rect 6733 32317 6745 32351
rect 6779 32348 6791 32351
rect 8386 32348 8392 32360
rect 6779 32320 8392 32348
rect 6779 32317 6791 32320
rect 6733 32311 6791 32317
rect 8386 32308 8392 32320
rect 8444 32308 8450 32360
rect 8754 32348 8760 32360
rect 8715 32320 8760 32348
rect 8754 32308 8760 32320
rect 8812 32348 8818 32360
rect 9398 32348 9404 32360
rect 8812 32320 9404 32348
rect 8812 32308 8818 32320
rect 9398 32308 9404 32320
rect 9456 32308 9462 32360
rect 12066 32348 12072 32360
rect 10704 32320 12072 32348
rect 5442 32240 5448 32292
rect 5500 32280 5506 32292
rect 7098 32280 7104 32292
rect 5500 32252 7104 32280
rect 5500 32240 5506 32252
rect 7098 32240 7104 32252
rect 7156 32240 7162 32292
rect 10704 32212 10732 32320
rect 12066 32308 12072 32320
rect 12124 32308 12130 32360
rect 11149 32283 11207 32289
rect 11149 32249 11161 32283
rect 11195 32280 11207 32283
rect 11514 32280 11520 32292
rect 11195 32252 11520 32280
rect 11195 32249 11207 32252
rect 11149 32243 11207 32249
rect 11514 32240 11520 32252
rect 11572 32240 11578 32292
rect 12176 32280 12204 32402
rect 12802 32308 12808 32360
rect 12860 32348 12866 32360
rect 13556 32357 13584 32456
rect 15102 32444 15108 32496
rect 15160 32444 15166 32496
rect 17405 32487 17463 32493
rect 17405 32453 17417 32487
rect 17451 32484 17463 32487
rect 17604 32484 17632 32524
rect 20165 32521 20177 32524
rect 20211 32521 20223 32555
rect 20165 32515 20223 32521
rect 22097 32555 22155 32561
rect 22097 32521 22109 32555
rect 22143 32552 22155 32555
rect 22186 32552 22192 32564
rect 22143 32524 22192 32552
rect 22143 32521 22155 32524
rect 22097 32515 22155 32521
rect 22186 32512 22192 32524
rect 22244 32512 22250 32564
rect 18322 32484 18328 32496
rect 17451 32456 17632 32484
rect 18283 32456 18328 32484
rect 17451 32453 17463 32456
rect 17405 32447 17463 32453
rect 18322 32444 18328 32456
rect 18380 32444 18386 32496
rect 18417 32487 18475 32493
rect 18417 32453 18429 32487
rect 18463 32484 18475 32487
rect 18690 32484 18696 32496
rect 18463 32456 18696 32484
rect 18463 32453 18475 32456
rect 18417 32447 18475 32453
rect 18690 32444 18696 32456
rect 18748 32444 18754 32496
rect 18782 32444 18788 32496
rect 18840 32484 18846 32496
rect 18969 32487 19027 32493
rect 18969 32484 18981 32487
rect 18840 32456 18981 32484
rect 18840 32444 18846 32456
rect 18969 32453 18981 32456
rect 19015 32453 19027 32487
rect 18969 32447 19027 32453
rect 19426 32376 19432 32428
rect 19484 32416 19490 32428
rect 19613 32419 19671 32425
rect 19613 32416 19625 32419
rect 19484 32388 19625 32416
rect 19484 32376 19490 32388
rect 19613 32385 19625 32388
rect 19659 32416 19671 32419
rect 19978 32416 19984 32428
rect 19659 32388 19984 32416
rect 19659 32385 19671 32388
rect 19613 32379 19671 32385
rect 19978 32376 19984 32388
rect 20036 32376 20042 32428
rect 20254 32416 20260 32428
rect 20167 32388 20260 32416
rect 20254 32376 20260 32388
rect 20312 32416 20318 32428
rect 20898 32416 20904 32428
rect 20312 32388 20904 32416
rect 20312 32376 20318 32388
rect 20898 32376 20904 32388
rect 20956 32376 20962 32428
rect 22186 32416 22192 32428
rect 22147 32388 22192 32416
rect 22186 32376 22192 32388
rect 22244 32376 22250 32428
rect 38010 32416 38016 32428
rect 37971 32388 38016 32416
rect 38010 32376 38016 32388
rect 38068 32376 38074 32428
rect 13265 32351 13323 32357
rect 13265 32348 13277 32351
rect 12860 32320 13277 32348
rect 12860 32308 12866 32320
rect 13265 32317 13277 32320
rect 13311 32317 13323 32351
rect 13265 32311 13323 32317
rect 13541 32351 13599 32357
rect 13541 32317 13553 32351
rect 13587 32348 13599 32351
rect 13587 32320 14596 32348
rect 13587 32317 13599 32320
rect 13541 32311 13599 32317
rect 11624 32252 12204 32280
rect 3804 32184 10732 32212
rect 10962 32172 10968 32224
rect 11020 32212 11026 32224
rect 11624 32212 11652 32252
rect 11020 32184 11652 32212
rect 11020 32172 11026 32184
rect 12066 32172 12072 32224
rect 12124 32212 12130 32224
rect 14093 32215 14151 32221
rect 14093 32212 14105 32215
rect 12124 32184 14105 32212
rect 12124 32172 12130 32184
rect 14093 32181 14105 32184
rect 14139 32181 14151 32215
rect 14568 32212 14596 32320
rect 15194 32308 15200 32360
rect 15252 32348 15258 32360
rect 15565 32351 15623 32357
rect 15565 32348 15577 32351
rect 15252 32320 15577 32348
rect 15252 32308 15258 32320
rect 15565 32317 15577 32320
rect 15611 32317 15623 32351
rect 15565 32311 15623 32317
rect 15841 32351 15899 32357
rect 15841 32317 15853 32351
rect 15887 32317 15899 32351
rect 17494 32348 17500 32360
rect 17455 32320 17500 32348
rect 15841 32311 15899 32317
rect 15856 32212 15884 32311
rect 17494 32308 17500 32320
rect 17552 32308 17558 32360
rect 17954 32308 17960 32360
rect 18012 32348 18018 32360
rect 19521 32351 19579 32357
rect 19521 32348 19533 32351
rect 18012 32320 19533 32348
rect 18012 32308 18018 32320
rect 19521 32317 19533 32320
rect 19567 32317 19579 32351
rect 20714 32348 20720 32360
rect 20675 32320 20720 32348
rect 19521 32311 19579 32317
rect 20714 32308 20720 32320
rect 20772 32308 20778 32360
rect 22094 32348 22100 32360
rect 22066 32308 22100 32348
rect 22152 32348 22158 32360
rect 22649 32351 22707 32357
rect 22649 32348 22661 32351
rect 22152 32320 22661 32348
rect 22152 32308 22158 32320
rect 22649 32317 22661 32320
rect 22695 32348 22707 32351
rect 23753 32351 23811 32357
rect 23753 32348 23765 32351
rect 22695 32320 23765 32348
rect 22695 32317 22707 32320
rect 22649 32311 22707 32317
rect 23753 32317 23765 32320
rect 23799 32348 23811 32351
rect 24026 32348 24032 32360
rect 23799 32320 24032 32348
rect 23799 32317 23811 32320
rect 23753 32311 23811 32317
rect 24026 32308 24032 32320
rect 24084 32348 24090 32360
rect 24305 32351 24363 32357
rect 24305 32348 24317 32351
rect 24084 32320 24317 32348
rect 24084 32308 24090 32320
rect 24305 32317 24317 32320
rect 24351 32317 24363 32351
rect 24305 32311 24363 32317
rect 16945 32283 17003 32289
rect 16945 32249 16957 32283
rect 16991 32280 17003 32283
rect 18414 32280 18420 32292
rect 16991 32252 18420 32280
rect 16991 32249 17003 32252
rect 16945 32243 17003 32249
rect 18414 32240 18420 32252
rect 18472 32240 18478 32292
rect 21361 32215 21419 32221
rect 21361 32212 21373 32215
rect 14568 32184 21373 32212
rect 14093 32175 14151 32181
rect 21361 32181 21373 32184
rect 21407 32212 21419 32215
rect 22066 32212 22094 32308
rect 21407 32184 22094 32212
rect 21407 32181 21419 32184
rect 21361 32175 21419 32181
rect 22278 32172 22284 32224
rect 22336 32212 22342 32224
rect 23201 32215 23259 32221
rect 23201 32212 23213 32215
rect 22336 32184 23213 32212
rect 22336 32172 22342 32184
rect 23201 32181 23213 32184
rect 23247 32181 23259 32215
rect 38194 32212 38200 32224
rect 38155 32184 38200 32212
rect 23201 32175 23259 32181
rect 38194 32172 38200 32184
rect 38252 32172 38258 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 1673 32011 1731 32017
rect 1673 31977 1685 32011
rect 1719 32008 1731 32011
rect 2774 32008 2780 32020
rect 1719 31980 2780 32008
rect 1719 31977 1731 31980
rect 1673 31971 1731 31977
rect 2774 31968 2780 31980
rect 2832 31968 2838 32020
rect 2958 31968 2964 32020
rect 3016 32008 3022 32020
rect 3418 32008 3424 32020
rect 3016 31980 3424 32008
rect 3016 31968 3022 31980
rect 3418 31968 3424 31980
rect 3476 31968 3482 32020
rect 4801 32011 4859 32017
rect 4801 31977 4813 32011
rect 4847 32008 4859 32011
rect 7098 32008 7104 32020
rect 4847 31980 7104 32008
rect 4847 31977 4859 31980
rect 4801 31971 4859 31977
rect 7098 31968 7104 31980
rect 7156 31968 7162 32020
rect 7282 31968 7288 32020
rect 7340 32008 7346 32020
rect 9306 32008 9312 32020
rect 7340 31980 9312 32008
rect 7340 31968 7346 31980
rect 9306 31968 9312 31980
rect 9364 31968 9370 32020
rect 10226 32008 10232 32020
rect 9508 31980 10232 32008
rect 7558 31900 7564 31952
rect 7616 31940 7622 31952
rect 9508 31949 9536 31980
rect 10226 31968 10232 31980
rect 10284 31968 10290 32020
rect 12066 32008 12072 32020
rect 10336 31980 12072 32008
rect 9493 31943 9551 31949
rect 7616 31912 9444 31940
rect 7616 31900 7622 31912
rect 3145 31875 3203 31881
rect 3145 31841 3157 31875
rect 3191 31872 3203 31875
rect 3602 31872 3608 31884
rect 3191 31844 3608 31872
rect 3191 31841 3203 31844
rect 3145 31835 3203 31841
rect 3602 31832 3608 31844
rect 3660 31832 3666 31884
rect 5534 31832 5540 31884
rect 5592 31872 5598 31884
rect 7377 31875 7435 31881
rect 7377 31872 7389 31875
rect 5592 31844 7389 31872
rect 5592 31832 5598 31844
rect 7377 31841 7389 31844
rect 7423 31872 7435 31875
rect 7837 31875 7895 31881
rect 7837 31872 7849 31875
rect 7423 31844 7849 31872
rect 7423 31841 7435 31844
rect 7377 31835 7435 31841
rect 7837 31841 7849 31844
rect 7883 31872 7895 31875
rect 8754 31872 8760 31884
rect 7883 31844 8760 31872
rect 7883 31841 7895 31844
rect 7837 31835 7895 31841
rect 8754 31832 8760 31844
rect 8812 31832 8818 31884
rect 3418 31764 3424 31816
rect 3476 31804 3482 31816
rect 4249 31807 4307 31813
rect 3476 31776 3521 31804
rect 3476 31764 3482 31776
rect 4249 31773 4261 31807
rect 4295 31804 4307 31807
rect 4709 31807 4767 31813
rect 4709 31804 4721 31807
rect 4295 31776 4721 31804
rect 4295 31773 4307 31776
rect 4249 31767 4307 31773
rect 4709 31773 4721 31776
rect 4755 31804 4767 31807
rect 5442 31804 5448 31816
rect 4755 31776 5448 31804
rect 4755 31773 4767 31776
rect 4709 31767 4767 31773
rect 5442 31764 5448 31776
rect 5500 31764 5506 31816
rect 5994 31764 6000 31816
rect 6052 31764 6058 31816
rect 8389 31807 8447 31813
rect 8389 31773 8401 31807
rect 8435 31773 8447 31807
rect 8389 31767 8447 31773
rect 8481 31807 8539 31813
rect 8481 31773 8493 31807
rect 8527 31804 8539 31807
rect 9306 31804 9312 31816
rect 8527 31776 9312 31804
rect 8527 31773 8539 31776
rect 8481 31767 8539 31773
rect 2130 31696 2136 31748
rect 2188 31696 2194 31748
rect 5353 31739 5411 31745
rect 5353 31705 5365 31739
rect 5399 31736 5411 31739
rect 5626 31736 5632 31748
rect 5399 31708 5632 31736
rect 5399 31705 5411 31708
rect 5353 31699 5411 31705
rect 5626 31696 5632 31708
rect 5684 31696 5690 31748
rect 7101 31739 7159 31745
rect 7101 31705 7113 31739
rect 7147 31736 7159 31739
rect 7190 31736 7196 31748
rect 7147 31708 7196 31736
rect 7147 31705 7159 31708
rect 7101 31699 7159 31705
rect 7190 31696 7196 31708
rect 7248 31696 7254 31748
rect 8404 31736 8432 31767
rect 9306 31764 9312 31776
rect 9364 31764 9370 31816
rect 9416 31813 9444 31912
rect 9493 31909 9505 31943
rect 9539 31909 9551 31943
rect 9493 31903 9551 31909
rect 10336 31872 10364 31980
rect 12066 31968 12072 31980
rect 12124 31968 12130 32020
rect 12434 31968 12440 32020
rect 12492 32008 12498 32020
rect 12989 32011 13047 32017
rect 12989 32008 13001 32011
rect 12492 31980 13001 32008
rect 12492 31968 12498 31980
rect 12989 31977 13001 31980
rect 13035 32008 13047 32011
rect 13446 32008 13452 32020
rect 13035 31980 13452 32008
rect 13035 31977 13047 31980
rect 12989 31971 13047 31977
rect 13446 31968 13452 31980
rect 13504 31968 13510 32020
rect 13538 31968 13544 32020
rect 13596 32008 13602 32020
rect 15378 32008 15384 32020
rect 13596 31980 15384 32008
rect 13596 31968 13602 31980
rect 15378 31968 15384 31980
rect 15436 31968 15442 32020
rect 15562 31968 15568 32020
rect 15620 32008 15626 32020
rect 19521 32011 19579 32017
rect 19521 32008 19533 32011
rect 15620 31980 19533 32008
rect 15620 31968 15626 31980
rect 19521 31977 19533 31980
rect 19567 31977 19579 32011
rect 19521 31971 19579 31977
rect 20806 31968 20812 32020
rect 20864 32008 20870 32020
rect 21729 32011 21787 32017
rect 21729 32008 21741 32011
rect 20864 31980 21741 32008
rect 20864 31968 20870 31980
rect 21729 31977 21741 31980
rect 21775 32008 21787 32011
rect 21818 32008 21824 32020
rect 21775 31980 21824 32008
rect 21775 31977 21787 31980
rect 21729 31971 21787 31977
rect 21818 31968 21824 31980
rect 21876 31968 21882 32020
rect 22094 31968 22100 32020
rect 22152 32008 22158 32020
rect 22281 32011 22339 32017
rect 22281 32008 22293 32011
rect 22152 31980 22293 32008
rect 22152 31968 22158 31980
rect 22281 31977 22293 31980
rect 22327 32008 22339 32011
rect 23385 32011 23443 32017
rect 23385 32008 23397 32011
rect 22327 31980 23397 32008
rect 22327 31977 22339 31980
rect 22281 31971 22339 31977
rect 23385 31977 23397 31980
rect 23431 31977 23443 32011
rect 23385 31971 23443 31977
rect 13630 31900 13636 31952
rect 13688 31940 13694 31952
rect 16022 31940 16028 31952
rect 13688 31912 13860 31940
rect 13688 31900 13694 31912
rect 10060 31844 10364 31872
rect 9401 31807 9459 31813
rect 9401 31773 9413 31807
rect 9447 31773 9459 31807
rect 9401 31767 9459 31773
rect 9582 31764 9588 31816
rect 9640 31804 9646 31816
rect 10060 31813 10088 31844
rect 10594 31832 10600 31884
rect 10652 31872 10658 31884
rect 10781 31875 10839 31881
rect 10781 31872 10793 31875
rect 10652 31844 10793 31872
rect 10652 31832 10658 31844
rect 10781 31841 10793 31844
rect 10827 31841 10839 31875
rect 10781 31835 10839 31841
rect 11054 31832 11060 31884
rect 11112 31872 11118 31884
rect 12529 31875 12587 31881
rect 12529 31872 12541 31875
rect 11112 31844 12541 31872
rect 11112 31832 11118 31844
rect 12529 31841 12541 31844
rect 12575 31872 12587 31875
rect 12986 31872 12992 31884
rect 12575 31844 12992 31872
rect 12575 31841 12587 31844
rect 12529 31835 12587 31841
rect 12986 31832 12992 31844
rect 13044 31832 13050 31884
rect 13354 31832 13360 31884
rect 13412 31872 13418 31884
rect 13412 31844 13768 31872
rect 13412 31832 13418 31844
rect 10045 31807 10103 31813
rect 10045 31804 10057 31807
rect 9640 31776 10057 31804
rect 9640 31764 9646 31776
rect 10045 31773 10057 31776
rect 10091 31773 10103 31807
rect 10045 31767 10103 31773
rect 10134 31764 10140 31816
rect 10192 31804 10198 31816
rect 13630 31804 13636 31816
rect 10192 31776 10237 31804
rect 13591 31776 13636 31804
rect 10192 31764 10198 31776
rect 13630 31764 13636 31776
rect 13688 31764 13694 31816
rect 13740 31813 13768 31844
rect 13725 31807 13783 31813
rect 13725 31773 13737 31807
rect 13771 31773 13783 31807
rect 13832 31804 13860 31912
rect 15304 31912 16028 31940
rect 13998 31832 14004 31884
rect 14056 31872 14062 31884
rect 14369 31875 14427 31881
rect 14369 31872 14381 31875
rect 14056 31844 14381 31872
rect 14056 31832 14062 31844
rect 14369 31841 14381 31844
rect 14415 31841 14427 31875
rect 14369 31835 14427 31841
rect 14642 31832 14648 31884
rect 14700 31872 14706 31884
rect 15304 31872 15332 31912
rect 16022 31900 16028 31912
rect 16080 31900 16086 31952
rect 16390 31940 16396 31952
rect 16351 31912 16396 31940
rect 16390 31900 16396 31912
rect 16448 31900 16454 31952
rect 16942 31900 16948 31952
rect 17000 31940 17006 31952
rect 20162 31940 20168 31952
rect 17000 31912 20168 31940
rect 17000 31900 17006 31912
rect 20162 31900 20168 31912
rect 20220 31900 20226 31952
rect 22830 31940 22836 31952
rect 22791 31912 22836 31940
rect 22830 31900 22836 31912
rect 22888 31900 22894 31952
rect 14700 31844 15332 31872
rect 14700 31832 14706 31844
rect 15378 31832 15384 31884
rect 15436 31872 15442 31884
rect 15746 31872 15752 31884
rect 15436 31844 15481 31872
rect 15707 31844 15752 31872
rect 15436 31832 15442 31844
rect 15746 31832 15752 31844
rect 15804 31832 15810 31884
rect 16574 31832 16580 31884
rect 16632 31872 16638 31884
rect 17586 31872 17592 31884
rect 16632 31844 17592 31872
rect 16632 31832 16638 31844
rect 17586 31832 17592 31844
rect 17644 31832 17650 31884
rect 17954 31832 17960 31884
rect 18012 31872 18018 31884
rect 21177 31875 21235 31881
rect 21177 31872 21189 31875
rect 18012 31844 21189 31872
rect 18012 31832 18018 31844
rect 21177 31841 21189 31844
rect 21223 31841 21235 31875
rect 22186 31872 22192 31884
rect 21177 31835 21235 31841
rect 21284 31844 22192 31872
rect 14277 31807 14335 31813
rect 14277 31804 14289 31807
rect 13832 31776 14289 31804
rect 13725 31767 13783 31773
rect 14277 31773 14289 31776
rect 14323 31773 14335 31807
rect 18782 31804 18788 31816
rect 18743 31776 18788 31804
rect 14277 31767 14335 31773
rect 18782 31764 18788 31776
rect 18840 31764 18846 31816
rect 18877 31807 18935 31813
rect 18877 31773 18889 31807
rect 18923 31804 18935 31807
rect 19426 31804 19432 31816
rect 18923 31776 19432 31804
rect 18923 31773 18935 31776
rect 18877 31767 18935 31773
rect 19426 31764 19432 31776
rect 19484 31764 19490 31816
rect 19613 31807 19671 31813
rect 19613 31773 19625 31807
rect 19659 31804 19671 31807
rect 19659 31776 19693 31804
rect 19659 31773 19671 31776
rect 19613 31767 19671 31773
rect 9490 31736 9496 31748
rect 8404 31708 9496 31736
rect 4157 31671 4215 31677
rect 4157 31637 4169 31671
rect 4203 31668 4215 31671
rect 4246 31668 4252 31680
rect 4203 31640 4252 31668
rect 4203 31637 4215 31640
rect 4157 31631 4215 31637
rect 4246 31628 4252 31640
rect 4304 31628 4310 31680
rect 6086 31628 6092 31680
rect 6144 31668 6150 31680
rect 8404 31668 8432 31708
rect 9490 31696 9496 31708
rect 9548 31696 9554 31748
rect 11822 31708 12204 31736
rect 6144 31640 8432 31668
rect 6144 31628 6150 31640
rect 8570 31628 8576 31680
rect 8628 31668 8634 31680
rect 11330 31668 11336 31680
rect 8628 31640 11336 31668
rect 8628 31628 8634 31640
rect 11330 31628 11336 31640
rect 11388 31628 11394 31680
rect 12176 31668 12204 31708
rect 12250 31696 12256 31748
rect 12308 31736 12314 31748
rect 13906 31736 13912 31748
rect 12308 31708 12353 31736
rect 12406 31708 13912 31736
rect 12308 31696 12314 31708
rect 12406 31668 12434 31708
rect 13906 31696 13912 31708
rect 13964 31696 13970 31748
rect 15654 31736 15660 31748
rect 15615 31708 15660 31736
rect 15654 31696 15660 31708
rect 15712 31696 15718 31748
rect 16758 31696 16764 31748
rect 16816 31736 16822 31748
rect 16853 31739 16911 31745
rect 16853 31736 16865 31739
rect 16816 31708 16865 31736
rect 16816 31696 16822 31708
rect 16853 31705 16865 31708
rect 16899 31705 16911 31739
rect 16853 31699 16911 31705
rect 16945 31739 17003 31745
rect 16945 31705 16957 31739
rect 16991 31705 17003 31739
rect 17586 31736 17592 31748
rect 17547 31708 17592 31736
rect 16945 31699 17003 31705
rect 12176 31640 12434 31668
rect 12526 31628 12532 31680
rect 12584 31668 12590 31680
rect 14182 31668 14188 31680
rect 12584 31640 14188 31668
rect 12584 31628 12590 31640
rect 14182 31628 14188 31640
rect 14240 31628 14246 31680
rect 16574 31628 16580 31680
rect 16632 31668 16638 31680
rect 16960 31668 16988 31699
rect 17586 31696 17592 31708
rect 17644 31696 17650 31748
rect 17678 31696 17684 31748
rect 17736 31736 17742 31748
rect 18230 31736 18236 31748
rect 17736 31708 17781 31736
rect 18191 31708 18236 31736
rect 17736 31696 17742 31708
rect 18230 31696 18236 31708
rect 18288 31696 18294 31748
rect 19334 31696 19340 31748
rect 19392 31736 19398 31748
rect 19628 31736 19656 31767
rect 20070 31764 20076 31816
rect 20128 31804 20134 31816
rect 20257 31807 20315 31813
rect 20128 31776 20208 31804
rect 20128 31764 20134 31776
rect 19978 31736 19984 31748
rect 19392 31708 19984 31736
rect 19392 31696 19398 31708
rect 19978 31696 19984 31708
rect 20036 31696 20042 31748
rect 20180 31745 20208 31776
rect 20257 31773 20269 31807
rect 20303 31804 20315 31807
rect 20714 31804 20720 31816
rect 20303 31776 20720 31804
rect 20303 31773 20315 31776
rect 20257 31767 20315 31773
rect 20714 31764 20720 31776
rect 20772 31764 20778 31816
rect 21284 31813 21312 31844
rect 22186 31832 22192 31844
rect 22244 31832 22250 31884
rect 21269 31807 21327 31813
rect 21269 31773 21281 31807
rect 21315 31773 21327 31807
rect 21269 31767 21327 31773
rect 20165 31739 20223 31745
rect 20165 31705 20177 31739
rect 20211 31736 20223 31739
rect 20211 31708 20245 31736
rect 20211 31705 20223 31708
rect 20165 31699 20223 31705
rect 16632 31640 16988 31668
rect 16632 31628 16638 31640
rect 17494 31628 17500 31680
rect 17552 31668 17558 31680
rect 20898 31668 20904 31680
rect 17552 31640 20904 31668
rect 17552 31628 17558 31640
rect 20898 31628 20904 31640
rect 20956 31628 20962 31680
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 5905 31467 5963 31473
rect 5905 31433 5917 31467
rect 5951 31464 5963 31467
rect 8294 31464 8300 31476
rect 5951 31436 8300 31464
rect 5951 31433 5963 31436
rect 5905 31427 5963 31433
rect 8294 31424 8300 31436
rect 8352 31424 8358 31476
rect 10686 31424 10692 31476
rect 10744 31464 10750 31476
rect 19150 31464 19156 31476
rect 10744 31436 14872 31464
rect 10744 31424 10750 31436
rect 3142 31356 3148 31408
rect 3200 31396 3206 31408
rect 3237 31399 3295 31405
rect 3237 31396 3249 31399
rect 3200 31368 3249 31396
rect 3200 31356 3206 31368
rect 3237 31365 3249 31368
rect 3283 31365 3295 31399
rect 3237 31359 3295 31365
rect 4246 31356 4252 31408
rect 4304 31356 4310 31408
rect 8478 31356 8484 31408
rect 8536 31356 8542 31408
rect 8846 31356 8852 31408
rect 8904 31396 8910 31408
rect 11698 31396 11704 31408
rect 8904 31368 11704 31396
rect 8904 31356 8910 31368
rect 1670 31328 1676 31340
rect 1583 31300 1676 31328
rect 1670 31288 1676 31300
rect 1728 31328 1734 31340
rect 2222 31328 2228 31340
rect 1728 31300 2228 31328
rect 1728 31288 1734 31300
rect 2222 31288 2228 31300
rect 2280 31288 2286 31340
rect 2501 31331 2559 31337
rect 2501 31297 2513 31331
rect 2547 31328 2559 31331
rect 2590 31328 2596 31340
rect 2547 31300 2596 31328
rect 2547 31297 2559 31300
rect 2501 31291 2559 31297
rect 2590 31288 2596 31300
rect 2648 31288 2654 31340
rect 5442 31288 5448 31340
rect 5500 31328 5506 31340
rect 5813 31331 5871 31337
rect 5813 31328 5825 31331
rect 5500 31300 5825 31328
rect 5500 31288 5506 31300
rect 5813 31297 5825 31300
rect 5859 31328 5871 31331
rect 6733 31331 6791 31337
rect 6733 31328 6745 31331
rect 5859 31300 6745 31328
rect 5859 31297 5871 31300
rect 5813 31291 5871 31297
rect 6733 31297 6745 31300
rect 6779 31328 6791 31331
rect 7466 31328 7472 31340
rect 6779 31300 7472 31328
rect 6779 31297 6791 31300
rect 6733 31291 6791 31297
rect 7466 31288 7472 31300
rect 7524 31288 7530 31340
rect 9398 31288 9404 31340
rect 9456 31328 9462 31340
rect 10336 31337 10364 31368
rect 11698 31356 11704 31368
rect 11756 31356 11762 31408
rect 12710 31356 12716 31408
rect 12768 31356 12774 31408
rect 13170 31356 13176 31408
rect 13228 31396 13234 31408
rect 14844 31396 14872 31436
rect 18248 31436 19156 31464
rect 18248 31408 18276 31436
rect 15013 31399 15071 31405
rect 15013 31396 15025 31399
rect 13228 31368 14228 31396
rect 14844 31368 15025 31396
rect 13228 31356 13234 31368
rect 10321 31331 10379 31337
rect 9456 31300 9501 31328
rect 9456 31288 9462 31300
rect 10321 31297 10333 31331
rect 10367 31297 10379 31331
rect 10321 31291 10379 31297
rect 10870 31288 10876 31340
rect 10928 31328 10934 31340
rect 14200 31337 14228 31368
rect 15013 31365 15025 31368
rect 15059 31365 15071 31399
rect 17310 31396 17316 31408
rect 17271 31368 17316 31396
rect 15013 31359 15071 31365
rect 17310 31356 17316 31368
rect 17368 31356 17374 31408
rect 17865 31399 17923 31405
rect 17865 31365 17877 31399
rect 17911 31396 17923 31399
rect 18230 31396 18236 31408
rect 17911 31368 18236 31396
rect 17911 31365 17923 31368
rect 17865 31359 17923 31365
rect 18230 31356 18236 31368
rect 18288 31356 18294 31408
rect 18506 31396 18512 31408
rect 18467 31368 18512 31396
rect 18506 31356 18512 31368
rect 18564 31356 18570 31408
rect 19076 31405 19104 31436
rect 19150 31424 19156 31436
rect 19208 31424 19214 31476
rect 19242 31424 19248 31476
rect 19300 31464 19306 31476
rect 20346 31464 20352 31476
rect 19300 31436 20352 31464
rect 19300 31424 19306 31436
rect 20346 31424 20352 31436
rect 20404 31424 20410 31476
rect 20898 31464 20904 31476
rect 20859 31436 20904 31464
rect 20898 31424 20904 31436
rect 20956 31424 20962 31476
rect 22094 31464 22100 31476
rect 22055 31436 22100 31464
rect 22094 31424 22100 31436
rect 22152 31464 22158 31476
rect 22554 31464 22560 31476
rect 22152 31436 22560 31464
rect 22152 31424 22158 31436
rect 22554 31424 22560 31436
rect 22612 31424 22618 31476
rect 23201 31467 23259 31473
rect 23201 31433 23213 31467
rect 23247 31464 23259 31467
rect 23658 31464 23664 31476
rect 23247 31436 23664 31464
rect 23247 31433 23259 31436
rect 23201 31427 23259 31433
rect 23658 31424 23664 31436
rect 23716 31424 23722 31476
rect 19061 31399 19119 31405
rect 19061 31365 19073 31399
rect 19107 31365 19119 31399
rect 19061 31359 19119 31365
rect 19334 31356 19340 31408
rect 19392 31396 19398 31408
rect 20254 31396 20260 31408
rect 19392 31368 20260 31396
rect 19392 31356 19398 31368
rect 20254 31356 20260 31368
rect 20312 31356 20318 31408
rect 10965 31331 11023 31337
rect 10965 31328 10977 31331
rect 10928 31300 10977 31328
rect 10928 31288 10934 31300
rect 10965 31297 10977 31300
rect 11011 31297 11023 31331
rect 10965 31291 11023 31297
rect 14185 31331 14243 31337
rect 14185 31297 14197 31331
rect 14231 31328 14243 31331
rect 14274 31328 14280 31340
rect 14231 31300 14280 31328
rect 14231 31297 14243 31300
rect 14185 31291 14243 31297
rect 14274 31288 14280 31300
rect 14332 31288 14338 31340
rect 16022 31328 16028 31340
rect 15983 31300 16028 31328
rect 16022 31288 16028 31300
rect 16080 31288 16086 31340
rect 19426 31288 19432 31340
rect 19484 31328 19490 31340
rect 19705 31331 19763 31337
rect 19705 31328 19717 31331
rect 19484 31300 19717 31328
rect 19484 31288 19490 31300
rect 19705 31297 19717 31300
rect 19751 31297 19763 31331
rect 19705 31291 19763 31297
rect 19978 31288 19984 31340
rect 20036 31328 20042 31340
rect 20349 31331 20407 31337
rect 20349 31328 20361 31331
rect 20036 31300 20361 31328
rect 20036 31288 20042 31300
rect 20349 31297 20361 31300
rect 20395 31328 20407 31331
rect 20809 31331 20867 31337
rect 20809 31328 20821 31331
rect 20395 31300 20821 31328
rect 20395 31297 20407 31300
rect 20349 31291 20407 31297
rect 20809 31297 20821 31300
rect 20855 31297 20867 31331
rect 20809 31291 20867 31297
rect 2961 31263 3019 31269
rect 2961 31229 2973 31263
rect 3007 31260 3019 31263
rect 3970 31260 3976 31272
rect 3007 31232 3976 31260
rect 3007 31229 3019 31232
rect 2961 31223 3019 31229
rect 3970 31220 3976 31232
rect 4028 31220 4034 31272
rect 4985 31263 5043 31269
rect 4985 31229 4997 31263
rect 5031 31229 5043 31263
rect 4985 31223 5043 31229
rect 1854 31192 1860 31204
rect 1815 31164 1860 31192
rect 1854 31152 1860 31164
rect 1912 31152 1918 31204
rect 5000 31192 5028 31223
rect 5994 31220 6000 31272
rect 6052 31260 6058 31272
rect 7377 31263 7435 31269
rect 7377 31260 7389 31263
rect 6052 31232 7389 31260
rect 6052 31220 6058 31232
rect 7377 31229 7389 31232
rect 7423 31229 7435 31263
rect 9122 31260 9128 31272
rect 9083 31232 9128 31260
rect 7377 31223 7435 31229
rect 9122 31220 9128 31232
rect 9180 31220 9186 31272
rect 11330 31220 11336 31272
rect 11388 31260 11394 31272
rect 11698 31260 11704 31272
rect 11388 31232 11704 31260
rect 11388 31220 11394 31232
rect 11698 31220 11704 31232
rect 11756 31260 11762 31272
rect 13170 31260 13176 31272
rect 11756 31232 13176 31260
rect 11756 31220 11762 31232
rect 13170 31220 13176 31232
rect 13228 31220 13234 31272
rect 13262 31220 13268 31272
rect 13320 31260 13326 31272
rect 13541 31263 13599 31269
rect 13541 31260 13553 31263
rect 13320 31232 13365 31260
rect 13464 31232 13553 31260
rect 13320 31220 13326 31232
rect 7742 31192 7748 31204
rect 5000 31164 7748 31192
rect 7742 31152 7748 31164
rect 7800 31152 7806 31204
rect 10962 31192 10968 31204
rect 9646 31164 10968 31192
rect 2314 31124 2320 31136
rect 2275 31096 2320 31124
rect 2314 31084 2320 31096
rect 2372 31084 2378 31136
rect 5166 31084 5172 31136
rect 5224 31124 5230 31136
rect 5442 31124 5448 31136
rect 5224 31096 5448 31124
rect 5224 31084 5230 31096
rect 5442 31084 5448 31096
rect 5500 31084 5506 31136
rect 6825 31127 6883 31133
rect 6825 31093 6837 31127
rect 6871 31124 6883 31127
rect 9646 31124 9674 31164
rect 10962 31152 10968 31164
rect 11020 31152 11026 31204
rect 10410 31124 10416 31136
rect 6871 31096 9674 31124
rect 10371 31096 10416 31124
rect 6871 31093 6883 31096
rect 6825 31087 6883 31093
rect 10410 31084 10416 31096
rect 10468 31084 10474 31136
rect 11057 31127 11115 31133
rect 11057 31093 11069 31127
rect 11103 31124 11115 31127
rect 11606 31124 11612 31136
rect 11103 31096 11612 31124
rect 11103 31093 11115 31096
rect 11057 31087 11115 31093
rect 11606 31084 11612 31096
rect 11664 31084 11670 31136
rect 11793 31127 11851 31133
rect 11793 31093 11805 31127
rect 11839 31124 11851 31127
rect 12802 31124 12808 31136
rect 11839 31096 12808 31124
rect 11839 31093 11851 31096
rect 11793 31087 11851 31093
rect 12802 31084 12808 31096
rect 12860 31084 12866 31136
rect 13078 31084 13084 31136
rect 13136 31124 13142 31136
rect 13464 31124 13492 31232
rect 13541 31229 13553 31232
rect 13587 31229 13599 31263
rect 13541 31223 13599 31229
rect 14921 31263 14979 31269
rect 14921 31229 14933 31263
rect 14967 31260 14979 31263
rect 15010 31260 15016 31272
rect 14967 31232 15016 31260
rect 14967 31229 14979 31232
rect 14921 31223 14979 31229
rect 15010 31220 15016 31232
rect 15068 31220 15074 31272
rect 15194 31260 15200 31272
rect 15155 31232 15200 31260
rect 15194 31220 15200 31232
rect 15252 31260 15258 31272
rect 15838 31260 15844 31272
rect 15252 31232 15844 31260
rect 15252 31220 15258 31232
rect 15838 31220 15844 31232
rect 15896 31220 15902 31272
rect 17218 31260 17224 31272
rect 17179 31232 17224 31260
rect 17218 31220 17224 31232
rect 17276 31220 17282 31272
rect 18417 31263 18475 31269
rect 18417 31229 18429 31263
rect 18463 31260 18475 31263
rect 20438 31260 20444 31272
rect 18463 31232 20444 31260
rect 18463 31229 18475 31232
rect 18417 31223 18475 31229
rect 20438 31220 20444 31232
rect 20496 31220 20502 31272
rect 13906 31152 13912 31204
rect 13964 31192 13970 31204
rect 20257 31195 20315 31201
rect 20257 31192 20269 31195
rect 13964 31164 20269 31192
rect 13964 31152 13970 31164
rect 20257 31161 20269 31164
rect 20303 31161 20315 31195
rect 20257 31155 20315 31161
rect 13136 31096 13492 31124
rect 14277 31127 14335 31133
rect 13136 31084 13142 31096
rect 14277 31093 14289 31127
rect 14323 31124 14335 31127
rect 15286 31124 15292 31136
rect 14323 31096 15292 31124
rect 14323 31093 14335 31096
rect 14277 31087 14335 31093
rect 15286 31084 15292 31096
rect 15344 31084 15350 31136
rect 15378 31084 15384 31136
rect 15436 31124 15442 31136
rect 16117 31127 16175 31133
rect 16117 31124 16129 31127
rect 15436 31096 16129 31124
rect 15436 31084 15442 31096
rect 16117 31093 16129 31096
rect 16163 31093 16175 31127
rect 16117 31087 16175 31093
rect 16206 31084 16212 31136
rect 16264 31124 16270 31136
rect 18138 31124 18144 31136
rect 16264 31096 18144 31124
rect 16264 31084 16270 31096
rect 18138 31084 18144 31096
rect 18196 31084 18202 31136
rect 19426 31084 19432 31136
rect 19484 31124 19490 31136
rect 19613 31127 19671 31133
rect 19613 31124 19625 31127
rect 19484 31096 19625 31124
rect 19484 31084 19490 31096
rect 19613 31093 19625 31096
rect 19659 31093 19671 31127
rect 19613 31087 19671 31093
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 4798 30880 4804 30932
rect 4856 30920 4862 30932
rect 5258 30920 5264 30932
rect 4856 30892 5264 30920
rect 4856 30880 4862 30892
rect 5258 30880 5264 30892
rect 5316 30880 5322 30932
rect 7650 30880 7656 30932
rect 7708 30920 7714 30932
rect 9217 30923 9275 30929
rect 7708 30892 9168 30920
rect 7708 30880 7714 30892
rect 8754 30852 8760 30864
rect 8496 30824 8760 30852
rect 4249 30787 4307 30793
rect 4249 30753 4261 30787
rect 4295 30784 4307 30787
rect 4706 30784 4712 30796
rect 4295 30756 4712 30784
rect 4295 30753 4307 30756
rect 4249 30747 4307 30753
rect 4706 30744 4712 30756
rect 4764 30784 4770 30796
rect 4890 30784 4896 30796
rect 4764 30756 4896 30784
rect 4764 30744 4770 30756
rect 4890 30744 4896 30756
rect 4948 30744 4954 30796
rect 5626 30744 5632 30796
rect 5684 30784 5690 30796
rect 8496 30784 8524 30824
rect 8754 30812 8760 30824
rect 8812 30812 8818 30864
rect 9140 30852 9168 30892
rect 9217 30889 9229 30923
rect 9263 30920 9275 30923
rect 9398 30920 9404 30932
rect 9263 30892 9404 30920
rect 9263 30889 9275 30892
rect 9217 30883 9275 30889
rect 9398 30880 9404 30892
rect 9456 30880 9462 30932
rect 10413 30923 10471 30929
rect 10413 30889 10425 30923
rect 10459 30920 10471 30923
rect 11054 30920 11060 30932
rect 10459 30892 11060 30920
rect 10459 30889 10471 30892
rect 10413 30883 10471 30889
rect 11054 30880 11060 30892
rect 11112 30880 11118 30932
rect 11238 30880 11244 30932
rect 11296 30920 11302 30932
rect 12342 30920 12348 30932
rect 11296 30892 12348 30920
rect 11296 30880 11302 30892
rect 12342 30880 12348 30892
rect 12400 30880 12406 30932
rect 12710 30880 12716 30932
rect 12768 30920 12774 30932
rect 20162 30920 20168 30932
rect 12768 30892 19656 30920
rect 20123 30892 20168 30920
rect 12768 30880 12774 30892
rect 9140 30824 9812 30852
rect 5684 30756 8524 30784
rect 8573 30787 8631 30793
rect 5684 30744 5690 30756
rect 8573 30753 8585 30787
rect 8619 30784 8631 30787
rect 9398 30784 9404 30796
rect 8619 30756 9404 30784
rect 8619 30753 8631 30756
rect 8573 30747 8631 30753
rect 9398 30744 9404 30756
rect 9456 30744 9462 30796
rect 9784 30784 9812 30824
rect 9858 30812 9864 30864
rect 9916 30852 9922 30864
rect 10502 30852 10508 30864
rect 9916 30824 10508 30852
rect 9916 30812 9922 30824
rect 10502 30812 10508 30824
rect 10560 30852 10566 30864
rect 10870 30852 10876 30864
rect 10560 30824 10876 30852
rect 10560 30812 10566 30824
rect 10870 30812 10876 30824
rect 10928 30812 10934 30864
rect 16206 30852 16212 30864
rect 16167 30824 16212 30852
rect 16206 30812 16212 30824
rect 16264 30812 16270 30864
rect 17954 30812 17960 30864
rect 18012 30852 18018 30864
rect 19521 30855 19579 30861
rect 19521 30852 19533 30855
rect 18012 30824 19533 30852
rect 18012 30812 18018 30824
rect 19521 30821 19533 30824
rect 19567 30821 19579 30855
rect 19628 30852 19656 30892
rect 20162 30880 20168 30892
rect 20220 30880 20226 30932
rect 20714 30920 20720 30932
rect 20675 30892 20720 30920
rect 20714 30880 20720 30892
rect 20772 30880 20778 30932
rect 21729 30855 21787 30861
rect 21729 30852 21741 30855
rect 19628 30824 21741 30852
rect 19521 30815 19579 30821
rect 21729 30821 21741 30824
rect 21775 30821 21787 30855
rect 21729 30815 21787 30821
rect 31113 30855 31171 30861
rect 31113 30821 31125 30855
rect 31159 30852 31171 30855
rect 37274 30852 37280 30864
rect 31159 30824 37280 30852
rect 31159 30821 31171 30824
rect 31113 30815 31171 30821
rect 37274 30812 37280 30824
rect 37332 30812 37338 30864
rect 9784 30756 10364 30784
rect 3418 30676 3424 30728
rect 3476 30716 3482 30728
rect 3970 30716 3976 30728
rect 3476 30688 3976 30716
rect 3476 30676 3482 30688
rect 3970 30676 3976 30688
rect 4028 30676 4034 30728
rect 5902 30676 5908 30728
rect 5960 30716 5966 30728
rect 5997 30719 6055 30725
rect 5997 30716 6009 30719
rect 5960 30688 6009 30716
rect 5960 30676 5966 30688
rect 5997 30685 6009 30688
rect 6043 30716 6055 30719
rect 6178 30716 6184 30728
rect 6043 30688 6184 30716
rect 6043 30685 6055 30688
rect 5997 30679 6055 30685
rect 6178 30676 6184 30688
rect 6236 30676 6242 30728
rect 9677 30719 9735 30725
rect 9677 30685 9689 30719
rect 9723 30716 9735 30719
rect 9950 30716 9956 30728
rect 9723 30688 9956 30716
rect 9723 30685 9735 30688
rect 9677 30679 9735 30685
rect 9950 30676 9956 30688
rect 10008 30676 10014 30728
rect 10336 30725 10364 30756
rect 10410 30744 10416 30796
rect 10468 30784 10474 30796
rect 15010 30784 15016 30796
rect 10468 30756 13676 30784
rect 14971 30756 15016 30784
rect 10468 30744 10474 30756
rect 10321 30719 10379 30725
rect 10321 30685 10333 30719
rect 10367 30685 10379 30719
rect 10321 30679 10379 30685
rect 10965 30719 11023 30725
rect 10965 30685 10977 30719
rect 11011 30716 11023 30719
rect 11238 30716 11244 30728
rect 11011 30688 11244 30716
rect 11011 30685 11023 30688
rect 10965 30679 11023 30685
rect 11238 30676 11244 30688
rect 11296 30676 11302 30728
rect 12986 30676 12992 30728
rect 13044 30716 13050 30728
rect 13044 30688 13089 30716
rect 13044 30676 13050 30688
rect 13170 30676 13176 30728
rect 13228 30716 13234 30728
rect 13541 30719 13599 30725
rect 13541 30716 13553 30719
rect 13228 30688 13553 30716
rect 13228 30676 13234 30688
rect 13541 30685 13553 30688
rect 13587 30685 13599 30719
rect 13541 30679 13599 30685
rect 2498 30608 2504 30660
rect 2556 30608 2562 30660
rect 3145 30651 3203 30657
rect 3145 30617 3157 30651
rect 3191 30648 3203 30651
rect 3191 30620 4660 30648
rect 3191 30617 3203 30620
rect 3145 30611 3203 30617
rect 1673 30583 1731 30589
rect 1673 30549 1685 30583
rect 1719 30580 1731 30583
rect 1762 30580 1768 30592
rect 1719 30552 1768 30580
rect 1719 30549 1731 30552
rect 1673 30543 1731 30549
rect 1762 30540 1768 30552
rect 1820 30580 1826 30592
rect 3234 30580 3240 30592
rect 1820 30552 3240 30580
rect 1820 30540 1826 30552
rect 3234 30540 3240 30552
rect 3292 30540 3298 30592
rect 4632 30580 4660 30620
rect 5258 30608 5264 30660
rect 5316 30608 5322 30660
rect 6549 30651 6607 30657
rect 6549 30617 6561 30651
rect 6595 30617 6607 30651
rect 6549 30611 6607 30617
rect 5626 30580 5632 30592
rect 4632 30552 5632 30580
rect 5626 30540 5632 30552
rect 5684 30540 5690 30592
rect 6564 30580 6592 30611
rect 6914 30608 6920 30660
rect 6972 30648 6978 30660
rect 8297 30651 8355 30657
rect 6972 30620 7130 30648
rect 6972 30608 6978 30620
rect 8297 30617 8309 30651
rect 8343 30648 8355 30651
rect 8570 30648 8576 30660
rect 8343 30620 8576 30648
rect 8343 30617 8355 30620
rect 8297 30611 8355 30617
rect 8570 30608 8576 30620
rect 8628 30648 8634 30660
rect 9582 30648 9588 30660
rect 8628 30620 9588 30648
rect 8628 30608 8634 30620
rect 9582 30608 9588 30620
rect 9640 30608 9646 30660
rect 9769 30651 9827 30657
rect 9769 30617 9781 30651
rect 9815 30648 9827 30651
rect 9815 30620 10916 30648
rect 9815 30617 9827 30620
rect 9769 30611 9827 30617
rect 8846 30580 8852 30592
rect 6564 30552 8852 30580
rect 8846 30540 8852 30552
rect 8904 30540 8910 30592
rect 10888 30580 10916 30620
rect 12250 30608 12256 30660
rect 12308 30608 12314 30660
rect 12713 30651 12771 30657
rect 12713 30617 12725 30651
rect 12759 30648 12771 30651
rect 12802 30648 12808 30660
rect 12759 30620 12808 30648
rect 12759 30617 12771 30620
rect 12713 30611 12771 30617
rect 12802 30608 12808 30620
rect 12860 30648 12866 30660
rect 13262 30648 13268 30660
rect 12860 30620 13268 30648
rect 12860 30608 12866 30620
rect 13262 30608 13268 30620
rect 13320 30608 13326 30660
rect 13648 30648 13676 30756
rect 15010 30744 15016 30756
rect 15068 30744 15074 30796
rect 16298 30744 16304 30796
rect 16356 30784 16362 30796
rect 16356 30756 19472 30784
rect 16356 30744 16362 30756
rect 14274 30716 14280 30728
rect 14235 30688 14280 30716
rect 14274 30676 14280 30688
rect 14332 30676 14338 30728
rect 18414 30676 18420 30728
rect 18472 30716 18478 30728
rect 19444 30725 19472 30756
rect 20346 30744 20352 30796
rect 20404 30784 20410 30796
rect 20404 30756 30972 30784
rect 20404 30744 20410 30756
rect 18601 30719 18659 30725
rect 18601 30716 18613 30719
rect 18472 30688 18613 30716
rect 18472 30676 18478 30688
rect 18601 30685 18613 30688
rect 18647 30685 18659 30719
rect 18601 30679 18659 30685
rect 19429 30719 19487 30725
rect 19429 30685 19441 30719
rect 19475 30685 19487 30719
rect 20254 30716 20260 30728
rect 20215 30688 20260 30716
rect 19429 30679 19487 30685
rect 20254 30676 20260 30688
rect 20312 30676 20318 30728
rect 21821 30719 21879 30725
rect 21821 30685 21833 30719
rect 21867 30716 21879 30719
rect 22186 30716 22192 30728
rect 21867 30688 22192 30716
rect 21867 30685 21879 30688
rect 21821 30679 21879 30685
rect 22186 30676 22192 30688
rect 22244 30716 22250 30728
rect 30944 30725 30972 30756
rect 22465 30719 22523 30725
rect 22465 30716 22477 30719
rect 22244 30688 22477 30716
rect 22244 30676 22250 30688
rect 22465 30685 22477 30688
rect 22511 30685 22523 30719
rect 22465 30679 22523 30685
rect 30929 30719 30987 30725
rect 30929 30685 30941 30719
rect 30975 30716 30987 30719
rect 31573 30719 31631 30725
rect 31573 30716 31585 30719
rect 30975 30688 31585 30716
rect 30975 30685 30987 30688
rect 30929 30679 30987 30685
rect 31573 30685 31585 30688
rect 31619 30685 31631 30719
rect 31573 30679 31631 30685
rect 15105 30651 15163 30657
rect 15105 30648 15117 30651
rect 13648 30620 15117 30648
rect 15105 30617 15117 30620
rect 15151 30617 15163 30651
rect 15105 30611 15163 30617
rect 15657 30651 15715 30657
rect 15657 30617 15669 30651
rect 15703 30648 15715 30651
rect 15838 30648 15844 30660
rect 15703 30620 15844 30648
rect 15703 30617 15715 30620
rect 15657 30611 15715 30617
rect 15838 30608 15844 30620
rect 15896 30608 15902 30660
rect 16669 30651 16727 30657
rect 16669 30617 16681 30651
rect 16715 30617 16727 30651
rect 16669 30611 16727 30617
rect 13078 30580 13084 30592
rect 10888 30552 13084 30580
rect 13078 30540 13084 30552
rect 13136 30540 13142 30592
rect 13633 30583 13691 30589
rect 13633 30549 13645 30583
rect 13679 30580 13691 30583
rect 14182 30580 14188 30592
rect 13679 30552 14188 30580
rect 13679 30549 13691 30552
rect 13633 30543 13691 30549
rect 14182 30540 14188 30552
rect 14240 30540 14246 30592
rect 14274 30540 14280 30592
rect 14332 30580 14338 30592
rect 14369 30583 14427 30589
rect 14369 30580 14381 30583
rect 14332 30552 14381 30580
rect 14332 30540 14338 30552
rect 14369 30549 14381 30552
rect 14415 30549 14427 30583
rect 14369 30543 14427 30549
rect 15010 30540 15016 30592
rect 15068 30580 15074 30592
rect 16114 30580 16120 30592
rect 15068 30552 16120 30580
rect 15068 30540 15074 30552
rect 16114 30540 16120 30552
rect 16172 30540 16178 30592
rect 16684 30580 16712 30611
rect 16758 30608 16764 30660
rect 16816 30648 16822 30660
rect 17313 30651 17371 30657
rect 16816 30620 16861 30648
rect 16816 30608 16822 30620
rect 17313 30617 17325 30651
rect 17359 30648 17371 30651
rect 17586 30648 17592 30660
rect 17359 30620 17592 30648
rect 17359 30617 17371 30620
rect 17313 30611 17371 30617
rect 17586 30608 17592 30620
rect 17644 30608 17650 30660
rect 17862 30648 17868 30660
rect 17823 30620 17868 30648
rect 17862 30608 17868 30620
rect 17920 30608 17926 30660
rect 17957 30651 18015 30657
rect 17957 30617 17969 30651
rect 18003 30648 18015 30651
rect 18509 30651 18567 30657
rect 18509 30648 18521 30651
rect 18003 30620 18521 30648
rect 18003 30617 18015 30620
rect 17957 30611 18015 30617
rect 18509 30617 18521 30620
rect 18555 30617 18567 30651
rect 20806 30648 20812 30660
rect 18509 30611 18567 30617
rect 19444 30620 20812 30648
rect 19444 30580 19472 30620
rect 20806 30608 20812 30620
rect 20864 30608 20870 30660
rect 16684 30552 19472 30580
rect 21818 30540 21824 30592
rect 21876 30580 21882 30592
rect 22373 30583 22431 30589
rect 22373 30580 22385 30583
rect 21876 30552 22385 30580
rect 21876 30540 21882 30552
rect 22373 30549 22385 30552
rect 22419 30549 22431 30583
rect 22373 30543 22431 30549
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 7282 30336 7288 30388
rect 7340 30376 7346 30388
rect 7650 30376 7656 30388
rect 7340 30348 7656 30376
rect 7340 30336 7346 30348
rect 7650 30336 7656 30348
rect 7708 30336 7714 30388
rect 9122 30336 9128 30388
rect 9180 30376 9186 30388
rect 9401 30379 9459 30385
rect 9401 30376 9413 30379
rect 9180 30348 9413 30376
rect 9180 30336 9186 30348
rect 9401 30345 9413 30348
rect 9447 30376 9459 30379
rect 9447 30348 10548 30376
rect 9447 30345 9459 30348
rect 9401 30339 9459 30345
rect 3145 30311 3203 30317
rect 3145 30277 3157 30311
rect 3191 30308 3203 30311
rect 3694 30308 3700 30320
rect 3191 30280 3700 30308
rect 3191 30277 3203 30280
rect 3145 30271 3203 30277
rect 3694 30268 3700 30280
rect 3752 30268 3758 30320
rect 5258 30308 5264 30320
rect 4922 30280 5264 30308
rect 5258 30268 5264 30280
rect 5316 30268 5322 30320
rect 5353 30311 5411 30317
rect 5353 30277 5365 30311
rect 5399 30308 5411 30311
rect 5994 30308 6000 30320
rect 5399 30280 6000 30308
rect 5399 30277 5411 30280
rect 5353 30271 5411 30277
rect 5994 30268 6000 30280
rect 6052 30268 6058 30320
rect 8294 30268 8300 30320
rect 8352 30268 8358 30320
rect 9214 30268 9220 30320
rect 9272 30308 9278 30320
rect 10520 30308 10548 30348
rect 12250 30336 12256 30388
rect 12308 30376 12314 30388
rect 21818 30376 21824 30388
rect 12308 30348 21824 30376
rect 12308 30336 12314 30348
rect 21818 30336 21824 30348
rect 21876 30336 21882 30388
rect 11330 30308 11336 30320
rect 9272 30280 9706 30308
rect 10520 30280 11336 30308
rect 9272 30268 9278 30280
rect 11330 30268 11336 30280
rect 11388 30268 11394 30320
rect 12710 30268 12716 30320
rect 12768 30268 12774 30320
rect 14918 30268 14924 30320
rect 14976 30308 14982 30320
rect 14976 30280 15021 30308
rect 14976 30268 14982 30280
rect 15286 30268 15292 30320
rect 15344 30308 15350 30320
rect 16117 30311 16175 30317
rect 16117 30308 16129 30311
rect 15344 30280 16129 30308
rect 15344 30268 15350 30280
rect 16117 30277 16129 30280
rect 16163 30277 16175 30311
rect 17034 30308 17040 30320
rect 16995 30280 17040 30308
rect 16117 30271 16175 30277
rect 17034 30268 17040 30280
rect 17092 30268 17098 30320
rect 20346 30308 20352 30320
rect 18064 30280 20352 30308
rect 2038 30200 2044 30252
rect 2096 30200 2102 30252
rect 3786 30200 3792 30252
rect 3844 30240 3850 30252
rect 4062 30240 4068 30252
rect 3844 30212 4068 30240
rect 3844 30200 3850 30212
rect 4062 30200 4068 30212
rect 4120 30200 4126 30252
rect 18064 30249 18092 30280
rect 20346 30268 20352 30280
rect 20404 30268 20410 30320
rect 18049 30243 18107 30249
rect 18049 30240 18061 30243
rect 17788 30212 18061 30240
rect 3418 30172 3424 30184
rect 3331 30144 3424 30172
rect 3418 30132 3424 30144
rect 3476 30172 3482 30184
rect 3970 30172 3976 30184
rect 3476 30144 3976 30172
rect 3476 30132 3482 30144
rect 3970 30132 3976 30144
rect 4028 30172 4034 30184
rect 5629 30175 5687 30181
rect 5629 30172 5641 30175
rect 4028 30144 5641 30172
rect 4028 30132 4034 30144
rect 5629 30141 5641 30144
rect 5675 30172 5687 30175
rect 5902 30172 5908 30184
rect 5675 30144 5908 30172
rect 5675 30141 5687 30144
rect 5629 30135 5687 30141
rect 5902 30132 5908 30144
rect 5960 30172 5966 30184
rect 7009 30175 7067 30181
rect 7009 30172 7021 30175
rect 5960 30144 7021 30172
rect 5960 30132 5966 30144
rect 7009 30141 7021 30144
rect 7055 30141 7067 30175
rect 7009 30135 7067 30141
rect 7285 30175 7343 30181
rect 7285 30141 7297 30175
rect 7331 30172 7343 30175
rect 7742 30172 7748 30184
rect 7331 30144 7748 30172
rect 7331 30141 7343 30144
rect 7285 30135 7343 30141
rect 7742 30132 7748 30144
rect 7800 30132 7806 30184
rect 8018 30132 8024 30184
rect 8076 30172 8082 30184
rect 10778 30172 10784 30184
rect 8076 30144 10784 30172
rect 8076 30132 8082 30144
rect 10778 30132 10784 30144
rect 10836 30132 10842 30184
rect 10870 30132 10876 30184
rect 10928 30172 10934 30184
rect 11149 30175 11207 30181
rect 10928 30144 10973 30172
rect 10928 30132 10934 30144
rect 11149 30141 11161 30175
rect 11195 30141 11207 30175
rect 11698 30172 11704 30184
rect 11659 30144 11704 30172
rect 11149 30135 11207 30141
rect 1670 30104 1676 30116
rect 1631 30076 1676 30104
rect 1670 30064 1676 30076
rect 1728 30064 1734 30116
rect 3602 29996 3608 30048
rect 3660 30036 3666 30048
rect 3786 30036 3792 30048
rect 3660 30008 3792 30036
rect 3660 29996 3666 30008
rect 3786 29996 3792 30008
rect 3844 30036 3850 30048
rect 3881 30039 3939 30045
rect 3881 30036 3893 30039
rect 3844 30008 3893 30036
rect 3844 29996 3850 30008
rect 3881 30005 3893 30008
rect 3927 30005 3939 30039
rect 3881 29999 3939 30005
rect 7466 29996 7472 30048
rect 7524 30036 7530 30048
rect 7926 30036 7932 30048
rect 7524 30008 7932 30036
rect 7524 29996 7530 30008
rect 7926 29996 7932 30008
rect 7984 29996 7990 30048
rect 8757 30039 8815 30045
rect 8757 30005 8769 30039
rect 8803 30036 8815 30039
rect 10686 30036 10692 30048
rect 8803 30008 10692 30036
rect 8803 30005 8815 30008
rect 8757 29999 8815 30005
rect 10686 29996 10692 30008
rect 10744 29996 10750 30048
rect 10870 29996 10876 30048
rect 10928 30036 10934 30048
rect 11164 30036 11192 30135
rect 11698 30132 11704 30144
rect 11756 30132 11762 30184
rect 12526 30172 12532 30184
rect 11808 30144 12532 30172
rect 11514 30064 11520 30116
rect 11572 30104 11578 30116
rect 11808 30104 11836 30144
rect 12526 30132 12532 30144
rect 12584 30132 12590 30184
rect 13170 30172 13176 30184
rect 13131 30144 13176 30172
rect 13170 30132 13176 30144
rect 13228 30132 13234 30184
rect 13449 30175 13507 30181
rect 13449 30141 13461 30175
rect 13495 30141 13507 30175
rect 13449 30135 13507 30141
rect 11572 30076 11836 30104
rect 11572 30064 11578 30076
rect 12986 30036 12992 30048
rect 10928 30008 12992 30036
rect 10928 29996 10934 30008
rect 12986 29996 12992 30008
rect 13044 30036 13050 30048
rect 13464 30036 13492 30135
rect 14090 30132 14096 30184
rect 14148 30172 14154 30184
rect 14369 30175 14427 30181
rect 14369 30172 14381 30175
rect 14148 30144 14381 30172
rect 14148 30132 14154 30144
rect 14369 30141 14381 30144
rect 14415 30141 14427 30175
rect 14369 30135 14427 30141
rect 15013 30175 15071 30181
rect 15013 30141 15025 30175
rect 15059 30141 15071 30175
rect 15013 30135 15071 30141
rect 15933 30175 15991 30181
rect 15933 30141 15945 30175
rect 15979 30172 15991 30175
rect 16114 30172 16120 30184
rect 15979 30144 16120 30172
rect 15979 30141 15991 30144
rect 15933 30135 15991 30141
rect 14826 30064 14832 30116
rect 14884 30104 14890 30116
rect 15028 30104 15056 30135
rect 16114 30132 16120 30144
rect 16172 30132 16178 30184
rect 16209 30175 16267 30181
rect 16209 30141 16221 30175
rect 16255 30172 16267 30175
rect 16574 30172 16580 30184
rect 16255 30144 16580 30172
rect 16255 30141 16267 30144
rect 16209 30135 16267 30141
rect 16574 30132 16580 30144
rect 16632 30132 16638 30184
rect 16942 30172 16948 30184
rect 16903 30144 16948 30172
rect 16942 30132 16948 30144
rect 17000 30132 17006 30184
rect 17402 30172 17408 30184
rect 17363 30144 17408 30172
rect 17402 30132 17408 30144
rect 17460 30132 17466 30184
rect 14884 30076 15056 30104
rect 14884 30064 14890 30076
rect 16482 30064 16488 30116
rect 16540 30104 16546 30116
rect 17788 30104 17816 30212
rect 18049 30209 18061 30212
rect 18095 30209 18107 30243
rect 18049 30203 18107 30209
rect 18874 30200 18880 30252
rect 18932 30240 18938 30252
rect 18969 30243 19027 30249
rect 18969 30240 18981 30243
rect 18932 30212 18981 30240
rect 18932 30200 18938 30212
rect 18969 30209 18981 30212
rect 19015 30209 19027 30243
rect 19610 30240 19616 30252
rect 19523 30212 19616 30240
rect 18969 30203 19027 30209
rect 19610 30200 19616 30212
rect 19668 30200 19674 30252
rect 20257 30243 20315 30249
rect 20257 30209 20269 30243
rect 20303 30240 20315 30243
rect 20714 30240 20720 30252
rect 20303 30212 20720 30240
rect 20303 30209 20315 30212
rect 20257 30203 20315 30209
rect 20714 30200 20720 30212
rect 20772 30200 20778 30252
rect 29549 30243 29607 30249
rect 29549 30209 29561 30243
rect 29595 30240 29607 30243
rect 29595 30212 30144 30240
rect 29595 30209 29607 30212
rect 29549 30203 29607 30209
rect 17862 30132 17868 30184
rect 17920 30172 17926 30184
rect 19426 30172 19432 30184
rect 17920 30144 19432 30172
rect 17920 30132 17926 30144
rect 19426 30132 19432 30144
rect 19484 30132 19490 30184
rect 19628 30172 19656 30200
rect 22097 30175 22155 30181
rect 22097 30172 22109 30175
rect 19628 30144 22109 30172
rect 22097 30141 22109 30144
rect 22143 30172 22155 30175
rect 29178 30172 29184 30184
rect 22143 30144 29184 30172
rect 22143 30141 22155 30144
rect 22097 30135 22155 30141
rect 29178 30132 29184 30144
rect 29236 30132 29242 30184
rect 30116 30181 30144 30212
rect 37274 30200 37280 30252
rect 37332 30240 37338 30252
rect 38013 30243 38071 30249
rect 38013 30240 38025 30243
rect 37332 30212 38025 30240
rect 37332 30200 37338 30212
rect 38013 30209 38025 30212
rect 38059 30209 38071 30243
rect 38013 30203 38071 30209
rect 30101 30175 30159 30181
rect 30101 30141 30113 30175
rect 30147 30172 30159 30175
rect 37642 30172 37648 30184
rect 30147 30144 37648 30172
rect 30147 30141 30159 30144
rect 30101 30135 30159 30141
rect 37642 30132 37648 30144
rect 37700 30132 37706 30184
rect 20165 30107 20223 30113
rect 20165 30104 20177 30107
rect 16540 30076 17816 30104
rect 17880 30076 20177 30104
rect 16540 30064 16546 30076
rect 13044 30008 13492 30036
rect 13044 29996 13050 30008
rect 14734 29996 14740 30048
rect 14792 30036 14798 30048
rect 17880 30036 17908 30076
rect 20165 30073 20177 30076
rect 20211 30073 20223 30107
rect 20165 30067 20223 30073
rect 20346 30064 20352 30116
rect 20404 30104 20410 30116
rect 20809 30107 20867 30113
rect 20809 30104 20821 30107
rect 20404 30076 20821 30104
rect 20404 30064 20410 30076
rect 20809 30073 20821 30076
rect 20855 30104 20867 30107
rect 22557 30107 22615 30113
rect 22557 30104 22569 30107
rect 20855 30076 22569 30104
rect 20855 30073 20867 30076
rect 20809 30067 20867 30073
rect 22557 30073 22569 30076
rect 22603 30073 22615 30107
rect 22557 30067 22615 30073
rect 14792 30008 17908 30036
rect 18141 30039 18199 30045
rect 14792 29996 14798 30008
rect 18141 30005 18153 30039
rect 18187 30036 18199 30039
rect 18230 30036 18236 30048
rect 18187 30008 18236 30036
rect 18187 30005 18199 30008
rect 18141 29999 18199 30005
rect 18230 29996 18236 30008
rect 18288 29996 18294 30048
rect 18690 29996 18696 30048
rect 18748 30036 18754 30048
rect 18877 30039 18935 30045
rect 18877 30036 18889 30039
rect 18748 30008 18889 30036
rect 18748 29996 18754 30008
rect 18877 30005 18889 30008
rect 18923 30005 18935 30039
rect 18877 29999 18935 30005
rect 18966 29996 18972 30048
rect 19024 30036 19030 30048
rect 19521 30039 19579 30045
rect 19521 30036 19533 30039
rect 19024 30008 19533 30036
rect 19024 29996 19030 30008
rect 19521 30005 19533 30008
rect 19567 30005 19579 30039
rect 19521 29999 19579 30005
rect 20254 29996 20260 30048
rect 20312 30036 20318 30048
rect 21269 30039 21327 30045
rect 21269 30036 21281 30039
rect 20312 30008 21281 30036
rect 20312 29996 20318 30008
rect 21269 30005 21281 30008
rect 21315 30005 21327 30039
rect 29454 30036 29460 30048
rect 29415 30008 29460 30036
rect 21269 29999 21327 30005
rect 29454 29996 29460 30008
rect 29512 29996 29518 30048
rect 38194 30036 38200 30048
rect 38155 30008 38200 30036
rect 38194 29996 38200 30008
rect 38252 29996 38258 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 1936 29835 1994 29841
rect 1936 29801 1948 29835
rect 1982 29832 1994 29835
rect 1982 29804 3832 29832
rect 1982 29801 1994 29804
rect 1936 29795 1994 29801
rect 3804 29764 3832 29804
rect 3878 29792 3884 29844
rect 3936 29832 3942 29844
rect 3973 29835 4031 29841
rect 3973 29832 3985 29835
rect 3936 29804 3985 29832
rect 3936 29792 3942 29804
rect 3973 29801 3985 29804
rect 4019 29801 4031 29835
rect 4798 29832 4804 29844
rect 3973 29795 4031 29801
rect 4080 29804 4804 29832
rect 4080 29764 4108 29804
rect 4798 29792 4804 29804
rect 4856 29792 4862 29844
rect 7742 29792 7748 29844
rect 7800 29832 7806 29844
rect 8018 29832 8024 29844
rect 7800 29804 8024 29832
rect 7800 29792 7806 29804
rect 8018 29792 8024 29804
rect 8076 29792 8082 29844
rect 8386 29792 8392 29844
rect 8444 29832 8450 29844
rect 9582 29832 9588 29844
rect 8444 29804 9588 29832
rect 8444 29792 8450 29804
rect 9582 29792 9588 29804
rect 9640 29792 9646 29844
rect 9950 29832 9956 29844
rect 9784 29804 9956 29832
rect 9674 29764 9680 29776
rect 3804 29736 4108 29764
rect 8404 29736 9680 29764
rect 3896 29708 3924 29736
rect 1673 29699 1731 29705
rect 1673 29665 1685 29699
rect 1719 29696 1731 29699
rect 3418 29696 3424 29708
rect 1719 29668 3424 29696
rect 1719 29665 1731 29668
rect 1673 29659 1731 29665
rect 3418 29656 3424 29668
rect 3476 29656 3482 29708
rect 3878 29656 3884 29708
rect 3936 29656 3942 29708
rect 5810 29696 5816 29708
rect 3988 29668 5816 29696
rect 3602 29588 3608 29640
rect 3660 29628 3666 29640
rect 3988 29628 4016 29668
rect 5810 29656 5816 29668
rect 5868 29656 5874 29708
rect 8404 29696 8432 29736
rect 9674 29724 9680 29736
rect 9732 29724 9738 29776
rect 9784 29773 9812 29804
rect 9950 29792 9956 29804
rect 10008 29832 10014 29844
rect 10008 29804 12020 29832
rect 10008 29792 10014 29804
rect 9769 29767 9827 29773
rect 9769 29733 9781 29767
rect 9815 29733 9827 29767
rect 9769 29727 9827 29733
rect 10410 29724 10416 29776
rect 10468 29764 10474 29776
rect 10468 29736 10732 29764
rect 10468 29724 10474 29736
rect 6748 29668 8432 29696
rect 8481 29699 8539 29705
rect 3660 29600 4016 29628
rect 5721 29631 5779 29637
rect 3660 29588 3666 29600
rect 5721 29597 5733 29631
rect 5767 29628 5779 29631
rect 5902 29628 5908 29640
rect 5767 29600 5908 29628
rect 5767 29597 5779 29600
rect 5721 29591 5779 29597
rect 5902 29588 5908 29600
rect 5960 29588 5966 29640
rect 3970 29560 3976 29572
rect 3174 29532 3976 29560
rect 3970 29520 3976 29532
rect 4028 29520 4034 29572
rect 4706 29520 4712 29572
rect 4764 29520 4770 29572
rect 5445 29563 5503 29569
rect 5445 29529 5457 29563
rect 5491 29560 5503 29563
rect 6362 29560 6368 29572
rect 5491 29532 6368 29560
rect 5491 29529 5503 29532
rect 5445 29523 5503 29529
rect 6362 29520 6368 29532
rect 6420 29560 6426 29572
rect 6748 29560 6776 29668
rect 8481 29665 8493 29699
rect 8527 29696 8539 29699
rect 10597 29699 10655 29705
rect 10597 29696 10609 29699
rect 8527 29668 10609 29696
rect 8527 29665 8539 29668
rect 8481 29659 8539 29665
rect 10597 29665 10609 29668
rect 10643 29665 10655 29699
rect 10704 29696 10732 29736
rect 10873 29699 10931 29705
rect 10873 29696 10885 29699
rect 10704 29668 10885 29696
rect 10597 29659 10655 29665
rect 10873 29665 10885 29668
rect 10919 29696 10931 29699
rect 11514 29696 11520 29708
rect 10919 29668 11520 29696
rect 10919 29665 10931 29668
rect 10873 29659 10931 29665
rect 7098 29588 7104 29640
rect 7156 29588 7162 29640
rect 6420 29532 6776 29560
rect 6420 29520 6426 29532
rect 3421 29495 3479 29501
rect 3421 29461 3433 29495
rect 3467 29492 3479 29495
rect 5534 29492 5540 29504
rect 3467 29464 5540 29492
rect 3467 29461 3479 29464
rect 3421 29455 3479 29461
rect 5534 29452 5540 29464
rect 5592 29452 5598 29504
rect 6748 29501 6776 29532
rect 8110 29520 8116 29572
rect 8168 29560 8174 29572
rect 8205 29563 8263 29569
rect 8205 29560 8217 29563
rect 8168 29532 8217 29560
rect 8168 29520 8174 29532
rect 8205 29529 8217 29532
rect 8251 29529 8263 29563
rect 9217 29563 9275 29569
rect 9217 29560 9229 29563
rect 8205 29523 8263 29529
rect 8312 29532 9229 29560
rect 6733 29495 6791 29501
rect 6733 29461 6745 29495
rect 6779 29461 6791 29495
rect 6733 29455 6791 29461
rect 6914 29452 6920 29504
rect 6972 29492 6978 29504
rect 8312 29492 8340 29532
rect 9217 29529 9229 29532
rect 9263 29529 9275 29563
rect 9217 29523 9275 29529
rect 9309 29563 9367 29569
rect 9309 29529 9321 29563
rect 9355 29560 9367 29563
rect 9398 29560 9404 29572
rect 9355 29532 9404 29560
rect 9355 29529 9367 29532
rect 9309 29523 9367 29529
rect 9398 29520 9404 29532
rect 9456 29520 9462 29572
rect 10612 29560 10640 29659
rect 11514 29656 11520 29668
rect 11572 29656 11578 29708
rect 11992 29696 12020 29804
rect 12526 29792 12532 29844
rect 12584 29832 12590 29844
rect 16482 29832 16488 29844
rect 12584 29804 16488 29832
rect 12584 29792 12590 29804
rect 16482 29792 16488 29804
rect 16540 29792 16546 29844
rect 16574 29792 16580 29844
rect 16632 29832 16638 29844
rect 16632 29804 19564 29832
rect 16632 29792 16638 29804
rect 12894 29724 12900 29776
rect 12952 29764 12958 29776
rect 14458 29764 14464 29776
rect 12952 29736 14464 29764
rect 12952 29724 12958 29736
rect 14458 29724 14464 29736
rect 14516 29724 14522 29776
rect 15930 29724 15936 29776
rect 15988 29764 15994 29776
rect 19426 29764 19432 29776
rect 15988 29736 19432 29764
rect 15988 29724 15994 29736
rect 19426 29724 19432 29736
rect 19484 29724 19490 29776
rect 19536 29764 19564 29804
rect 19610 29792 19616 29844
rect 19668 29832 19674 29844
rect 20165 29835 20223 29841
rect 20165 29832 20177 29835
rect 19668 29804 20177 29832
rect 19668 29792 19674 29804
rect 20165 29801 20177 29804
rect 20211 29801 20223 29835
rect 20806 29832 20812 29844
rect 20767 29804 20812 29832
rect 20165 29795 20223 29801
rect 20806 29792 20812 29804
rect 20864 29792 20870 29844
rect 21453 29835 21511 29841
rect 21453 29801 21465 29835
rect 21499 29832 21511 29835
rect 21542 29832 21548 29844
rect 21499 29804 21548 29832
rect 21499 29801 21511 29804
rect 21453 29795 21511 29801
rect 21542 29792 21548 29804
rect 21600 29792 21606 29844
rect 22554 29832 22560 29844
rect 22515 29804 22560 29832
rect 22554 29792 22560 29804
rect 22612 29792 22618 29844
rect 38010 29832 38016 29844
rect 37971 29804 38016 29832
rect 38010 29792 38016 29804
rect 38068 29792 38074 29844
rect 29454 29764 29460 29776
rect 19536 29736 29460 29764
rect 29454 29724 29460 29736
rect 29512 29724 29518 29776
rect 13633 29699 13691 29705
rect 13633 29696 13645 29699
rect 11992 29668 13645 29696
rect 13633 29665 13645 29668
rect 13679 29696 13691 29699
rect 14553 29699 14611 29705
rect 14553 29696 14565 29699
rect 13679 29668 14565 29696
rect 13679 29665 13691 29668
rect 13633 29659 13691 29665
rect 14553 29665 14565 29668
rect 14599 29665 14611 29699
rect 15562 29696 15568 29708
rect 15523 29668 15568 29696
rect 14553 29659 14611 29665
rect 15562 29656 15568 29668
rect 15620 29656 15626 29708
rect 21542 29696 21548 29708
rect 17972 29668 18828 29696
rect 17129 29631 17187 29637
rect 17129 29597 17141 29631
rect 17175 29628 17187 29631
rect 17310 29628 17316 29640
rect 17175 29600 17316 29628
rect 17175 29597 17187 29600
rect 17129 29591 17187 29597
rect 17310 29588 17316 29600
rect 17368 29588 17374 29640
rect 10870 29560 10876 29572
rect 10612 29532 10876 29560
rect 10870 29520 10876 29532
rect 10928 29520 10934 29572
rect 11514 29520 11520 29572
rect 11572 29520 11578 29572
rect 12989 29563 13047 29569
rect 12989 29529 13001 29563
rect 13035 29529 13047 29563
rect 12989 29523 13047 29529
rect 6972 29464 8340 29492
rect 6972 29452 6978 29464
rect 12250 29452 12256 29504
rect 12308 29492 12314 29504
rect 12345 29495 12403 29501
rect 12345 29492 12357 29495
rect 12308 29464 12357 29492
rect 12308 29452 12314 29464
rect 12345 29461 12357 29464
rect 12391 29492 12403 29495
rect 12434 29492 12440 29504
rect 12391 29464 12440 29492
rect 12391 29461 12403 29464
rect 12345 29455 12403 29461
rect 12434 29452 12440 29464
rect 12492 29452 12498 29504
rect 12802 29452 12808 29504
rect 12860 29492 12866 29504
rect 13004 29492 13032 29523
rect 13078 29520 13084 29572
rect 13136 29560 13142 29572
rect 13136 29532 13181 29560
rect 13136 29520 13142 29532
rect 13354 29520 13360 29572
rect 13412 29560 13418 29572
rect 14550 29560 14556 29572
rect 13412 29532 14556 29560
rect 13412 29520 13418 29532
rect 14550 29520 14556 29532
rect 14608 29520 14614 29572
rect 14645 29563 14703 29569
rect 14645 29529 14657 29563
rect 14691 29560 14703 29563
rect 14734 29560 14740 29572
rect 14691 29532 14740 29560
rect 14691 29529 14703 29532
rect 14645 29523 14703 29529
rect 14734 29520 14740 29532
rect 14792 29520 14798 29572
rect 14918 29520 14924 29572
rect 14976 29560 14982 29572
rect 16485 29563 16543 29569
rect 16485 29560 16497 29563
rect 14976 29532 16497 29560
rect 14976 29520 14982 29532
rect 16485 29529 16497 29532
rect 16531 29529 16543 29563
rect 16485 29523 16543 29529
rect 16577 29563 16635 29569
rect 16577 29529 16589 29563
rect 16623 29560 16635 29563
rect 17972 29560 18000 29668
rect 18800 29628 18828 29668
rect 20272 29668 21548 29696
rect 19334 29628 19340 29640
rect 18800 29600 19340 29628
rect 19306 29594 19340 29600
rect 19334 29588 19340 29594
rect 19392 29588 19398 29640
rect 19426 29588 19432 29640
rect 19484 29628 19490 29640
rect 20272 29637 20300 29668
rect 21542 29656 21548 29668
rect 21600 29656 21606 29708
rect 27338 29696 27344 29708
rect 22066 29668 27344 29696
rect 20257 29631 20315 29637
rect 19484 29600 19529 29628
rect 19484 29588 19490 29600
rect 20257 29597 20269 29631
rect 20303 29597 20315 29631
rect 20714 29628 20720 29640
rect 20675 29600 20720 29628
rect 20257 29591 20315 29597
rect 20714 29588 20720 29600
rect 20772 29588 20778 29640
rect 18138 29560 18144 29572
rect 16623 29532 18000 29560
rect 18099 29532 18144 29560
rect 16623 29529 16635 29532
rect 16577 29523 16635 29529
rect 18138 29520 18144 29532
rect 18196 29520 18202 29572
rect 18230 29520 18236 29572
rect 18288 29560 18294 29572
rect 18288 29532 18333 29560
rect 18288 29520 18294 29532
rect 18414 29520 18420 29572
rect 18472 29560 18478 29572
rect 18782 29560 18788 29572
rect 18472 29532 18788 29560
rect 18472 29520 18478 29532
rect 18782 29520 18788 29532
rect 18840 29520 18846 29572
rect 18874 29520 18880 29572
rect 18932 29560 18938 29572
rect 21913 29563 21971 29569
rect 21913 29560 21925 29563
rect 18932 29532 21925 29560
rect 18932 29520 18938 29532
rect 21913 29529 21925 29532
rect 21959 29560 21971 29563
rect 22066 29560 22094 29668
rect 27338 29656 27344 29668
rect 27396 29656 27402 29708
rect 37829 29631 37887 29637
rect 37829 29628 37841 29631
rect 21959 29532 22094 29560
rect 37660 29600 37841 29628
rect 21959 29529 21971 29532
rect 21913 29523 21971 29529
rect 37660 29504 37688 29600
rect 37829 29597 37841 29600
rect 37875 29597 37887 29631
rect 37829 29591 37887 29597
rect 15470 29492 15476 29504
rect 12860 29464 15476 29492
rect 12860 29452 12866 29464
rect 15470 29452 15476 29464
rect 15528 29452 15534 29504
rect 17494 29452 17500 29504
rect 17552 29492 17558 29504
rect 19521 29495 19579 29501
rect 19521 29492 19533 29495
rect 17552 29464 19533 29492
rect 17552 29452 17558 29464
rect 19521 29461 19533 29464
rect 19567 29461 19579 29495
rect 19521 29455 19579 29461
rect 37369 29495 37427 29501
rect 37369 29461 37381 29495
rect 37415 29492 37427 29495
rect 37642 29492 37648 29504
rect 37415 29464 37648 29492
rect 37415 29461 37427 29464
rect 37369 29455 37427 29461
rect 37642 29452 37648 29464
rect 37700 29452 37706 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 2685 29291 2743 29297
rect 2685 29257 2697 29291
rect 2731 29288 2743 29291
rect 5905 29291 5963 29297
rect 2731 29260 5396 29288
rect 2731 29257 2743 29260
rect 2685 29251 2743 29257
rect 1670 29220 1676 29232
rect 1631 29192 1676 29220
rect 1670 29180 1676 29192
rect 1728 29180 1734 29232
rect 3050 29180 3056 29232
rect 3108 29220 3114 29232
rect 5368 29220 5396 29260
rect 5905 29257 5917 29291
rect 5951 29288 5963 29291
rect 9490 29288 9496 29300
rect 5951 29260 9496 29288
rect 5951 29257 5963 29260
rect 5905 29251 5963 29257
rect 9490 29248 9496 29260
rect 9548 29248 9554 29300
rect 13354 29288 13360 29300
rect 10060 29260 13360 29288
rect 7926 29220 7932 29232
rect 3108 29192 3542 29220
rect 5368 29192 7932 29220
rect 3108 29180 3114 29192
rect 7926 29180 7932 29192
rect 7984 29180 7990 29232
rect 8202 29220 8208 29232
rect 8163 29192 8208 29220
rect 8202 29180 8208 29192
rect 8260 29180 8266 29232
rect 8386 29180 8392 29232
rect 8444 29220 8450 29232
rect 8757 29223 8815 29229
rect 8757 29220 8769 29223
rect 8444 29192 8769 29220
rect 8444 29180 8450 29192
rect 8757 29189 8769 29192
rect 8803 29189 8815 29223
rect 8757 29183 8815 29189
rect 9306 29180 9312 29232
rect 9364 29220 9370 29232
rect 9401 29223 9459 29229
rect 9401 29220 9413 29223
rect 9364 29192 9413 29220
rect 9364 29180 9370 29192
rect 9401 29189 9413 29192
rect 9447 29189 9459 29223
rect 9401 29183 9459 29189
rect 1762 29112 1768 29164
rect 1820 29152 1826 29164
rect 2593 29155 2651 29161
rect 2593 29152 2605 29155
rect 1820 29124 2605 29152
rect 1820 29112 1826 29124
rect 2593 29121 2605 29124
rect 2639 29121 2651 29155
rect 2593 29115 2651 29121
rect 5534 29112 5540 29164
rect 5592 29152 5598 29164
rect 5813 29155 5871 29161
rect 5813 29152 5825 29155
rect 5592 29124 5825 29152
rect 5592 29112 5598 29124
rect 5813 29121 5825 29124
rect 5859 29152 5871 29155
rect 5859 29124 6040 29152
rect 5859 29121 5871 29124
rect 5813 29115 5871 29121
rect 3142 29044 3148 29096
rect 3200 29084 3206 29096
rect 3237 29087 3295 29093
rect 3237 29084 3249 29087
rect 3200 29056 3249 29084
rect 3200 29044 3206 29056
rect 3237 29053 3249 29056
rect 3283 29084 3295 29087
rect 4985 29087 5043 29093
rect 3283 29056 4936 29084
rect 3283 29053 3295 29056
rect 3237 29047 3295 29053
rect 842 28976 848 29028
rect 900 29016 906 29028
rect 1857 29019 1915 29025
rect 1857 29016 1869 29019
rect 900 28988 1869 29016
rect 900 28976 906 28988
rect 1857 28985 1869 28988
rect 1903 28985 1915 29019
rect 4908 29016 4936 29056
rect 4985 29053 4997 29087
rect 5031 29084 5043 29087
rect 5902 29084 5908 29096
rect 5031 29056 5908 29084
rect 5031 29053 5043 29056
rect 4985 29047 5043 29053
rect 5902 29044 5908 29056
rect 5960 29044 5966 29096
rect 6012 29084 6040 29124
rect 6086 29112 6092 29164
rect 6144 29152 6150 29164
rect 7101 29155 7159 29161
rect 7101 29152 7113 29155
rect 6144 29124 7113 29152
rect 6144 29112 6150 29124
rect 7101 29121 7113 29124
rect 7147 29121 7159 29155
rect 7101 29115 7159 29121
rect 6270 29084 6276 29096
rect 6012 29056 6276 29084
rect 6270 29044 6276 29056
rect 6328 29044 6334 29096
rect 6914 29084 6920 29096
rect 6875 29056 6920 29084
rect 6914 29044 6920 29056
rect 6972 29044 6978 29096
rect 8113 29087 8171 29093
rect 8113 29053 8125 29087
rect 8159 29084 8171 29087
rect 9309 29087 9367 29093
rect 8159 29056 8708 29084
rect 8159 29053 8171 29056
rect 8113 29047 8171 29053
rect 8680 29028 8708 29056
rect 9309 29053 9321 29087
rect 9355 29084 9367 29087
rect 9398 29084 9404 29096
rect 9355 29056 9404 29084
rect 9355 29053 9367 29056
rect 9309 29047 9367 29053
rect 9398 29044 9404 29056
rect 9456 29084 9462 29096
rect 10060 29084 10088 29260
rect 13354 29248 13360 29260
rect 13412 29248 13418 29300
rect 16942 29288 16948 29300
rect 13924 29260 16948 29288
rect 10134 29180 10140 29232
rect 10192 29220 10198 29232
rect 10597 29223 10655 29229
rect 10597 29220 10609 29223
rect 10192 29192 10609 29220
rect 10192 29180 10198 29192
rect 10597 29189 10609 29192
rect 10643 29189 10655 29223
rect 10597 29183 10655 29189
rect 10870 29180 10876 29232
rect 10928 29220 10934 29232
rect 11974 29220 11980 29232
rect 10928 29192 11744 29220
rect 11935 29192 11980 29220
rect 10928 29180 10934 29192
rect 11146 29112 11152 29164
rect 11204 29152 11210 29164
rect 11716 29161 11744 29192
rect 11974 29180 11980 29192
rect 12032 29180 12038 29232
rect 13814 29220 13820 29232
rect 13202 29192 13820 29220
rect 13814 29180 13820 29192
rect 13872 29180 13878 29232
rect 11701 29155 11759 29161
rect 11204 29124 11249 29152
rect 11204 29112 11210 29124
rect 11701 29121 11713 29155
rect 11747 29121 11759 29155
rect 11701 29115 11759 29121
rect 9456 29056 10088 29084
rect 9456 29044 9462 29056
rect 10318 29044 10324 29096
rect 10376 29084 10382 29096
rect 10505 29087 10563 29093
rect 10505 29084 10517 29087
rect 10376 29056 10517 29084
rect 10376 29044 10382 29056
rect 10505 29053 10517 29056
rect 10551 29084 10563 29087
rect 13924 29084 13952 29260
rect 16942 29248 16948 29260
rect 17000 29248 17006 29300
rect 18874 29288 18880 29300
rect 17328 29260 18880 29288
rect 14182 29220 14188 29232
rect 14143 29192 14188 29220
rect 14182 29180 14188 29192
rect 14240 29180 14246 29232
rect 15378 29220 15384 29232
rect 15339 29192 15384 29220
rect 15378 29180 15384 29192
rect 15436 29180 15442 29232
rect 15933 29223 15991 29229
rect 15933 29189 15945 29223
rect 15979 29220 15991 29223
rect 16114 29220 16120 29232
rect 15979 29192 16120 29220
rect 15979 29189 15991 29192
rect 15933 29183 15991 29189
rect 16114 29180 16120 29192
rect 16172 29180 16178 29232
rect 16206 29180 16212 29232
rect 16264 29220 16270 29232
rect 17328 29220 17356 29260
rect 18874 29248 18880 29260
rect 18932 29248 18938 29300
rect 19613 29291 19671 29297
rect 19613 29257 19625 29291
rect 19659 29288 19671 29291
rect 22922 29288 22928 29300
rect 19659 29260 22928 29288
rect 19659 29257 19671 29260
rect 19613 29251 19671 29257
rect 22922 29248 22928 29260
rect 22980 29248 22986 29300
rect 17494 29220 17500 29232
rect 16264 29192 17356 29220
rect 17455 29192 17500 29220
rect 16264 29180 16270 29192
rect 17494 29180 17500 29192
rect 17552 29180 17558 29232
rect 17586 29180 17592 29232
rect 17644 29220 17650 29232
rect 18325 29223 18383 29229
rect 17644 29192 17689 29220
rect 17644 29180 17650 29192
rect 18325 29189 18337 29223
rect 18371 29220 18383 29223
rect 18966 29220 18972 29232
rect 18371 29192 18972 29220
rect 18371 29189 18383 29192
rect 18325 29183 18383 29189
rect 18966 29180 18972 29192
rect 19024 29180 19030 29232
rect 37366 29220 37372 29232
rect 19444 29192 20392 29220
rect 19444 29164 19472 29192
rect 19426 29152 19432 29164
rect 19387 29124 19432 29152
rect 19426 29112 19432 29124
rect 19484 29112 19490 29164
rect 20254 29152 20260 29164
rect 20215 29124 20260 29152
rect 20254 29112 20260 29124
rect 20312 29112 20318 29164
rect 20364 29152 20392 29192
rect 21376 29192 37372 29220
rect 20364 29124 20852 29152
rect 14090 29084 14096 29096
rect 10551 29056 13952 29084
rect 14052 29056 14096 29084
rect 10551 29053 10563 29056
rect 10505 29047 10563 29053
rect 14090 29044 14096 29056
rect 14148 29044 14154 29096
rect 15286 29084 15292 29096
rect 14200 29056 14780 29084
rect 15247 29056 15292 29084
rect 8202 29016 8208 29028
rect 4908 28988 5764 29016
rect 1857 28979 1915 28985
rect 3418 28908 3424 28960
rect 3476 28948 3482 28960
rect 4062 28948 4068 28960
rect 3476 28920 4068 28948
rect 3476 28908 3482 28920
rect 4062 28908 4068 28920
rect 4120 28908 4126 28960
rect 4727 28951 4785 28957
rect 4727 28917 4739 28951
rect 4773 28948 4785 28951
rect 5074 28948 5080 28960
rect 4773 28920 5080 28948
rect 4773 28917 4785 28920
rect 4727 28911 4785 28917
rect 5074 28908 5080 28920
rect 5132 28948 5138 28960
rect 5626 28948 5632 28960
rect 5132 28920 5632 28948
rect 5132 28908 5138 28920
rect 5626 28908 5632 28920
rect 5684 28908 5690 28960
rect 5736 28948 5764 28988
rect 6288 28988 8208 29016
rect 6288 28960 6316 28988
rect 8202 28976 8208 28988
rect 8260 28976 8266 29028
rect 8662 28976 8668 29028
rect 8720 29016 8726 29028
rect 9861 29019 9919 29025
rect 9861 29016 9873 29019
rect 8720 28988 9873 29016
rect 8720 28976 8726 28988
rect 9861 28985 9873 28988
rect 9907 28985 9919 29019
rect 9861 28979 9919 28985
rect 10226 28976 10232 29028
rect 10284 29016 10290 29028
rect 11238 29016 11244 29028
rect 10284 28988 11244 29016
rect 10284 28976 10290 28988
rect 11238 28976 11244 28988
rect 11296 28976 11302 29028
rect 13170 28976 13176 29028
rect 13228 29016 13234 29028
rect 13449 29019 13507 29025
rect 13449 29016 13461 29019
rect 13228 28988 13461 29016
rect 13228 28976 13234 28988
rect 13449 28985 13461 28988
rect 13495 29016 13507 29019
rect 13495 28988 13676 29016
rect 13495 28985 13507 28988
rect 13449 28979 13507 28985
rect 5810 28948 5816 28960
rect 5736 28920 5816 28948
rect 5810 28908 5816 28920
rect 5868 28908 5874 28960
rect 6270 28908 6276 28960
rect 6328 28908 6334 28960
rect 7561 28951 7619 28957
rect 7561 28917 7573 28951
rect 7607 28948 7619 28951
rect 7650 28948 7656 28960
rect 7607 28920 7656 28948
rect 7607 28917 7619 28920
rect 7561 28911 7619 28917
rect 7650 28908 7656 28920
rect 7708 28908 7714 28960
rect 7742 28908 7748 28960
rect 7800 28948 7806 28960
rect 10134 28948 10140 28960
rect 7800 28920 10140 28948
rect 7800 28908 7806 28920
rect 10134 28908 10140 28920
rect 10192 28908 10198 28960
rect 11974 28908 11980 28960
rect 12032 28948 12038 28960
rect 13354 28948 13360 28960
rect 12032 28920 13360 28948
rect 12032 28908 12038 28920
rect 13354 28908 13360 28920
rect 13412 28908 13418 28960
rect 13648 28948 13676 28988
rect 14200 28948 14228 29056
rect 14642 29016 14648 29028
rect 14603 28988 14648 29016
rect 14642 28976 14648 28988
rect 14700 28976 14706 29028
rect 14752 29016 14780 29056
rect 15286 29044 15292 29056
rect 15344 29044 15350 29096
rect 17310 29044 17316 29096
rect 17368 29084 17374 29096
rect 17862 29084 17868 29096
rect 17368 29056 17868 29084
rect 17368 29044 17374 29056
rect 17862 29044 17868 29056
rect 17920 29044 17926 29096
rect 18230 29084 18236 29096
rect 18191 29056 18236 29084
rect 18230 29044 18236 29056
rect 18288 29044 18294 29096
rect 18506 29084 18512 29096
rect 18467 29056 18512 29084
rect 18506 29044 18512 29056
rect 18564 29044 18570 29096
rect 20714 29084 20720 29096
rect 18616 29056 20720 29084
rect 18616 29016 18644 29056
rect 20714 29044 20720 29056
rect 20772 29044 20778 29096
rect 20824 29084 20852 29124
rect 20898 29112 20904 29164
rect 20956 29152 20962 29164
rect 21376 29161 21404 29192
rect 37366 29180 37372 29192
rect 37424 29180 37430 29232
rect 21361 29155 21419 29161
rect 21361 29152 21373 29155
rect 20956 29124 21373 29152
rect 20956 29112 20962 29124
rect 21361 29121 21373 29124
rect 21407 29121 21419 29155
rect 21361 29115 21419 29121
rect 34514 29112 34520 29164
rect 34572 29152 34578 29164
rect 38013 29155 38071 29161
rect 38013 29152 38025 29155
rect 34572 29124 38025 29152
rect 34572 29112 34578 29124
rect 38013 29121 38025 29124
rect 38059 29121 38071 29155
rect 38013 29115 38071 29121
rect 22005 29087 22063 29093
rect 22005 29084 22017 29087
rect 20824 29056 22017 29084
rect 22005 29053 22017 29056
rect 22051 29053 22063 29087
rect 22005 29047 22063 29053
rect 14752 28988 18644 29016
rect 18966 28976 18972 29028
rect 19024 29016 19030 29028
rect 20809 29019 20867 29025
rect 20809 29016 20821 29019
rect 19024 28988 20821 29016
rect 19024 28976 19030 28988
rect 20809 28985 20821 28988
rect 20855 28985 20867 29019
rect 38194 29016 38200 29028
rect 38155 28988 38200 29016
rect 20809 28979 20867 28985
rect 38194 28976 38200 28988
rect 38252 28976 38258 29028
rect 13648 28920 14228 28948
rect 16206 28908 16212 28960
rect 16264 28948 16270 28960
rect 20165 28951 20223 28957
rect 20165 28948 20177 28951
rect 16264 28920 20177 28948
rect 16264 28908 16270 28920
rect 20165 28917 20177 28920
rect 20211 28917 20223 28951
rect 20165 28911 20223 28917
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 2685 28747 2743 28753
rect 2685 28713 2697 28747
rect 2731 28744 2743 28747
rect 6914 28744 6920 28756
rect 2731 28716 6920 28744
rect 2731 28713 2743 28716
rect 2685 28707 2743 28713
rect 6914 28704 6920 28716
rect 6972 28704 6978 28756
rect 7558 28704 7564 28756
rect 7616 28744 7622 28756
rect 11882 28744 11888 28756
rect 7616 28716 11888 28744
rect 7616 28704 7622 28716
rect 11882 28704 11888 28716
rect 11940 28704 11946 28756
rect 13354 28704 13360 28756
rect 13412 28744 13418 28756
rect 16022 28744 16028 28756
rect 13412 28716 16028 28744
rect 13412 28704 13418 28716
rect 16022 28704 16028 28716
rect 16080 28704 16086 28756
rect 16850 28744 16856 28756
rect 16316 28716 16856 28744
rect 3329 28679 3387 28685
rect 3329 28645 3341 28679
rect 3375 28676 3387 28679
rect 9858 28676 9864 28688
rect 3375 28648 9864 28676
rect 3375 28645 3387 28648
rect 3329 28639 3387 28645
rect 9858 28636 9864 28648
rect 9916 28636 9922 28688
rect 9953 28679 10011 28685
rect 9953 28645 9965 28679
rect 9999 28676 10011 28679
rect 10962 28676 10968 28688
rect 9999 28648 10968 28676
rect 9999 28645 10011 28648
rect 9953 28639 10011 28645
rect 10962 28636 10968 28648
rect 11020 28676 11026 28688
rect 11698 28676 11704 28688
rect 11020 28648 11704 28676
rect 11020 28636 11026 28648
rect 11698 28636 11704 28648
rect 11756 28636 11762 28688
rect 11974 28636 11980 28688
rect 12032 28676 12038 28688
rect 13538 28676 13544 28688
rect 12032 28648 13544 28676
rect 12032 28636 12038 28648
rect 13538 28636 13544 28648
rect 13596 28636 13602 28688
rect 15562 28676 15568 28688
rect 14752 28648 15568 28676
rect 2041 28611 2099 28617
rect 2041 28577 2053 28611
rect 2087 28608 2099 28611
rect 2087 28580 3556 28608
rect 2087 28577 2099 28580
rect 2041 28571 2099 28577
rect 2133 28543 2191 28549
rect 2133 28509 2145 28543
rect 2179 28509 2191 28543
rect 2590 28540 2596 28552
rect 2551 28512 2596 28540
rect 2133 28503 2191 28509
rect 1854 28432 1860 28484
rect 1912 28472 1918 28484
rect 2148 28472 2176 28503
rect 2590 28500 2596 28512
rect 2648 28500 2654 28552
rect 3418 28540 3424 28552
rect 3379 28512 3424 28540
rect 3418 28500 3424 28512
rect 3476 28500 3482 28552
rect 2866 28472 2872 28484
rect 1912 28444 2872 28472
rect 1912 28432 1918 28444
rect 2866 28432 2872 28444
rect 2924 28432 2930 28484
rect 3528 28404 3556 28580
rect 4154 28568 4160 28620
rect 4212 28608 4218 28620
rect 6178 28608 6184 28620
rect 4212 28580 6184 28608
rect 4212 28568 4218 28580
rect 6178 28568 6184 28580
rect 6236 28568 6242 28620
rect 6549 28611 6607 28617
rect 6549 28577 6561 28611
rect 6595 28608 6607 28611
rect 7742 28608 7748 28620
rect 6595 28580 7748 28608
rect 6595 28577 6607 28580
rect 6549 28571 6607 28577
rect 7742 28568 7748 28580
rect 7800 28568 7806 28620
rect 7929 28611 7987 28617
rect 7929 28577 7941 28611
rect 7975 28608 7987 28611
rect 7975 28580 10088 28608
rect 7975 28577 7987 28580
rect 7929 28571 7987 28577
rect 7377 28543 7435 28549
rect 7377 28509 7389 28543
rect 7423 28540 7435 28543
rect 7558 28540 7564 28552
rect 7423 28512 7564 28540
rect 7423 28509 7435 28512
rect 7377 28503 7435 28509
rect 7558 28500 7564 28512
rect 7616 28500 7622 28552
rect 10060 28540 10088 28580
rect 10134 28568 10140 28620
rect 10192 28608 10198 28620
rect 10505 28611 10563 28617
rect 10505 28608 10517 28611
rect 10192 28580 10517 28608
rect 10192 28568 10198 28580
rect 10505 28577 10517 28580
rect 10551 28577 10563 28611
rect 10505 28571 10563 28577
rect 11238 28568 11244 28620
rect 11296 28608 11302 28620
rect 12618 28608 12624 28620
rect 11296 28580 11744 28608
rect 11296 28568 11302 28580
rect 10594 28540 10600 28552
rect 10060 28512 10600 28540
rect 10594 28500 10600 28512
rect 10652 28500 10658 28552
rect 11716 28540 11744 28580
rect 11900 28580 12624 28608
rect 11900 28540 11928 28580
rect 12618 28568 12624 28580
rect 12676 28568 12682 28620
rect 13449 28611 13507 28617
rect 13449 28577 13461 28611
rect 13495 28608 13507 28611
rect 14752 28608 14780 28648
rect 15562 28636 15568 28648
rect 15620 28676 15626 28688
rect 15930 28676 15936 28688
rect 15620 28648 15936 28676
rect 15620 28636 15626 28648
rect 15930 28636 15936 28648
rect 15988 28636 15994 28688
rect 13495 28580 14780 28608
rect 13495 28577 13507 28580
rect 13449 28571 13507 28577
rect 14826 28568 14832 28620
rect 14884 28608 14890 28620
rect 14921 28611 14979 28617
rect 14921 28608 14933 28611
rect 14884 28580 14933 28608
rect 14884 28568 14890 28580
rect 14921 28577 14933 28580
rect 14967 28577 14979 28611
rect 14921 28571 14979 28577
rect 16025 28611 16083 28617
rect 16025 28577 16037 28611
rect 16071 28608 16083 28611
rect 16114 28608 16120 28620
rect 16071 28580 16120 28608
rect 16071 28577 16083 28580
rect 16025 28571 16083 28577
rect 16114 28568 16120 28580
rect 16172 28568 16178 28620
rect 16316 28617 16344 28716
rect 16850 28704 16856 28716
rect 16908 28744 16914 28756
rect 17034 28744 17040 28756
rect 16908 28716 17040 28744
rect 16908 28704 16914 28716
rect 17034 28704 17040 28716
rect 17092 28704 17098 28756
rect 17310 28704 17316 28756
rect 17368 28744 17374 28756
rect 22830 28744 22836 28756
rect 17368 28716 22836 28744
rect 17368 28704 17374 28716
rect 22830 28704 22836 28716
rect 22888 28704 22894 28756
rect 33962 28744 33968 28756
rect 33923 28716 33968 28744
rect 33962 28704 33968 28716
rect 34020 28704 34026 28756
rect 16666 28636 16672 28688
rect 16724 28676 16730 28688
rect 20809 28679 20867 28685
rect 20809 28676 20821 28679
rect 16724 28648 20821 28676
rect 16724 28636 16730 28648
rect 20809 28645 20821 28648
rect 20855 28645 20867 28679
rect 20809 28639 20867 28645
rect 30929 28679 30987 28685
rect 30929 28645 30941 28679
rect 30975 28676 30987 28679
rect 34514 28676 34520 28688
rect 30975 28648 34520 28676
rect 30975 28645 30987 28648
rect 30929 28639 30987 28645
rect 34514 28636 34520 28648
rect 34572 28636 34578 28688
rect 16301 28611 16359 28617
rect 16301 28577 16313 28611
rect 16347 28577 16359 28611
rect 16942 28608 16948 28620
rect 16855 28580 16948 28608
rect 16301 28571 16359 28577
rect 16942 28568 16948 28580
rect 17000 28608 17006 28620
rect 18966 28608 18972 28620
rect 17000 28580 18972 28608
rect 17000 28568 17006 28580
rect 18966 28568 18972 28580
rect 19024 28568 19030 28620
rect 11716 28512 11928 28540
rect 19150 28500 19156 28552
rect 19208 28540 19214 28552
rect 20901 28543 20959 28549
rect 20901 28540 20913 28543
rect 19208 28512 20913 28540
rect 19208 28500 19214 28512
rect 20901 28509 20913 28512
rect 20947 28540 20959 28543
rect 21361 28543 21419 28549
rect 21361 28540 21373 28543
rect 20947 28512 21373 28540
rect 20947 28509 20959 28512
rect 20901 28503 20959 28509
rect 21361 28509 21373 28512
rect 21407 28509 21419 28543
rect 30742 28540 30748 28552
rect 30703 28512 30748 28540
rect 21361 28503 21419 28509
rect 30742 28500 30748 28512
rect 30800 28540 30806 28552
rect 31389 28543 31447 28549
rect 31389 28540 31401 28543
rect 30800 28512 31401 28540
rect 30800 28500 30806 28512
rect 31389 28509 31401 28512
rect 31435 28509 31447 28543
rect 34146 28540 34152 28552
rect 34107 28512 34152 28540
rect 31389 28503 31447 28509
rect 34146 28500 34152 28512
rect 34204 28540 34210 28552
rect 34885 28543 34943 28549
rect 34885 28540 34897 28543
rect 34204 28512 34897 28540
rect 34204 28500 34210 28512
rect 34885 28509 34897 28512
rect 34931 28509 34943 28543
rect 34885 28503 34943 28509
rect 4062 28472 4068 28484
rect 4023 28444 4068 28472
rect 4062 28432 4068 28444
rect 4120 28432 4126 28484
rect 4157 28475 4215 28481
rect 4157 28441 4169 28475
rect 4203 28441 4215 28475
rect 4157 28435 4215 28441
rect 4709 28475 4767 28481
rect 4709 28441 4721 28475
rect 4755 28472 4767 28475
rect 5074 28472 5080 28484
rect 4755 28444 5080 28472
rect 4755 28441 4767 28444
rect 4709 28435 4767 28441
rect 4172 28404 4200 28435
rect 5074 28432 5080 28444
rect 5132 28472 5138 28484
rect 5537 28475 5595 28481
rect 5537 28472 5549 28475
rect 5132 28444 5549 28472
rect 5132 28432 5138 28444
rect 5537 28441 5549 28444
rect 5583 28441 5595 28475
rect 5537 28435 5595 28441
rect 5629 28475 5687 28481
rect 5629 28441 5641 28475
rect 5675 28441 5687 28475
rect 5629 28435 5687 28441
rect 3528 28376 4200 28404
rect 4614 28364 4620 28416
rect 4672 28404 4678 28416
rect 5637 28404 5665 28435
rect 6638 28432 6644 28484
rect 6696 28472 6702 28484
rect 6696 28444 7880 28472
rect 6696 28432 6702 28444
rect 4672 28376 5665 28404
rect 4672 28364 4678 28376
rect 5718 28364 5724 28416
rect 5776 28404 5782 28416
rect 6270 28404 6276 28416
rect 5776 28376 6276 28404
rect 5776 28364 5782 28376
rect 6270 28364 6276 28376
rect 6328 28364 6334 28416
rect 7285 28407 7343 28413
rect 7285 28373 7297 28407
rect 7331 28404 7343 28407
rect 7742 28404 7748 28416
rect 7331 28376 7748 28404
rect 7331 28373 7343 28376
rect 7285 28367 7343 28373
rect 7742 28364 7748 28376
rect 7800 28364 7806 28416
rect 7852 28404 7880 28444
rect 7926 28432 7932 28484
rect 7984 28472 7990 28484
rect 8021 28475 8079 28481
rect 8021 28472 8033 28475
rect 7984 28444 8033 28472
rect 7984 28432 7990 28444
rect 8021 28441 8033 28444
rect 8067 28441 8079 28475
rect 8021 28435 8079 28441
rect 8386 28432 8392 28484
rect 8444 28472 8450 28484
rect 8573 28475 8631 28481
rect 8573 28472 8585 28475
rect 8444 28444 8585 28472
rect 8444 28432 8450 28444
rect 8573 28441 8585 28444
rect 8619 28441 8631 28475
rect 9398 28472 9404 28484
rect 9359 28444 9404 28472
rect 8573 28435 8631 28441
rect 9398 28432 9404 28444
rect 9456 28432 9462 28484
rect 9490 28432 9496 28484
rect 9548 28472 9554 28484
rect 11422 28472 11428 28484
rect 9548 28444 9593 28472
rect 11383 28444 11428 28472
rect 9548 28432 9554 28444
rect 11422 28432 11428 28444
rect 11480 28432 11486 28484
rect 11514 28432 11520 28484
rect 11572 28472 11578 28484
rect 11572 28444 11617 28472
rect 11572 28432 11578 28444
rect 11698 28432 11704 28484
rect 11756 28472 11762 28484
rect 12529 28475 12587 28481
rect 12529 28472 12541 28475
rect 11756 28444 12541 28472
rect 11756 28432 11762 28444
rect 12529 28441 12541 28444
rect 12575 28441 12587 28475
rect 12529 28435 12587 28441
rect 12618 28432 12624 28484
rect 12676 28472 12682 28484
rect 12676 28444 12721 28472
rect 12676 28432 12682 28444
rect 13630 28432 13636 28484
rect 13688 28472 13694 28484
rect 14277 28475 14335 28481
rect 14277 28472 14289 28475
rect 13688 28444 14289 28472
rect 13688 28432 13694 28444
rect 14277 28441 14289 28444
rect 14323 28441 14335 28475
rect 14277 28435 14335 28441
rect 14829 28475 14887 28481
rect 14829 28441 14841 28475
rect 14875 28441 14887 28475
rect 16206 28472 16212 28484
rect 16167 28444 16212 28472
rect 14829 28435 14887 28441
rect 10318 28404 10324 28416
rect 7852 28376 10324 28404
rect 10318 28364 10324 28376
rect 10376 28364 10382 28416
rect 11054 28364 11060 28416
rect 11112 28404 11118 28416
rect 14844 28404 14872 28435
rect 16206 28432 16212 28444
rect 16264 28432 16270 28484
rect 17037 28475 17095 28481
rect 17037 28441 17049 28475
rect 17083 28441 17095 28475
rect 17037 28435 17095 28441
rect 17589 28475 17647 28481
rect 17589 28441 17601 28475
rect 17635 28441 17647 28475
rect 17589 28435 17647 28441
rect 18141 28475 18199 28481
rect 18141 28441 18153 28475
rect 18187 28472 18199 28475
rect 18506 28472 18512 28484
rect 18187 28444 18512 28472
rect 18187 28441 18199 28444
rect 18141 28435 18199 28441
rect 11112 28376 14872 28404
rect 11112 28364 11118 28376
rect 16390 28364 16396 28416
rect 16448 28404 16454 28416
rect 17052 28404 17080 28435
rect 16448 28376 17080 28404
rect 17604 28404 17632 28435
rect 18506 28432 18512 28444
rect 18564 28432 18570 28484
rect 18690 28472 18696 28484
rect 18651 28444 18696 28472
rect 18690 28432 18696 28444
rect 18748 28432 18754 28484
rect 18785 28475 18843 28481
rect 18785 28441 18797 28475
rect 18831 28472 18843 28475
rect 19242 28472 19248 28484
rect 18831 28444 19248 28472
rect 18831 28441 18843 28444
rect 18785 28435 18843 28441
rect 19242 28432 19248 28444
rect 19300 28432 19306 28484
rect 18230 28404 18236 28416
rect 17604 28376 18236 28404
rect 16448 28364 16454 28376
rect 18230 28364 18236 28376
rect 18288 28404 18294 28416
rect 18414 28404 18420 28416
rect 18288 28376 18420 28404
rect 18288 28364 18294 28376
rect 18414 28364 18420 28376
rect 18472 28364 18478 28416
rect 19613 28407 19671 28413
rect 19613 28373 19625 28407
rect 19659 28404 19671 28407
rect 19978 28404 19984 28416
rect 19659 28376 19984 28404
rect 19659 28373 19671 28376
rect 19613 28367 19671 28373
rect 19978 28364 19984 28376
rect 20036 28364 20042 28416
rect 20070 28364 20076 28416
rect 20128 28404 20134 28416
rect 20128 28376 20173 28404
rect 20128 28364 20134 28376
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 2685 28203 2743 28209
rect 2685 28169 2697 28203
rect 2731 28169 2743 28203
rect 2685 28163 2743 28169
rect 2700 28132 2728 28163
rect 4062 28160 4068 28212
rect 4120 28200 4126 28212
rect 4525 28203 4583 28209
rect 4525 28200 4537 28203
rect 4120 28172 4537 28200
rect 4120 28160 4126 28172
rect 4525 28169 4537 28172
rect 4571 28169 4583 28203
rect 4525 28163 4583 28169
rect 5261 28203 5319 28209
rect 5261 28169 5273 28203
rect 5307 28200 5319 28203
rect 5307 28172 7880 28200
rect 5307 28169 5319 28172
rect 5261 28163 5319 28169
rect 4982 28132 4988 28144
rect 2700 28104 4988 28132
rect 4982 28092 4988 28104
rect 5040 28092 5046 28144
rect 5534 28092 5540 28144
rect 5592 28132 5598 28144
rect 7745 28135 7803 28141
rect 7745 28132 7757 28135
rect 5592 28104 7757 28132
rect 5592 28092 5598 28104
rect 7745 28101 7757 28104
rect 7791 28101 7803 28135
rect 7852 28132 7880 28172
rect 9582 28160 9588 28212
rect 9640 28200 9646 28212
rect 11974 28200 11980 28212
rect 9640 28172 11980 28200
rect 9640 28160 9646 28172
rect 11974 28160 11980 28172
rect 12032 28160 12038 28212
rect 16209 28203 16267 28209
rect 16209 28169 16221 28203
rect 16255 28200 16267 28203
rect 16390 28200 16396 28212
rect 16255 28172 16396 28200
rect 16255 28169 16267 28172
rect 16209 28163 16267 28169
rect 16390 28160 16396 28172
rect 16448 28160 16454 28212
rect 18138 28160 18144 28212
rect 18196 28200 18202 28212
rect 18233 28203 18291 28209
rect 18233 28200 18245 28203
rect 18196 28172 18245 28200
rect 18196 28160 18202 28172
rect 18233 28169 18245 28172
rect 18279 28169 18291 28203
rect 21085 28203 21143 28209
rect 21085 28200 21097 28203
rect 18233 28163 18291 28169
rect 18340 28172 21097 28200
rect 9401 28135 9459 28141
rect 9401 28132 9413 28135
rect 7852 28104 9413 28132
rect 7745 28095 7803 28101
rect 9401 28101 9413 28104
rect 9447 28101 9459 28135
rect 9401 28095 9459 28101
rect 9674 28092 9680 28144
rect 9732 28132 9738 28144
rect 10597 28135 10655 28141
rect 10597 28132 10609 28135
rect 9732 28104 10609 28132
rect 9732 28092 9738 28104
rect 10597 28101 10609 28104
rect 10643 28101 10655 28135
rect 10597 28095 10655 28101
rect 10686 28092 10692 28144
rect 10744 28132 10750 28144
rect 12897 28135 12955 28141
rect 12897 28132 12909 28135
rect 10744 28104 12909 28132
rect 10744 28092 10750 28104
rect 12897 28101 12909 28104
rect 12943 28101 12955 28135
rect 12897 28095 12955 28101
rect 13449 28135 13507 28141
rect 13449 28101 13461 28135
rect 13495 28132 13507 28135
rect 13630 28132 13636 28144
rect 13495 28104 13636 28132
rect 13495 28101 13507 28104
rect 13449 28095 13507 28101
rect 1857 28067 1915 28073
rect 1857 28033 1869 28067
rect 1903 28064 1915 28067
rect 2314 28064 2320 28076
rect 1903 28036 2320 28064
rect 1903 28033 1915 28036
rect 1857 28027 1915 28033
rect 2314 28024 2320 28036
rect 2372 28024 2378 28076
rect 2501 28067 2559 28073
rect 2501 28033 2513 28067
rect 2547 28033 2559 28067
rect 3326 28064 3332 28076
rect 3287 28036 3332 28064
rect 2501 28027 2559 28033
rect 2516 27996 2544 28027
rect 3326 28024 3332 28036
rect 3384 28024 3390 28076
rect 3973 28067 4031 28073
rect 3973 28033 3985 28067
rect 4019 28064 4031 28067
rect 4062 28064 4068 28076
rect 4019 28036 4068 28064
rect 4019 28033 4031 28036
rect 3973 28027 4031 28033
rect 4062 28024 4068 28036
rect 4120 28024 4126 28076
rect 4522 28064 4528 28076
rect 4483 28036 4528 28064
rect 4522 28024 4528 28036
rect 4580 28024 4586 28076
rect 5169 28067 5227 28073
rect 5169 28033 5181 28067
rect 5215 28064 5227 28067
rect 5442 28064 5448 28076
rect 5215 28036 5448 28064
rect 5215 28033 5227 28036
rect 5169 28027 5227 28033
rect 5442 28024 5448 28036
rect 5500 28024 5506 28076
rect 5813 28067 5871 28073
rect 5813 28033 5825 28067
rect 5859 28033 5871 28067
rect 5813 28027 5871 28033
rect 5905 28067 5963 28073
rect 5905 28033 5917 28067
rect 5951 28064 5963 28067
rect 6638 28064 6644 28076
rect 5951 28036 6644 28064
rect 5951 28033 5963 28036
rect 5905 28027 5963 28033
rect 3142 27996 3148 28008
rect 2516 27968 3148 27996
rect 3142 27956 3148 27968
rect 3200 27956 3206 28008
rect 3237 27999 3295 28005
rect 3237 27965 3249 27999
rect 3283 27996 3295 27999
rect 5718 27996 5724 28008
rect 3283 27968 5724 27996
rect 3283 27965 3295 27968
rect 3237 27959 3295 27965
rect 5718 27956 5724 27968
rect 5776 27956 5782 28008
rect 5828 27996 5856 28027
rect 6638 28024 6644 28036
rect 6696 28024 6702 28076
rect 6914 28064 6920 28076
rect 6827 28036 6920 28064
rect 6914 28024 6920 28036
rect 6972 28064 6978 28076
rect 7466 28064 7472 28076
rect 6972 28036 7472 28064
rect 6972 28024 6978 28036
rect 7466 28024 7472 28036
rect 7524 28024 7530 28076
rect 9950 28024 9956 28076
rect 10008 28064 10014 28076
rect 12250 28064 12256 28076
rect 10008 28036 10053 28064
rect 12211 28036 12256 28064
rect 10008 28024 10014 28036
rect 12250 28024 12256 28036
rect 12308 28024 12314 28076
rect 6178 27996 6184 28008
rect 5828 27968 6184 27996
rect 6178 27956 6184 27968
rect 6236 27956 6242 28008
rect 7650 27956 7656 28008
rect 7708 27996 7714 28008
rect 8297 27999 8355 28005
rect 7708 27968 7753 27996
rect 7708 27956 7714 27968
rect 8297 27965 8309 27999
rect 8343 27996 8355 27999
rect 8386 27996 8392 28008
rect 8343 27968 8392 27996
rect 8343 27965 8355 27968
rect 8297 27959 8355 27965
rect 8386 27956 8392 27968
rect 8444 27956 8450 28008
rect 9030 27956 9036 28008
rect 9088 27996 9094 28008
rect 9309 27999 9367 28005
rect 9309 27996 9321 27999
rect 9088 27968 9321 27996
rect 9088 27956 9094 27968
rect 9309 27965 9321 27968
rect 9355 27965 9367 27999
rect 9309 27959 9367 27965
rect 10318 27956 10324 28008
rect 10376 27996 10382 28008
rect 10505 27999 10563 28005
rect 10505 27996 10517 27999
rect 10376 27968 10517 27996
rect 10376 27956 10382 27968
rect 10505 27965 10517 27968
rect 10551 27965 10563 27999
rect 10505 27959 10563 27965
rect 12805 27999 12863 28005
rect 12805 27965 12817 27999
rect 12851 27996 12863 27999
rect 12894 27996 12900 28008
rect 12851 27968 12900 27996
rect 12851 27965 12863 27968
rect 12805 27959 12863 27965
rect 12894 27956 12900 27968
rect 12952 27956 12958 28008
rect 1670 27928 1676 27940
rect 1631 27900 1676 27928
rect 1670 27888 1676 27900
rect 1728 27888 1734 27940
rect 3881 27931 3939 27937
rect 3881 27897 3893 27931
rect 3927 27928 3939 27931
rect 7558 27928 7564 27940
rect 3927 27900 7564 27928
rect 3927 27897 3939 27900
rect 3881 27891 3939 27897
rect 7558 27888 7564 27900
rect 7616 27888 7622 27940
rect 10778 27928 10784 27940
rect 9646 27900 10784 27928
rect 5902 27820 5908 27872
rect 5960 27860 5966 27872
rect 6546 27860 6552 27872
rect 5960 27832 6552 27860
rect 5960 27820 5966 27832
rect 6546 27820 6552 27832
rect 6604 27820 6610 27872
rect 7009 27863 7067 27869
rect 7009 27829 7021 27863
rect 7055 27860 7067 27863
rect 9646 27860 9674 27900
rect 10778 27888 10784 27900
rect 10836 27888 10842 27940
rect 11054 27928 11060 27940
rect 11015 27900 11060 27928
rect 11054 27888 11060 27900
rect 11112 27928 11118 27940
rect 13464 27928 13492 28095
rect 13630 28092 13636 28104
rect 13688 28092 13694 28144
rect 14274 28132 14280 28144
rect 14235 28104 14280 28132
rect 14274 28092 14280 28104
rect 14332 28092 14338 28144
rect 14458 28092 14464 28144
rect 14516 28132 14522 28144
rect 14516 28104 16160 28132
rect 14516 28092 14522 28104
rect 15473 28067 15531 28073
rect 15473 28033 15485 28067
rect 15519 28064 15531 28067
rect 16022 28064 16028 28076
rect 15519 28036 16028 28064
rect 15519 28033 15531 28036
rect 15473 28027 15531 28033
rect 16022 28024 16028 28036
rect 16080 28024 16086 28076
rect 16132 28073 16160 28104
rect 16574 28092 16580 28144
rect 16632 28132 16638 28144
rect 17037 28135 17095 28141
rect 17037 28132 17049 28135
rect 16632 28104 17049 28132
rect 16632 28092 16638 28104
rect 17037 28101 17049 28104
rect 17083 28101 17095 28135
rect 17037 28095 17095 28101
rect 16117 28067 16175 28073
rect 16117 28033 16129 28067
rect 16163 28064 16175 28067
rect 16482 28064 16488 28076
rect 16163 28036 16488 28064
rect 16163 28033 16175 28036
rect 16117 28027 16175 28033
rect 16482 28024 16488 28036
rect 16540 28024 16546 28076
rect 18340 28073 18368 28172
rect 21085 28169 21097 28172
rect 21131 28200 21143 28203
rect 23566 28200 23572 28212
rect 21131 28172 23572 28200
rect 21131 28169 21143 28172
rect 21085 28163 21143 28169
rect 23566 28160 23572 28172
rect 23624 28160 23630 28212
rect 18598 28092 18604 28144
rect 18656 28132 18662 28144
rect 18969 28135 19027 28141
rect 18969 28132 18981 28135
rect 18656 28104 18981 28132
rect 18656 28092 18662 28104
rect 18969 28101 18981 28104
rect 19015 28101 19027 28135
rect 18969 28095 19027 28101
rect 22097 28135 22155 28141
rect 22097 28101 22109 28135
rect 22143 28132 22155 28135
rect 22646 28132 22652 28144
rect 22143 28104 22652 28132
rect 22143 28101 22155 28104
rect 22097 28095 22155 28101
rect 22646 28092 22652 28104
rect 22704 28092 22710 28144
rect 18325 28067 18383 28073
rect 18325 28033 18337 28067
rect 18371 28033 18383 28067
rect 19978 28064 19984 28076
rect 19939 28036 19984 28064
rect 18325 28027 18383 28033
rect 19978 28024 19984 28036
rect 20036 28024 20042 28076
rect 14185 27999 14243 28005
rect 14185 27965 14197 27999
rect 14231 27965 14243 27999
rect 14642 27996 14648 28008
rect 14603 27968 14648 27996
rect 14185 27959 14243 27965
rect 11112 27900 13492 27928
rect 14200 27928 14228 27959
rect 14642 27956 14648 27968
rect 14700 27956 14706 28008
rect 15010 27956 15016 28008
rect 15068 27996 15074 28008
rect 16942 27996 16948 28008
rect 15068 27968 16804 27996
rect 16903 27968 16948 27996
rect 15068 27956 15074 27968
rect 15562 27928 15568 27940
rect 14200 27900 15568 27928
rect 11112 27888 11118 27900
rect 15562 27888 15568 27900
rect 15620 27888 15626 27940
rect 7055 27832 9674 27860
rect 12161 27863 12219 27869
rect 7055 27829 7067 27832
rect 7009 27823 7067 27829
rect 12161 27829 12173 27863
rect 12207 27860 12219 27863
rect 14366 27860 14372 27872
rect 12207 27832 14372 27860
rect 12207 27829 12219 27832
rect 12161 27823 12219 27829
rect 14366 27820 14372 27832
rect 14424 27820 14430 27872
rect 15194 27820 15200 27872
rect 15252 27860 15258 27872
rect 15381 27863 15439 27869
rect 15381 27860 15393 27863
rect 15252 27832 15393 27860
rect 15252 27820 15258 27832
rect 15381 27829 15393 27832
rect 15427 27829 15439 27863
rect 16776 27860 16804 27968
rect 16942 27956 16948 27968
rect 17000 27956 17006 28008
rect 17221 27999 17279 28005
rect 17221 27965 17233 27999
rect 17267 27996 17279 27999
rect 18690 27996 18696 28008
rect 17267 27968 18696 27996
rect 17267 27965 17279 27968
rect 17221 27959 17279 27965
rect 16850 27888 16856 27940
rect 16908 27928 16914 27940
rect 17236 27928 17264 27959
rect 18690 27956 18696 27968
rect 18748 27956 18754 28008
rect 18874 27996 18880 28008
rect 18835 27968 18880 27996
rect 18874 27956 18880 27968
rect 18932 27956 18938 28008
rect 19334 27956 19340 28008
rect 19392 27996 19398 28008
rect 20165 27999 20223 28005
rect 20165 27996 20177 27999
rect 19392 27968 20177 27996
rect 19392 27956 19398 27968
rect 20165 27965 20177 27968
rect 20211 27965 20223 27999
rect 20165 27959 20223 27965
rect 16908 27900 17264 27928
rect 16908 27888 16914 27900
rect 18506 27888 18512 27940
rect 18564 27928 18570 27940
rect 19429 27931 19487 27937
rect 19429 27928 19441 27931
rect 18564 27900 19441 27928
rect 18564 27888 18570 27900
rect 19429 27897 19441 27900
rect 19475 27928 19487 27931
rect 26234 27928 26240 27940
rect 19475 27900 26240 27928
rect 19475 27897 19487 27900
rect 19429 27891 19487 27897
rect 26234 27888 26240 27900
rect 26292 27888 26298 27940
rect 19150 27860 19156 27872
rect 16776 27832 19156 27860
rect 15381 27823 15439 27829
rect 19150 27820 19156 27832
rect 19208 27820 19214 27872
rect 19242 27820 19248 27872
rect 19300 27860 19306 27872
rect 20349 27863 20407 27869
rect 20349 27860 20361 27863
rect 19300 27832 20361 27860
rect 19300 27820 19306 27832
rect 20349 27829 20361 27832
rect 20395 27829 20407 27863
rect 20349 27823 20407 27829
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 2866 27616 2872 27668
rect 2924 27656 2930 27668
rect 8110 27656 8116 27668
rect 2924 27628 8116 27656
rect 2924 27616 2930 27628
rect 8110 27616 8116 27628
rect 8168 27616 8174 27668
rect 8481 27659 8539 27665
rect 8481 27625 8493 27659
rect 8527 27656 8539 27659
rect 10686 27656 10692 27668
rect 8527 27628 10692 27656
rect 8527 27625 8539 27628
rect 8481 27619 8539 27625
rect 10686 27616 10692 27628
rect 10744 27616 10750 27668
rect 11514 27616 11520 27668
rect 11572 27656 11578 27668
rect 16850 27656 16856 27668
rect 11572 27628 16856 27656
rect 11572 27616 11578 27628
rect 16850 27616 16856 27628
rect 16908 27616 16914 27668
rect 18874 27656 18880 27668
rect 18835 27628 18880 27656
rect 18874 27616 18880 27628
rect 18932 27616 18938 27668
rect 22373 27659 22431 27665
rect 22373 27625 22385 27659
rect 22419 27656 22431 27659
rect 22646 27656 22652 27668
rect 22419 27628 22652 27656
rect 22419 27625 22431 27628
rect 22373 27619 22431 27625
rect 22646 27616 22652 27628
rect 22704 27616 22710 27668
rect 22830 27656 22836 27668
rect 22791 27628 22836 27656
rect 22830 27616 22836 27628
rect 22888 27616 22894 27668
rect 1949 27591 2007 27597
rect 1949 27557 1961 27591
rect 1995 27588 2007 27591
rect 2038 27588 2044 27600
rect 1995 27560 2044 27588
rect 1995 27557 2007 27560
rect 1949 27551 2007 27557
rect 2038 27548 2044 27560
rect 2096 27548 2102 27600
rect 2685 27591 2743 27597
rect 2685 27557 2697 27591
rect 2731 27588 2743 27591
rect 4614 27588 4620 27600
rect 2731 27560 4620 27588
rect 2731 27557 2743 27560
rect 2685 27551 2743 27557
rect 4614 27548 4620 27560
rect 4672 27548 4678 27600
rect 10318 27588 10324 27600
rect 5368 27560 10324 27588
rect 2866 27480 2872 27532
rect 2924 27520 2930 27532
rect 5368 27529 5396 27560
rect 10318 27548 10324 27560
rect 10376 27548 10382 27600
rect 14642 27588 14648 27600
rect 14603 27560 14648 27588
rect 14642 27548 14648 27560
rect 14700 27548 14706 27600
rect 15212 27560 22094 27588
rect 3329 27523 3387 27529
rect 2924 27492 3280 27520
rect 2924 27480 2930 27492
rect 3252 27461 3280 27492
rect 3329 27489 3341 27523
rect 3375 27520 3387 27523
rect 5353 27523 5411 27529
rect 3375 27492 5304 27520
rect 3375 27489 3387 27492
rect 3329 27483 3387 27489
rect 1857 27455 1915 27461
rect 1857 27421 1869 27455
rect 1903 27421 1915 27455
rect 1857 27415 1915 27421
rect 2777 27455 2835 27461
rect 2777 27421 2789 27455
rect 2823 27452 2835 27455
rect 3237 27455 3295 27461
rect 2823 27424 2912 27452
rect 2823 27421 2835 27424
rect 2777 27415 2835 27421
rect 1872 27384 1900 27415
rect 2884 27384 2912 27424
rect 3237 27421 3249 27455
rect 3283 27421 3295 27455
rect 3237 27415 3295 27421
rect 3694 27412 3700 27464
rect 3752 27452 3758 27464
rect 4525 27455 4583 27461
rect 4525 27452 4537 27455
rect 3752 27424 4537 27452
rect 3752 27412 3758 27424
rect 4525 27421 4537 27424
rect 4571 27421 4583 27455
rect 5276 27452 5304 27492
rect 5353 27489 5365 27523
rect 5399 27489 5411 27523
rect 5353 27483 5411 27489
rect 6549 27523 6607 27529
rect 6549 27489 6561 27523
rect 6595 27520 6607 27523
rect 12069 27523 12127 27529
rect 6595 27492 11468 27520
rect 6595 27489 6607 27492
rect 6549 27483 6607 27489
rect 5534 27452 5540 27464
rect 5276 27424 5540 27452
rect 4525 27415 4583 27421
rect 5534 27412 5540 27424
rect 5592 27412 5598 27464
rect 5997 27455 6055 27461
rect 5997 27421 6009 27455
rect 6043 27452 6055 27455
rect 6454 27452 6460 27464
rect 6043 27424 6316 27452
rect 6415 27424 6460 27452
rect 6043 27421 6055 27424
rect 5997 27415 6055 27421
rect 4617 27387 4675 27393
rect 1872 27356 2774 27384
rect 2884 27356 4568 27384
rect 2746 27316 2774 27356
rect 3602 27316 3608 27328
rect 2746 27288 3608 27316
rect 3602 27276 3608 27288
rect 3660 27276 3666 27328
rect 3878 27276 3884 27328
rect 3936 27316 3942 27328
rect 3973 27319 4031 27325
rect 3973 27316 3985 27319
rect 3936 27288 3985 27316
rect 3936 27276 3942 27288
rect 3973 27285 3985 27288
rect 4019 27285 4031 27319
rect 4540 27316 4568 27356
rect 4617 27353 4629 27387
rect 4663 27384 4675 27387
rect 6086 27384 6092 27396
rect 4663 27356 6092 27384
rect 4663 27353 4675 27356
rect 4617 27347 4675 27353
rect 6086 27344 6092 27356
rect 6144 27344 6150 27396
rect 6288 27384 6316 27424
rect 6454 27412 6460 27424
rect 6512 27412 6518 27464
rect 7098 27452 7104 27464
rect 7059 27424 7104 27452
rect 7098 27412 7104 27424
rect 7156 27412 7162 27464
rect 7374 27412 7380 27464
rect 7432 27452 7438 27464
rect 7737 27455 7795 27461
rect 7737 27452 7749 27455
rect 7432 27424 7749 27452
rect 7432 27412 7438 27424
rect 7737 27421 7749 27424
rect 7783 27421 7795 27455
rect 7737 27415 7795 27421
rect 8389 27455 8447 27461
rect 8389 27421 8401 27455
rect 8435 27452 8447 27455
rect 8754 27452 8760 27464
rect 8435 27424 8760 27452
rect 8435 27421 8447 27424
rect 8389 27415 8447 27421
rect 8754 27412 8760 27424
rect 8812 27412 8818 27464
rect 9030 27412 9036 27464
rect 9088 27452 9094 27464
rect 9125 27455 9183 27461
rect 9125 27452 9137 27455
rect 9088 27424 9137 27452
rect 9088 27412 9094 27424
rect 9125 27421 9137 27424
rect 9171 27421 9183 27455
rect 9306 27452 9312 27464
rect 9267 27424 9312 27452
rect 9125 27415 9183 27421
rect 9306 27412 9312 27424
rect 9364 27412 9370 27464
rect 9398 27412 9404 27464
rect 9456 27452 9462 27464
rect 9456 27424 10364 27452
rect 9456 27412 9462 27424
rect 6914 27384 6920 27396
rect 6288 27356 6920 27384
rect 6914 27344 6920 27356
rect 6972 27344 6978 27396
rect 7837 27387 7895 27393
rect 7837 27353 7849 27387
rect 7883 27384 7895 27387
rect 7883 27356 10088 27384
rect 7883 27353 7895 27356
rect 7837 27347 7895 27353
rect 4890 27316 4896 27328
rect 4540 27288 4896 27316
rect 3973 27279 4031 27285
rect 4890 27276 4896 27288
rect 4948 27276 4954 27328
rect 5905 27319 5963 27325
rect 5905 27285 5917 27319
rect 5951 27316 5963 27319
rect 6454 27316 6460 27328
rect 5951 27288 6460 27316
rect 5951 27285 5963 27288
rect 5905 27279 5963 27285
rect 6454 27276 6460 27288
rect 6512 27276 6518 27328
rect 7193 27319 7251 27325
rect 7193 27285 7205 27319
rect 7239 27316 7251 27319
rect 7558 27316 7564 27328
rect 7239 27288 7564 27316
rect 7239 27285 7251 27288
rect 7193 27279 7251 27285
rect 7558 27276 7564 27288
rect 7616 27276 7622 27328
rect 8294 27276 8300 27328
rect 8352 27316 8358 27328
rect 9674 27316 9680 27328
rect 8352 27288 9680 27316
rect 8352 27276 8358 27288
rect 9674 27276 9680 27288
rect 9732 27276 9738 27328
rect 9766 27276 9772 27328
rect 9824 27316 9830 27328
rect 10060 27316 10088 27356
rect 10134 27344 10140 27396
rect 10192 27384 10198 27396
rect 10229 27387 10287 27393
rect 10229 27384 10241 27387
rect 10192 27356 10241 27384
rect 10192 27344 10198 27356
rect 10229 27353 10241 27356
rect 10275 27353 10287 27387
rect 10336 27384 10364 27424
rect 11149 27387 11207 27393
rect 11149 27384 11161 27387
rect 10336 27356 11161 27384
rect 10229 27347 10287 27353
rect 11149 27353 11161 27356
rect 11195 27353 11207 27387
rect 11149 27347 11207 27353
rect 11238 27344 11244 27396
rect 11296 27384 11302 27396
rect 11440 27384 11468 27492
rect 12069 27489 12081 27523
rect 12115 27520 12127 27523
rect 12434 27520 12440 27532
rect 12115 27492 12440 27520
rect 12115 27489 12127 27492
rect 12069 27483 12127 27489
rect 12434 27480 12440 27492
rect 12492 27480 12498 27532
rect 12894 27480 12900 27532
rect 12952 27520 12958 27532
rect 15212 27529 15240 27560
rect 15197 27523 15255 27529
rect 15197 27520 15209 27523
rect 12952 27492 15209 27520
rect 12952 27480 12958 27492
rect 15197 27489 15209 27492
rect 15243 27489 15255 27523
rect 15838 27520 15844 27532
rect 15799 27492 15844 27520
rect 15197 27483 15255 27489
rect 15838 27480 15844 27492
rect 15896 27480 15902 27532
rect 16482 27480 16488 27532
rect 16540 27520 16546 27532
rect 17681 27523 17739 27529
rect 16540 27492 17632 27520
rect 16540 27480 16546 27492
rect 13725 27455 13783 27461
rect 13725 27421 13737 27455
rect 13771 27452 13783 27455
rect 14550 27452 14556 27464
rect 13771 27424 14556 27452
rect 13771 27421 13783 27424
rect 13725 27415 13783 27421
rect 14550 27412 14556 27424
rect 14608 27412 14614 27464
rect 17604 27461 17632 27492
rect 17681 27489 17693 27523
rect 17727 27520 17739 27523
rect 18417 27523 18475 27529
rect 18417 27520 18429 27523
rect 17727 27492 18429 27520
rect 17727 27489 17739 27492
rect 17681 27483 17739 27489
rect 18417 27489 18429 27492
rect 18463 27489 18475 27523
rect 18417 27483 18475 27489
rect 19981 27523 20039 27529
rect 19981 27489 19993 27523
rect 20027 27520 20039 27523
rect 20070 27520 20076 27532
rect 20027 27492 20076 27520
rect 20027 27489 20039 27492
rect 19981 27483 20039 27489
rect 20070 27480 20076 27492
rect 20128 27480 20134 27532
rect 20438 27520 20444 27532
rect 20399 27492 20444 27520
rect 20438 27480 20444 27492
rect 20496 27480 20502 27532
rect 22066 27520 22094 27560
rect 24673 27523 24731 27529
rect 24673 27520 24685 27523
rect 22066 27492 24685 27520
rect 24673 27489 24685 27492
rect 24719 27489 24731 27523
rect 24673 27483 24731 27489
rect 17589 27455 17647 27461
rect 17589 27421 17601 27455
rect 17635 27421 17647 27455
rect 18230 27452 18236 27464
rect 18191 27424 18236 27452
rect 17589 27415 17647 27421
rect 12161 27387 12219 27393
rect 12161 27384 12173 27387
rect 11296 27356 11341 27384
rect 11440 27356 12173 27384
rect 11296 27344 11302 27356
rect 12161 27353 12173 27356
rect 12207 27353 12219 27387
rect 13078 27384 13084 27396
rect 12991 27356 13084 27384
rect 12161 27347 12219 27353
rect 13078 27344 13084 27356
rect 13136 27384 13142 27396
rect 15102 27384 15108 27396
rect 13136 27356 14964 27384
rect 15063 27356 15108 27384
rect 13136 27344 13142 27356
rect 11882 27316 11888 27328
rect 9824 27288 9869 27316
rect 10060 27288 11888 27316
rect 9824 27276 9830 27288
rect 11882 27276 11888 27288
rect 11940 27276 11946 27328
rect 12986 27276 12992 27328
rect 13044 27316 13050 27328
rect 13541 27319 13599 27325
rect 13541 27316 13553 27319
rect 13044 27288 13553 27316
rect 13044 27276 13050 27288
rect 13541 27285 13553 27288
rect 13587 27285 13599 27319
rect 14936 27316 14964 27356
rect 15102 27344 15108 27356
rect 15160 27344 15166 27396
rect 15933 27387 15991 27393
rect 15933 27353 15945 27387
rect 15979 27384 15991 27387
rect 16666 27384 16672 27396
rect 15979 27356 16672 27384
rect 15979 27353 15991 27356
rect 15933 27347 15991 27353
rect 16666 27344 16672 27356
rect 16724 27344 16730 27396
rect 16850 27384 16856 27396
rect 16811 27356 16856 27384
rect 16850 27344 16856 27356
rect 16908 27344 16914 27396
rect 17604 27384 17632 27415
rect 18230 27412 18236 27424
rect 18288 27412 18294 27464
rect 21269 27455 21327 27461
rect 21269 27452 21281 27455
rect 20640 27424 21281 27452
rect 17678 27384 17684 27396
rect 17604 27356 17684 27384
rect 17678 27344 17684 27356
rect 17736 27344 17742 27396
rect 20073 27387 20131 27393
rect 20073 27353 20085 27387
rect 20119 27384 20131 27387
rect 20346 27384 20352 27396
rect 20119 27356 20352 27384
rect 20119 27353 20131 27356
rect 20073 27347 20131 27353
rect 20346 27344 20352 27356
rect 20404 27344 20410 27396
rect 16868 27316 16896 27344
rect 14936 27288 16896 27316
rect 13541 27279 13599 27285
rect 16942 27276 16948 27328
rect 17000 27316 17006 27328
rect 20640 27316 20668 27424
rect 21269 27421 21281 27424
rect 21315 27452 21327 27455
rect 21729 27455 21787 27461
rect 21729 27452 21741 27455
rect 21315 27424 21741 27452
rect 21315 27421 21327 27424
rect 21269 27415 21327 27421
rect 21729 27421 21741 27424
rect 21775 27452 21787 27455
rect 24765 27455 24823 27461
rect 21775 27424 22094 27452
rect 21775 27421 21787 27424
rect 21729 27415 21787 27421
rect 21174 27316 21180 27328
rect 17000 27288 20668 27316
rect 21135 27288 21180 27316
rect 17000 27276 17006 27288
rect 21174 27276 21180 27288
rect 21232 27276 21238 27328
rect 22066 27316 22094 27424
rect 24765 27421 24777 27455
rect 24811 27452 24823 27455
rect 24811 27424 25360 27452
rect 24811 27421 24823 27424
rect 24765 27415 24823 27421
rect 25332 27393 25360 27424
rect 25317 27387 25375 27393
rect 25317 27353 25329 27387
rect 25363 27384 25375 27387
rect 34146 27384 34152 27396
rect 25363 27356 34152 27384
rect 25363 27353 25375 27356
rect 25317 27347 25375 27353
rect 34146 27344 34152 27356
rect 34204 27384 34210 27396
rect 34790 27384 34796 27396
rect 34204 27356 34796 27384
rect 34204 27344 34210 27356
rect 34790 27344 34796 27356
rect 34848 27344 34854 27396
rect 37918 27316 37924 27328
rect 22066 27288 37924 27316
rect 37918 27276 37924 27288
rect 37976 27276 37982 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 2409 27115 2467 27121
rect 2409 27081 2421 27115
rect 2455 27112 2467 27115
rect 2498 27112 2504 27124
rect 2455 27084 2504 27112
rect 2455 27081 2467 27084
rect 2409 27075 2467 27081
rect 2498 27072 2504 27084
rect 2556 27072 2562 27124
rect 3050 27112 3056 27124
rect 3011 27084 3056 27112
rect 3050 27072 3056 27084
rect 3108 27072 3114 27124
rect 3878 27072 3884 27124
rect 3936 27112 3942 27124
rect 5442 27112 5448 27124
rect 3936 27084 5448 27112
rect 3936 27072 3942 27084
rect 3973 27047 4031 27053
rect 3973 27013 3985 27047
rect 4019 27044 4031 27047
rect 4890 27044 4896 27056
rect 4019 27016 4896 27044
rect 4019 27013 4031 27016
rect 3973 27007 4031 27013
rect 4890 27004 4896 27016
rect 4948 27004 4954 27056
rect 1762 26936 1768 26988
rect 1820 26976 1826 26988
rect 1857 26979 1915 26985
rect 1857 26976 1869 26979
rect 1820 26948 1869 26976
rect 1820 26936 1826 26948
rect 1857 26945 1869 26948
rect 1903 26945 1915 26979
rect 2498 26976 2504 26988
rect 2459 26948 2504 26976
rect 1857 26939 1915 26945
rect 2498 26936 2504 26948
rect 2556 26936 2562 26988
rect 2958 26976 2964 26988
rect 2746 26948 2964 26976
rect 2314 26868 2320 26920
rect 2372 26908 2378 26920
rect 2746 26908 2774 26948
rect 2958 26936 2964 26948
rect 3016 26936 3022 26988
rect 3234 26936 3240 26988
rect 3292 26976 3298 26988
rect 3881 26979 3939 26985
rect 3881 26976 3893 26979
rect 3292 26948 3893 26976
rect 3292 26936 3298 26948
rect 3881 26945 3893 26948
rect 3927 26945 3939 26979
rect 3881 26939 3939 26945
rect 4525 26979 4583 26985
rect 4525 26945 4537 26979
rect 4571 26976 4583 26979
rect 5074 26976 5080 26988
rect 4571 26948 5080 26976
rect 4571 26945 4583 26948
rect 4525 26939 4583 26945
rect 5074 26936 5080 26948
rect 5132 26936 5138 26988
rect 5169 26979 5227 26985
rect 5169 26945 5181 26979
rect 5215 26976 5227 26979
rect 5276 26976 5304 27084
rect 5442 27072 5448 27084
rect 5500 27112 5506 27124
rect 5500 27084 6040 27112
rect 5500 27072 5506 27084
rect 5215 26948 5304 26976
rect 5215 26945 5227 26948
rect 5169 26939 5227 26945
rect 5818 26942 5824 26994
rect 5876 26982 5882 26994
rect 5876 26954 5921 26982
rect 6012 26976 6040 27084
rect 6178 27072 6184 27124
rect 6236 27112 6242 27124
rect 8202 27112 8208 27124
rect 6236 27084 8208 27112
rect 6236 27072 6242 27084
rect 8202 27072 8208 27084
rect 8260 27072 8266 27124
rect 9306 27072 9312 27124
rect 9364 27112 9370 27124
rect 11054 27112 11060 27124
rect 9364 27084 11060 27112
rect 9364 27072 9370 27084
rect 11054 27072 11060 27084
rect 11112 27072 11118 27124
rect 11238 27072 11244 27124
rect 11296 27112 11302 27124
rect 16114 27112 16120 27124
rect 11296 27084 16120 27112
rect 11296 27072 11302 27084
rect 16114 27072 16120 27084
rect 16172 27072 16178 27124
rect 16209 27115 16267 27121
rect 16209 27081 16221 27115
rect 16255 27112 16267 27115
rect 16574 27112 16580 27124
rect 16255 27084 16580 27112
rect 16255 27081 16267 27084
rect 16209 27075 16267 27081
rect 16574 27072 16580 27084
rect 16632 27072 16638 27124
rect 18230 27072 18236 27124
rect 18288 27112 18294 27124
rect 20346 27112 20352 27124
rect 18288 27084 19840 27112
rect 20307 27084 20352 27112
rect 18288 27072 18294 27084
rect 7834 27004 7840 27056
rect 7892 27044 7898 27056
rect 8021 27047 8079 27053
rect 8021 27044 8033 27047
rect 7892 27016 8033 27044
rect 7892 27004 7898 27016
rect 8021 27013 8033 27016
rect 8067 27013 8079 27047
rect 8021 27007 8079 27013
rect 8113 27047 8171 27053
rect 8113 27013 8125 27047
rect 8159 27044 8171 27047
rect 9122 27044 9128 27056
rect 8159 27016 9128 27044
rect 8159 27013 8171 27016
rect 8113 27007 8171 27013
rect 9122 27004 9128 27016
rect 9180 27004 9186 27056
rect 9214 27004 9220 27056
rect 9272 27044 9278 27056
rect 10413 27047 10471 27053
rect 10413 27044 10425 27047
rect 9272 27016 9317 27044
rect 9784 27016 10425 27044
rect 9272 27004 9278 27016
rect 6825 26979 6883 26985
rect 6825 26976 6837 26979
rect 5876 26942 5882 26954
rect 6012 26948 6837 26976
rect 6825 26945 6837 26948
rect 6871 26945 6883 26979
rect 6825 26939 6883 26945
rect 7374 26936 7380 26988
rect 7432 26976 7438 26988
rect 7469 26979 7527 26985
rect 7469 26976 7481 26979
rect 7432 26948 7481 26976
rect 7432 26936 7438 26948
rect 7469 26945 7481 26948
rect 7515 26945 7527 26979
rect 7469 26939 7527 26945
rect 2372 26880 2774 26908
rect 4617 26911 4675 26917
rect 2372 26868 2378 26880
rect 4617 26877 4629 26911
rect 4663 26908 4675 26911
rect 8018 26908 8024 26920
rect 4663 26880 8024 26908
rect 4663 26877 4675 26880
rect 4617 26871 4675 26877
rect 8018 26868 8024 26880
rect 8076 26868 8082 26920
rect 9122 26908 9128 26920
rect 9083 26880 9128 26908
rect 9122 26868 9128 26880
rect 9180 26868 9186 26920
rect 5905 26843 5963 26849
rect 5905 26809 5917 26843
rect 5951 26840 5963 26843
rect 9030 26840 9036 26852
rect 5951 26812 9036 26840
rect 5951 26809 5963 26812
rect 5905 26803 5963 26809
rect 9030 26800 9036 26812
rect 9088 26800 9094 26852
rect 9674 26840 9680 26852
rect 9635 26812 9680 26840
rect 9674 26800 9680 26812
rect 9732 26800 9738 26852
rect 1670 26772 1676 26784
rect 1631 26744 1676 26772
rect 1670 26732 1676 26744
rect 1728 26732 1734 26784
rect 3050 26732 3056 26784
rect 3108 26772 3114 26784
rect 4890 26772 4896 26784
rect 3108 26744 4896 26772
rect 3108 26732 3114 26744
rect 4890 26732 4896 26744
rect 4948 26732 4954 26784
rect 5261 26775 5319 26781
rect 5261 26741 5273 26775
rect 5307 26772 5319 26775
rect 6178 26772 6184 26784
rect 5307 26744 6184 26772
rect 5307 26741 5319 26744
rect 5261 26735 5319 26741
rect 6178 26732 6184 26744
rect 6236 26732 6242 26784
rect 6917 26775 6975 26781
rect 6917 26741 6929 26775
rect 6963 26772 6975 26775
rect 9784 26772 9812 27016
rect 10413 27013 10425 27016
rect 10459 27013 10471 27047
rect 10413 27007 10471 27013
rect 10594 27004 10600 27056
rect 10652 27044 10658 27056
rect 10962 27044 10968 27056
rect 10652 27016 10968 27044
rect 10652 27004 10658 27016
rect 10962 27004 10968 27016
rect 11020 27004 11026 27056
rect 11882 27044 11888 27056
rect 11843 27016 11888 27044
rect 11882 27004 11888 27016
rect 11940 27004 11946 27056
rect 12805 27047 12863 27053
rect 12805 27013 12817 27047
rect 12851 27044 12863 27047
rect 13078 27044 13084 27056
rect 12851 27016 13084 27044
rect 12851 27013 12863 27016
rect 12805 27007 12863 27013
rect 13078 27004 13084 27016
rect 13136 27004 13142 27056
rect 14366 27044 14372 27056
rect 14327 27016 14372 27044
rect 14366 27004 14372 27016
rect 14424 27004 14430 27056
rect 14918 27044 14924 27056
rect 14879 27016 14924 27044
rect 14918 27004 14924 27016
rect 14976 27004 14982 27056
rect 15102 27004 15108 27056
rect 15160 27044 15166 27056
rect 16945 27047 17003 27053
rect 16945 27044 16957 27047
rect 15160 27016 16957 27044
rect 15160 27004 15166 27016
rect 16945 27013 16957 27016
rect 16991 27013 17003 27047
rect 16945 27007 17003 27013
rect 17037 27047 17095 27053
rect 17037 27013 17049 27047
rect 17083 27044 17095 27047
rect 17954 27044 17960 27056
rect 17083 27016 17960 27044
rect 17083 27013 17095 27016
rect 17037 27007 17095 27013
rect 17954 27004 17960 27016
rect 18012 27004 18018 27056
rect 18325 27047 18383 27053
rect 18325 27013 18337 27047
rect 18371 27044 18383 27047
rect 19334 27044 19340 27056
rect 18371 27016 19340 27044
rect 18371 27013 18383 27016
rect 18325 27007 18383 27013
rect 19334 27004 19340 27016
rect 19392 27004 19398 27056
rect 19429 27047 19487 27053
rect 19429 27013 19441 27047
rect 19475 27044 19487 27047
rect 19518 27044 19524 27056
rect 19475 27016 19524 27044
rect 19475 27013 19487 27016
rect 19429 27007 19487 27013
rect 19518 27004 19524 27016
rect 19576 27004 19582 27056
rect 19812 27044 19840 27084
rect 20346 27072 20352 27084
rect 20404 27072 20410 27124
rect 22097 27115 22155 27121
rect 22097 27081 22109 27115
rect 22143 27112 22155 27115
rect 22646 27112 22652 27124
rect 22143 27084 22652 27112
rect 22143 27081 22155 27084
rect 22097 27075 22155 27081
rect 21174 27044 21180 27056
rect 19812 27016 21180 27044
rect 13446 26936 13452 26988
rect 13504 26976 13510 26988
rect 13725 26979 13783 26985
rect 13725 26976 13737 26979
rect 13504 26948 13737 26976
rect 13504 26936 13510 26948
rect 13725 26945 13737 26948
rect 13771 26945 13783 26979
rect 13725 26939 13783 26945
rect 15565 26979 15623 26985
rect 15565 26945 15577 26979
rect 15611 26945 15623 26979
rect 16114 26976 16120 26988
rect 16075 26948 16120 26976
rect 15565 26939 15623 26945
rect 10318 26908 10324 26920
rect 10279 26880 10324 26908
rect 10318 26868 10324 26880
rect 10376 26868 10382 26920
rect 11793 26911 11851 26917
rect 11793 26908 11805 26911
rect 10704 26880 11805 26908
rect 9858 26800 9864 26852
rect 9916 26840 9922 26852
rect 10704 26840 10732 26880
rect 11793 26877 11805 26880
rect 11839 26877 11851 26911
rect 11793 26871 11851 26877
rect 12250 26868 12256 26920
rect 12308 26908 12314 26920
rect 12308 26880 13860 26908
rect 12308 26868 12314 26880
rect 9916 26812 10732 26840
rect 13832 26840 13860 26880
rect 14090 26868 14096 26920
rect 14148 26908 14154 26920
rect 14277 26911 14335 26917
rect 14277 26908 14289 26911
rect 14148 26880 14289 26908
rect 14148 26868 14154 26880
rect 14277 26877 14289 26880
rect 14323 26877 14335 26911
rect 14277 26871 14335 26877
rect 15580 26840 15608 26939
rect 16114 26936 16120 26948
rect 16172 26936 16178 26988
rect 17678 26936 17684 26988
rect 17736 26976 17742 26988
rect 18233 26979 18291 26985
rect 18233 26976 18245 26979
rect 17736 26948 18245 26976
rect 17736 26936 17742 26948
rect 18233 26945 18245 26948
rect 18279 26976 18291 26979
rect 18598 26976 18604 26988
rect 18279 26948 18604 26976
rect 18279 26945 18291 26948
rect 18233 26939 18291 26945
rect 18598 26936 18604 26948
rect 18656 26936 18662 26988
rect 17218 26868 17224 26920
rect 17276 26908 17282 26920
rect 18877 26911 18935 26917
rect 18877 26908 18889 26911
rect 17276 26880 18184 26908
rect 17276 26868 17282 26880
rect 13832 26812 15608 26840
rect 17497 26843 17555 26849
rect 9916 26800 9922 26812
rect 17497 26809 17509 26843
rect 17543 26840 17555 26843
rect 17862 26840 17868 26852
rect 17543 26812 17868 26840
rect 17543 26809 17555 26812
rect 17497 26803 17555 26809
rect 17862 26800 17868 26812
rect 17920 26800 17926 26852
rect 18156 26840 18184 26880
rect 18524 26880 18889 26908
rect 18524 26840 18552 26880
rect 18877 26877 18889 26880
rect 18923 26908 18935 26911
rect 19334 26908 19340 26920
rect 18923 26880 19340 26908
rect 18923 26877 18935 26880
rect 18877 26871 18935 26877
rect 19334 26868 19340 26880
rect 19392 26868 19398 26920
rect 19521 26911 19579 26917
rect 19521 26877 19533 26911
rect 19567 26908 19579 26911
rect 19812 26908 19840 27016
rect 21174 27004 21180 27016
rect 21232 27004 21238 27056
rect 20441 26979 20499 26985
rect 20441 26945 20453 26979
rect 20487 26976 20499 26979
rect 20714 26976 20720 26988
rect 20487 26948 20720 26976
rect 20487 26945 20499 26948
rect 20441 26939 20499 26945
rect 20714 26936 20720 26948
rect 20772 26976 20778 26988
rect 20901 26979 20959 26985
rect 20901 26976 20913 26979
rect 20772 26948 20913 26976
rect 20772 26936 20778 26948
rect 20901 26945 20913 26948
rect 20947 26976 20959 26979
rect 21634 26976 21640 26988
rect 20947 26948 21640 26976
rect 20947 26945 20959 26948
rect 20901 26939 20959 26945
rect 21634 26936 21640 26948
rect 21692 26936 21698 26988
rect 19567 26880 19840 26908
rect 19567 26877 19579 26880
rect 19521 26871 19579 26877
rect 18156 26812 18552 26840
rect 18598 26800 18604 26852
rect 18656 26840 18662 26852
rect 22112 26840 22140 27075
rect 22646 27072 22652 27084
rect 22704 27072 22710 27124
rect 23753 27115 23811 27121
rect 23753 27081 23765 27115
rect 23799 27112 23811 27115
rect 25314 27112 25320 27124
rect 23799 27084 25320 27112
rect 23799 27081 23811 27084
rect 23753 27075 23811 27081
rect 25314 27072 25320 27084
rect 25372 27072 25378 27124
rect 22278 27004 22284 27056
rect 22336 27044 22342 27056
rect 22557 27047 22615 27053
rect 22557 27044 22569 27047
rect 22336 27016 22569 27044
rect 22336 27004 22342 27016
rect 22557 27013 22569 27016
rect 22603 27013 22615 27047
rect 22557 27007 22615 27013
rect 37734 27004 37740 27056
rect 37792 27044 37798 27056
rect 38013 27047 38071 27053
rect 38013 27044 38025 27047
rect 37792 27016 38025 27044
rect 37792 27004 37798 27016
rect 38013 27013 38025 27016
rect 38059 27013 38071 27047
rect 38013 27007 38071 27013
rect 23566 26976 23572 26988
rect 23527 26948 23572 26976
rect 23566 26936 23572 26948
rect 23624 26976 23630 26988
rect 24213 26979 24271 26985
rect 24213 26976 24225 26979
rect 23624 26948 24225 26976
rect 23624 26936 23630 26948
rect 24213 26945 24225 26948
rect 24259 26976 24271 26979
rect 37553 26979 37611 26985
rect 24259 26948 26234 26976
rect 24259 26945 24271 26948
rect 24213 26939 24271 26945
rect 18656 26812 22140 26840
rect 26206 26840 26234 26948
rect 37553 26945 37565 26979
rect 37599 26976 37611 26979
rect 38194 26976 38200 26988
rect 37599 26948 38200 26976
rect 37599 26945 37611 26948
rect 37553 26939 37611 26945
rect 38194 26936 38200 26948
rect 38252 26936 38258 26988
rect 38286 26840 38292 26852
rect 26206 26812 38292 26840
rect 18656 26800 18662 26812
rect 38286 26800 38292 26812
rect 38344 26800 38350 26852
rect 6963 26744 9812 26772
rect 6963 26741 6975 26744
rect 6917 26735 6975 26741
rect 10318 26732 10324 26784
rect 10376 26772 10382 26784
rect 12802 26772 12808 26784
rect 10376 26744 12808 26772
rect 10376 26732 10382 26744
rect 12802 26732 12808 26744
rect 12860 26732 12866 26784
rect 13630 26772 13636 26784
rect 13591 26744 13636 26772
rect 13630 26732 13636 26744
rect 13688 26732 13694 26784
rect 15378 26732 15384 26784
rect 15436 26772 15442 26784
rect 15473 26775 15531 26781
rect 15473 26772 15485 26775
rect 15436 26744 15485 26772
rect 15436 26732 15442 26744
rect 15473 26741 15485 26744
rect 15519 26741 15531 26775
rect 15473 26735 15531 26741
rect 16114 26732 16120 26784
rect 16172 26772 16178 26784
rect 22278 26772 22284 26784
rect 16172 26744 22284 26772
rect 16172 26732 16178 26744
rect 22278 26732 22284 26744
rect 22336 26732 22342 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 1949 26571 2007 26577
rect 1949 26537 1961 26571
rect 1995 26568 2007 26571
rect 2130 26568 2136 26580
rect 1995 26540 2136 26568
rect 1995 26537 2007 26540
rect 1949 26531 2007 26537
rect 2130 26528 2136 26540
rect 2188 26528 2194 26580
rect 2406 26528 2412 26580
rect 2464 26568 2470 26580
rect 2464 26540 4660 26568
rect 2464 26528 2470 26540
rect 1302 26460 1308 26512
rect 1360 26500 1366 26512
rect 2593 26503 2651 26509
rect 2593 26500 2605 26503
rect 1360 26472 2605 26500
rect 1360 26460 1366 26472
rect 2593 26469 2605 26472
rect 2639 26469 2651 26503
rect 2593 26463 2651 26469
rect 842 26392 848 26444
rect 900 26432 906 26444
rect 3050 26432 3056 26444
rect 900 26404 3056 26432
rect 900 26392 906 26404
rect 3050 26392 3056 26404
rect 3108 26392 3114 26444
rect 3142 26392 3148 26444
rect 3200 26432 3206 26444
rect 3878 26432 3884 26444
rect 3200 26404 3884 26432
rect 3200 26392 3206 26404
rect 3878 26392 3884 26404
rect 3936 26432 3942 26444
rect 3936 26404 4016 26432
rect 3936 26392 3942 26404
rect 1857 26367 1915 26373
rect 1857 26333 1869 26367
rect 1903 26364 1915 26367
rect 2314 26364 2320 26376
rect 1903 26336 2320 26364
rect 1903 26333 1915 26336
rect 1857 26327 1915 26333
rect 2314 26324 2320 26336
rect 2372 26324 2378 26376
rect 2501 26367 2559 26373
rect 2501 26333 2513 26367
rect 2547 26333 2559 26367
rect 2501 26327 2559 26333
rect 1946 26256 1952 26308
rect 2004 26296 2010 26308
rect 2130 26296 2136 26308
rect 2004 26268 2136 26296
rect 2004 26256 2010 26268
rect 2130 26256 2136 26268
rect 2188 26256 2194 26308
rect 2406 26188 2412 26240
rect 2464 26228 2470 26240
rect 2516 26228 2544 26327
rect 2774 26324 2780 26376
rect 2832 26364 2838 26376
rect 3237 26367 3295 26373
rect 3237 26364 3249 26367
rect 2832 26336 3249 26364
rect 2832 26324 2838 26336
rect 3237 26333 3249 26336
rect 3283 26364 3295 26367
rect 3602 26364 3608 26376
rect 3283 26336 3608 26364
rect 3283 26333 3295 26336
rect 3237 26327 3295 26333
rect 3602 26324 3608 26336
rect 3660 26324 3666 26376
rect 3988 26373 4016 26404
rect 3973 26367 4031 26373
rect 3973 26333 3985 26367
rect 4019 26333 4031 26367
rect 3973 26327 4031 26333
rect 4065 26367 4123 26373
rect 4065 26333 4077 26367
rect 4111 26364 4123 26367
rect 4522 26364 4528 26376
rect 4111 26336 4528 26364
rect 4111 26333 4123 26336
rect 4065 26327 4123 26333
rect 4522 26324 4528 26336
rect 4580 26324 4586 26376
rect 4632 26373 4660 26540
rect 5074 26528 5080 26580
rect 5132 26568 5138 26580
rect 7006 26568 7012 26580
rect 5132 26540 7012 26568
rect 5132 26528 5138 26540
rect 7006 26528 7012 26540
rect 7064 26528 7070 26580
rect 7374 26528 7380 26580
rect 7432 26568 7438 26580
rect 7558 26568 7564 26580
rect 7432 26540 7564 26568
rect 7432 26528 7438 26540
rect 7558 26528 7564 26540
rect 7616 26528 7622 26580
rect 7650 26528 7656 26580
rect 7708 26568 7714 26580
rect 9493 26571 9551 26577
rect 9493 26568 9505 26571
rect 7708 26540 9505 26568
rect 7708 26528 7714 26540
rect 9493 26537 9505 26540
rect 9539 26568 9551 26571
rect 9766 26568 9772 26580
rect 9539 26540 9772 26568
rect 9539 26537 9551 26540
rect 9493 26531 9551 26537
rect 9766 26528 9772 26540
rect 9824 26528 9830 26580
rect 10042 26528 10048 26580
rect 10100 26568 10106 26580
rect 11882 26568 11888 26580
rect 10100 26540 11888 26568
rect 10100 26528 10106 26540
rect 11882 26528 11888 26540
rect 11940 26528 11946 26580
rect 12434 26568 12440 26580
rect 12084 26540 12440 26568
rect 12084 26509 12112 26540
rect 12434 26528 12440 26540
rect 12492 26568 12498 26580
rect 13722 26568 13728 26580
rect 12492 26540 13728 26568
rect 12492 26528 12498 26540
rect 13722 26528 13728 26540
rect 13780 26528 13786 26580
rect 15102 26568 15108 26580
rect 15063 26540 15108 26568
rect 15102 26528 15108 26540
rect 15160 26528 15166 26580
rect 17126 26568 17132 26580
rect 17087 26540 17132 26568
rect 17126 26528 17132 26540
rect 17184 26528 17190 26580
rect 17218 26528 17224 26580
rect 17276 26568 17282 26580
rect 18690 26568 18696 26580
rect 17276 26540 18696 26568
rect 17276 26528 17282 26540
rect 18690 26528 18696 26540
rect 18748 26528 18754 26580
rect 18874 26568 18880 26580
rect 18835 26540 18880 26568
rect 18874 26528 18880 26540
rect 18932 26568 18938 26580
rect 19521 26571 19579 26577
rect 19521 26568 19533 26571
rect 18932 26540 19533 26568
rect 18932 26528 18938 26540
rect 19521 26537 19533 26540
rect 19567 26537 19579 26571
rect 19521 26531 19579 26537
rect 19610 26528 19616 26580
rect 19668 26568 19674 26580
rect 20530 26568 20536 26580
rect 19668 26540 20536 26568
rect 19668 26528 19674 26540
rect 20530 26528 20536 26540
rect 20588 26528 20594 26580
rect 20714 26528 20720 26580
rect 20772 26568 20778 26580
rect 20809 26571 20867 26577
rect 20809 26568 20821 26571
rect 20772 26540 20821 26568
rect 20772 26528 20778 26540
rect 20809 26537 20821 26540
rect 20855 26537 20867 26571
rect 20809 26531 20867 26537
rect 7285 26503 7343 26509
rect 7285 26469 7297 26503
rect 7331 26500 7343 26503
rect 11241 26503 11299 26509
rect 7331 26472 11192 26500
rect 7331 26469 7343 26472
rect 7285 26463 7343 26469
rect 4709 26435 4767 26441
rect 4709 26401 4721 26435
rect 4755 26432 4767 26435
rect 4755 26404 8616 26432
rect 4755 26401 4767 26404
rect 4709 26395 4767 26401
rect 4617 26367 4675 26373
rect 4617 26333 4629 26367
rect 4663 26333 4675 26367
rect 4617 26327 4675 26333
rect 4890 26324 4896 26376
rect 4948 26364 4954 26376
rect 5261 26367 5319 26373
rect 5261 26364 5273 26367
rect 4948 26336 5273 26364
rect 4948 26324 4954 26336
rect 5261 26333 5273 26336
rect 5307 26333 5319 26367
rect 5261 26327 5319 26333
rect 5626 26324 5632 26376
rect 5684 26364 5690 26376
rect 5905 26367 5963 26373
rect 5905 26364 5917 26367
rect 5684 26336 5917 26364
rect 5684 26324 5690 26336
rect 5905 26333 5917 26336
rect 5951 26333 5963 26367
rect 6638 26364 6644 26376
rect 6599 26336 6644 26364
rect 5905 26327 5963 26333
rect 6638 26324 6644 26336
rect 6696 26324 6702 26376
rect 6733 26367 6791 26373
rect 6733 26333 6745 26367
rect 6779 26333 6791 26367
rect 6733 26327 6791 26333
rect 3329 26299 3387 26305
rect 3329 26265 3341 26299
rect 3375 26296 3387 26299
rect 4798 26296 4804 26308
rect 3375 26268 4804 26296
rect 3375 26265 3387 26268
rect 3329 26259 3387 26265
rect 4798 26256 4804 26268
rect 4856 26256 4862 26308
rect 5353 26299 5411 26305
rect 5353 26265 5365 26299
rect 5399 26296 5411 26299
rect 5997 26299 6055 26305
rect 5399 26268 5948 26296
rect 5399 26265 5411 26268
rect 5353 26259 5411 26265
rect 2464 26200 2544 26228
rect 2464 26188 2470 26200
rect 3142 26188 3148 26240
rect 3200 26228 3206 26240
rect 5074 26228 5080 26240
rect 3200 26200 5080 26228
rect 3200 26188 3206 26200
rect 5074 26188 5080 26200
rect 5132 26188 5138 26240
rect 5920 26228 5948 26268
rect 5997 26265 6009 26299
rect 6043 26296 6055 26299
rect 6454 26296 6460 26308
rect 6043 26268 6460 26296
rect 6043 26265 6055 26268
rect 5997 26259 6055 26265
rect 6454 26256 6460 26268
rect 6512 26256 6518 26308
rect 6748 26296 6776 26327
rect 7006 26324 7012 26376
rect 7064 26364 7070 26376
rect 7193 26367 7251 26373
rect 7193 26364 7205 26367
rect 7064 26336 7205 26364
rect 7064 26324 7070 26336
rect 7193 26333 7205 26336
rect 7239 26364 7251 26367
rect 7282 26364 7288 26376
rect 7239 26336 7288 26364
rect 7239 26333 7251 26336
rect 7193 26327 7251 26333
rect 7282 26324 7288 26336
rect 7340 26324 7346 26376
rect 8588 26364 8616 26404
rect 9030 26392 9036 26444
rect 9088 26432 9094 26444
rect 10137 26435 10195 26441
rect 9088 26404 10088 26432
rect 9088 26392 9094 26404
rect 9398 26364 9404 26376
rect 8588 26336 9404 26364
rect 9398 26324 9404 26336
rect 9456 26324 9462 26376
rect 9950 26364 9956 26376
rect 9911 26336 9956 26364
rect 9950 26324 9956 26336
rect 10008 26324 10014 26376
rect 10060 26364 10088 26404
rect 10137 26401 10149 26435
rect 10183 26432 10195 26435
rect 10318 26432 10324 26444
rect 10183 26404 10324 26432
rect 10183 26401 10195 26404
rect 10137 26395 10195 26401
rect 10318 26392 10324 26404
rect 10376 26392 10382 26444
rect 10778 26432 10784 26444
rect 10739 26404 10784 26432
rect 10778 26392 10784 26404
rect 10836 26392 10842 26444
rect 11164 26432 11192 26472
rect 11241 26469 11253 26503
rect 11287 26500 11299 26503
rect 12069 26503 12127 26509
rect 12069 26500 12081 26503
rect 11287 26472 12081 26500
rect 11287 26469 11299 26472
rect 11241 26463 11299 26469
rect 12069 26469 12081 26472
rect 12115 26469 12127 26503
rect 13078 26500 13084 26512
rect 12069 26463 12127 26469
rect 12176 26472 13084 26500
rect 12176 26432 12204 26472
rect 13078 26460 13084 26472
rect 13136 26460 13142 26512
rect 16390 26500 16396 26512
rect 15488 26472 16396 26500
rect 13725 26435 13783 26441
rect 11164 26404 12204 26432
rect 12406 26404 12848 26432
rect 10597 26367 10655 26373
rect 10597 26364 10609 26367
rect 10060 26336 10609 26364
rect 10597 26333 10609 26336
rect 10643 26333 10655 26367
rect 10597 26327 10655 26333
rect 11514 26324 11520 26376
rect 11572 26364 11578 26376
rect 11701 26367 11759 26373
rect 11701 26364 11713 26367
rect 11572 26336 11713 26364
rect 11572 26324 11578 26336
rect 11701 26333 11713 26336
rect 11747 26333 11759 26367
rect 11882 26364 11888 26376
rect 11843 26336 11888 26364
rect 11701 26327 11759 26333
rect 11882 26324 11888 26336
rect 11940 26324 11946 26376
rect 7650 26296 7656 26308
rect 6748 26268 7656 26296
rect 7650 26256 7656 26268
rect 7708 26256 7714 26308
rect 7926 26296 7932 26308
rect 7887 26268 7932 26296
rect 7926 26256 7932 26268
rect 7984 26256 7990 26308
rect 8018 26256 8024 26308
rect 8076 26296 8082 26308
rect 8076 26268 8121 26296
rect 8076 26256 8082 26268
rect 8294 26256 8300 26308
rect 8352 26296 8358 26308
rect 8573 26299 8631 26305
rect 8573 26296 8585 26299
rect 8352 26268 8585 26296
rect 8352 26256 8358 26268
rect 8573 26265 8585 26268
rect 8619 26265 8631 26299
rect 8573 26259 8631 26265
rect 8754 26256 8760 26308
rect 8812 26296 8818 26308
rect 9306 26296 9312 26308
rect 8812 26268 9312 26296
rect 8812 26256 8818 26268
rect 9306 26256 9312 26268
rect 9364 26256 9370 26308
rect 9674 26256 9680 26308
rect 9732 26296 9738 26308
rect 12406 26296 12434 26404
rect 9732 26268 12434 26296
rect 9732 26256 9738 26268
rect 9214 26228 9220 26240
rect 5920 26200 9220 26228
rect 9214 26188 9220 26200
rect 9272 26188 9278 26240
rect 9490 26188 9496 26240
rect 9548 26228 9554 26240
rect 12710 26228 12716 26240
rect 9548 26200 12716 26228
rect 9548 26188 9554 26200
rect 12710 26188 12716 26200
rect 12768 26188 12774 26240
rect 12820 26228 12848 26404
rect 13725 26401 13737 26435
rect 13771 26432 13783 26435
rect 14918 26432 14924 26444
rect 13771 26404 14924 26432
rect 13771 26401 13783 26404
rect 13725 26395 13783 26401
rect 14918 26392 14924 26404
rect 14976 26392 14982 26444
rect 15289 26435 15347 26441
rect 15289 26401 15301 26435
rect 15335 26432 15347 26435
rect 15378 26432 15384 26444
rect 15335 26404 15384 26432
rect 15335 26401 15347 26404
rect 15289 26395 15347 26401
rect 15378 26392 15384 26404
rect 15436 26392 15442 26444
rect 15488 26441 15516 26472
rect 16390 26460 16396 26472
rect 16448 26500 16454 26512
rect 16448 26472 22094 26500
rect 16448 26460 16454 26472
rect 15473 26435 15531 26441
rect 15473 26401 15485 26435
rect 15519 26401 15531 26435
rect 15473 26395 15531 26401
rect 16040 26404 16988 26432
rect 12894 26324 12900 26376
rect 12952 26324 12958 26376
rect 14369 26367 14427 26373
rect 14369 26333 14381 26367
rect 14415 26364 14427 26367
rect 16040 26364 16068 26404
rect 16960 26376 16988 26404
rect 18138 26392 18144 26444
rect 18196 26432 18202 26444
rect 18233 26435 18291 26441
rect 18233 26432 18245 26435
rect 18196 26404 18245 26432
rect 18196 26392 18202 26404
rect 18233 26401 18245 26404
rect 18279 26401 18291 26435
rect 18233 26395 18291 26401
rect 18322 26392 18328 26444
rect 18380 26432 18386 26444
rect 19981 26435 20039 26441
rect 19981 26432 19993 26435
rect 18380 26404 19993 26432
rect 18380 26392 18386 26404
rect 19981 26401 19993 26404
rect 20027 26401 20039 26435
rect 21913 26435 21971 26441
rect 21913 26432 21925 26435
rect 19981 26395 20039 26401
rect 20088 26404 21925 26432
rect 14415 26336 16068 26364
rect 16117 26367 16175 26373
rect 14415 26333 14427 26336
rect 14369 26327 14427 26333
rect 16117 26333 16129 26367
rect 16163 26333 16175 26367
rect 16942 26364 16948 26376
rect 16903 26336 16948 26364
rect 16117 26327 16175 26333
rect 12912 26296 12940 26324
rect 13081 26299 13139 26305
rect 13081 26296 13093 26299
rect 12912 26268 13093 26296
rect 13081 26265 13093 26268
rect 13127 26265 13139 26299
rect 13081 26259 13139 26265
rect 13173 26299 13231 26305
rect 13173 26265 13185 26299
rect 13219 26265 13231 26299
rect 13173 26259 13231 26265
rect 13188 26228 13216 26259
rect 14550 26256 14556 26308
rect 14608 26296 14614 26308
rect 16025 26299 16083 26305
rect 16025 26296 16037 26299
rect 14608 26268 16037 26296
rect 14608 26256 14614 26268
rect 16025 26265 16037 26268
rect 16071 26265 16083 26299
rect 16025 26259 16083 26265
rect 12820 26200 13216 26228
rect 13906 26188 13912 26240
rect 13964 26228 13970 26240
rect 14642 26228 14648 26240
rect 13964 26200 14648 26228
rect 13964 26188 13970 26200
rect 14642 26188 14648 26200
rect 14700 26188 14706 26240
rect 15470 26188 15476 26240
rect 15528 26228 15534 26240
rect 16132 26228 16160 26327
rect 16942 26324 16948 26336
rect 17000 26324 17006 26376
rect 17494 26324 17500 26376
rect 17552 26364 17558 26376
rect 17589 26367 17647 26373
rect 17589 26364 17601 26367
rect 17552 26336 17601 26364
rect 17552 26324 17558 26336
rect 17589 26333 17601 26336
rect 17635 26333 17647 26367
rect 18414 26364 18420 26376
rect 18375 26336 18420 26364
rect 17589 26327 17647 26333
rect 18414 26324 18420 26336
rect 18472 26324 18478 26376
rect 20088 26364 20116 26404
rect 21913 26401 21925 26404
rect 21959 26401 21971 26435
rect 22066 26432 22094 26472
rect 30469 26435 30527 26441
rect 30469 26432 30481 26435
rect 22066 26404 30481 26432
rect 21913 26395 21971 26401
rect 30469 26401 30481 26404
rect 30515 26401 30527 26435
rect 30469 26395 30527 26401
rect 18524 26336 20116 26364
rect 20165 26367 20223 26373
rect 17681 26299 17739 26305
rect 17681 26265 17693 26299
rect 17727 26296 17739 26299
rect 17954 26296 17960 26308
rect 17727 26268 17960 26296
rect 17727 26265 17739 26268
rect 17681 26259 17739 26265
rect 17954 26256 17960 26268
rect 18012 26256 18018 26308
rect 16298 26228 16304 26240
rect 15528 26200 16304 26228
rect 15528 26188 15534 26200
rect 16298 26188 16304 26200
rect 16356 26228 16362 26240
rect 18524 26228 18552 26336
rect 20165 26333 20177 26367
rect 20211 26364 20223 26367
rect 20622 26364 20628 26376
rect 20211 26336 20628 26364
rect 20211 26333 20223 26336
rect 20165 26327 20223 26333
rect 20622 26324 20628 26336
rect 20680 26364 20686 26376
rect 21361 26367 21419 26373
rect 21361 26364 21373 26367
rect 20680 26336 21373 26364
rect 20680 26324 20686 26336
rect 21361 26333 21373 26336
rect 21407 26333 21419 26367
rect 29825 26367 29883 26373
rect 29825 26364 29837 26367
rect 21361 26327 21419 26333
rect 22066 26336 29837 26364
rect 18690 26256 18696 26308
rect 18748 26296 18754 26308
rect 22066 26296 22094 26336
rect 29825 26333 29837 26336
rect 29871 26333 29883 26367
rect 29825 26327 29883 26333
rect 29917 26367 29975 26373
rect 29917 26333 29929 26367
rect 29963 26333 29975 26367
rect 29917 26327 29975 26333
rect 30561 26367 30619 26373
rect 30561 26333 30573 26367
rect 30607 26364 30619 26367
rect 31113 26367 31171 26373
rect 31113 26364 31125 26367
rect 30607 26336 31125 26364
rect 30607 26333 30619 26336
rect 30561 26327 30619 26333
rect 31113 26333 31125 26336
rect 31159 26364 31171 26367
rect 31159 26336 38240 26364
rect 31159 26333 31171 26336
rect 31113 26327 31171 26333
rect 18748 26268 22094 26296
rect 29932 26296 29960 26327
rect 37734 26296 37740 26308
rect 29932 26268 37740 26296
rect 18748 26256 18754 26268
rect 37734 26256 37740 26268
rect 37792 26256 37798 26308
rect 18598 26228 18604 26240
rect 16356 26200 18604 26228
rect 16356 26188 16362 26200
rect 18598 26188 18604 26200
rect 18656 26188 18662 26240
rect 38212 26237 38240 26336
rect 38197 26231 38255 26237
rect 38197 26228 38209 26231
rect 38107 26200 38209 26228
rect 38197 26197 38209 26200
rect 38243 26228 38255 26231
rect 38378 26228 38384 26240
rect 38243 26200 38384 26228
rect 38243 26197 38255 26200
rect 38197 26191 38255 26197
rect 38378 26188 38384 26200
rect 38436 26188 38442 26240
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 1949 26027 2007 26033
rect 1949 25993 1961 26027
rect 1995 26024 2007 26027
rect 2038 26024 2044 26036
rect 1995 25996 2044 26024
rect 1995 25993 2007 25996
rect 1949 25987 2007 25993
rect 2038 25984 2044 25996
rect 2096 25984 2102 26036
rect 4062 26024 4068 26036
rect 4023 25996 4068 26024
rect 4062 25984 4068 25996
rect 4120 25984 4126 26036
rect 4617 26027 4675 26033
rect 4617 25993 4629 26027
rect 4663 26024 4675 26027
rect 4982 26024 4988 26036
rect 4663 25996 4988 26024
rect 4663 25993 4675 25996
rect 4617 25987 4675 25993
rect 4982 25984 4988 25996
rect 5040 25984 5046 26036
rect 6733 26027 6791 26033
rect 6733 25993 6745 26027
rect 6779 26024 6791 26027
rect 13722 26024 13728 26036
rect 6779 25996 9897 26024
rect 13683 25996 13728 26024
rect 6779 25993 6791 25996
rect 6733 25987 6791 25993
rect 3237 25959 3295 25965
rect 3237 25925 3249 25959
rect 3283 25956 3295 25959
rect 4706 25956 4712 25968
rect 3283 25928 4712 25956
rect 3283 25925 3295 25928
rect 3237 25919 3295 25925
rect 4706 25916 4712 25928
rect 4764 25916 4770 25968
rect 6178 25916 6184 25968
rect 6236 25956 6242 25968
rect 7469 25959 7527 25965
rect 7469 25956 7481 25959
rect 6236 25928 7481 25956
rect 6236 25916 6242 25928
rect 7469 25925 7481 25928
rect 7515 25925 7527 25959
rect 9030 25956 9036 25968
rect 8991 25928 9036 25956
rect 7469 25919 7527 25925
rect 9030 25916 9036 25928
rect 9088 25916 9094 25968
rect 9306 25916 9312 25968
rect 9364 25956 9370 25968
rect 9766 25956 9772 25968
rect 9364 25928 9772 25956
rect 9364 25916 9370 25928
rect 9766 25916 9772 25928
rect 9824 25916 9830 25968
rect 9869 25965 9897 25996
rect 13722 25984 13728 25996
rect 13780 25984 13786 26036
rect 13906 25984 13912 26036
rect 13964 26024 13970 26036
rect 17221 26027 17279 26033
rect 13964 25996 17172 26024
rect 13964 25984 13970 25996
rect 9861 25959 9919 25965
rect 9861 25925 9873 25959
rect 9907 25925 9919 25959
rect 13078 25956 13084 25968
rect 13039 25928 13084 25956
rect 9861 25919 9919 25925
rect 13078 25916 13084 25928
rect 13136 25916 13142 25968
rect 13173 25959 13231 25965
rect 13173 25925 13185 25959
rect 13219 25956 13231 25959
rect 14090 25956 14096 25968
rect 13219 25928 14096 25956
rect 13219 25925 13231 25928
rect 13173 25919 13231 25925
rect 14090 25916 14096 25928
rect 14148 25916 14154 25968
rect 17144 25956 17172 25996
rect 17221 25993 17233 26027
rect 17267 26024 17279 26027
rect 18322 26024 18328 26036
rect 17267 25996 18328 26024
rect 17267 25993 17279 25996
rect 17221 25987 17279 25993
rect 18322 25984 18328 25996
rect 18380 25984 18386 26036
rect 18414 25984 18420 26036
rect 18472 26024 18478 26036
rect 19153 26027 19211 26033
rect 19153 26024 19165 26027
rect 18472 25996 19165 26024
rect 18472 25984 18478 25996
rect 19153 25993 19165 25996
rect 19199 25993 19211 26027
rect 19153 25987 19211 25993
rect 20530 25984 20536 26036
rect 20588 26024 20594 26036
rect 21085 26027 21143 26033
rect 21085 26024 21097 26027
rect 20588 25996 21097 26024
rect 20588 25984 20594 25996
rect 21085 25993 21097 25996
rect 21131 25993 21143 26027
rect 37826 26024 37832 26036
rect 37787 25996 37832 26024
rect 21085 25987 21143 25993
rect 37826 25984 37832 25996
rect 37884 25984 37890 26036
rect 19426 25956 19432 25968
rect 17144 25928 19432 25956
rect 19426 25916 19432 25928
rect 19484 25916 19490 25968
rect 20714 25916 20720 25968
rect 20772 25956 20778 25968
rect 22557 25959 22615 25965
rect 22557 25956 22569 25959
rect 20772 25928 21220 25956
rect 20772 25916 20778 25928
rect 1857 25891 1915 25897
rect 1857 25857 1869 25891
rect 1903 25857 1915 25891
rect 1857 25851 1915 25857
rect 2501 25891 2559 25897
rect 2501 25857 2513 25891
rect 2547 25888 2559 25891
rect 2774 25888 2780 25900
rect 2547 25860 2780 25888
rect 2547 25857 2559 25860
rect 2501 25851 2559 25857
rect 1872 25684 1900 25851
rect 2774 25848 2780 25860
rect 2832 25848 2838 25900
rect 3142 25888 3148 25900
rect 3103 25860 3148 25888
rect 3142 25848 3148 25860
rect 3200 25848 3206 25900
rect 3973 25891 4031 25897
rect 3973 25888 3985 25891
rect 3436 25860 3985 25888
rect 2958 25780 2964 25832
rect 3016 25820 3022 25832
rect 3436 25820 3464 25860
rect 3973 25857 3985 25860
rect 4019 25888 4031 25891
rect 4062 25888 4068 25900
rect 4019 25860 4068 25888
rect 4019 25857 4031 25860
rect 3973 25851 4031 25857
rect 4062 25848 4068 25860
rect 4120 25848 4126 25900
rect 4614 25848 4620 25900
rect 4672 25888 4678 25900
rect 5074 25888 5080 25900
rect 4672 25860 5080 25888
rect 4672 25848 4678 25860
rect 5074 25848 5080 25860
rect 5132 25848 5138 25900
rect 5169 25891 5227 25897
rect 5169 25857 5181 25891
rect 5215 25857 5227 25891
rect 5169 25851 5227 25857
rect 3016 25792 3464 25820
rect 3016 25780 3022 25792
rect 3786 25780 3792 25832
rect 3844 25820 3850 25832
rect 5184 25820 5212 25851
rect 5718 25848 5724 25900
rect 5776 25888 5782 25900
rect 5813 25891 5871 25897
rect 5813 25888 5825 25891
rect 5776 25860 5825 25888
rect 5776 25848 5782 25860
rect 5813 25857 5825 25860
rect 5859 25857 5871 25891
rect 5813 25851 5871 25857
rect 6641 25891 6699 25897
rect 6641 25857 6653 25891
rect 6687 25888 6699 25891
rect 6730 25888 6736 25900
rect 6687 25860 6736 25888
rect 6687 25857 6699 25860
rect 6641 25851 6699 25857
rect 6730 25848 6736 25860
rect 6788 25848 6794 25900
rect 10962 25888 10968 25900
rect 10923 25860 10968 25888
rect 10962 25848 10968 25860
rect 11020 25848 11026 25900
rect 11790 25848 11796 25900
rect 11848 25888 11854 25900
rect 11885 25891 11943 25897
rect 11885 25888 11897 25891
rect 11848 25860 11897 25888
rect 11848 25848 11854 25860
rect 11885 25857 11897 25860
rect 11931 25857 11943 25891
rect 11885 25851 11943 25857
rect 13630 25848 13636 25900
rect 13688 25888 13694 25900
rect 14369 25891 14427 25897
rect 14369 25888 14381 25891
rect 13688 25860 14381 25888
rect 13688 25848 13694 25860
rect 14369 25857 14381 25860
rect 14415 25857 14427 25891
rect 14369 25851 14427 25857
rect 14826 25848 14832 25900
rect 14884 25888 14890 25900
rect 15013 25891 15071 25897
rect 15013 25888 15025 25891
rect 14884 25860 15025 25888
rect 14884 25848 14890 25860
rect 15013 25857 15025 25860
rect 15059 25857 15071 25891
rect 15654 25888 15660 25900
rect 15615 25860 15660 25888
rect 15013 25851 15071 25857
rect 15654 25848 15660 25860
rect 15712 25848 15718 25900
rect 16298 25888 16304 25900
rect 16259 25860 16304 25888
rect 16298 25848 16304 25860
rect 16356 25848 16362 25900
rect 17129 25891 17187 25897
rect 17129 25857 17141 25891
rect 17175 25888 17187 25891
rect 17494 25888 17500 25900
rect 17175 25860 17500 25888
rect 17175 25857 17187 25860
rect 17129 25851 17187 25857
rect 17494 25848 17500 25860
rect 17552 25848 17558 25900
rect 17954 25888 17960 25900
rect 17915 25860 17960 25888
rect 17954 25848 17960 25860
rect 18012 25848 18018 25900
rect 19245 25891 19303 25897
rect 19245 25888 19257 25891
rect 18340 25860 19257 25888
rect 3844 25792 5212 25820
rect 3844 25780 3850 25792
rect 5626 25780 5632 25832
rect 5684 25820 5690 25832
rect 7377 25823 7435 25829
rect 7377 25820 7389 25823
rect 5684 25792 7389 25820
rect 5684 25780 5690 25792
rect 7377 25789 7389 25792
rect 7423 25789 7435 25823
rect 7377 25783 7435 25789
rect 7558 25780 7564 25832
rect 7616 25820 7622 25832
rect 8294 25820 8300 25832
rect 7616 25792 8300 25820
rect 7616 25780 7622 25792
rect 8294 25780 8300 25792
rect 8352 25820 8358 25832
rect 8481 25823 8539 25829
rect 8481 25820 8493 25823
rect 8352 25792 8493 25820
rect 8352 25780 8358 25792
rect 8481 25789 8493 25792
rect 8527 25789 8539 25823
rect 8481 25783 8539 25789
rect 9125 25823 9183 25829
rect 9125 25789 9137 25823
rect 9171 25789 9183 25823
rect 9766 25820 9772 25832
rect 9727 25792 9772 25820
rect 9125 25783 9183 25789
rect 2593 25755 2651 25761
rect 2593 25721 2605 25755
rect 2639 25752 2651 25755
rect 5166 25752 5172 25764
rect 2639 25724 5172 25752
rect 2639 25721 2651 25724
rect 2593 25715 2651 25721
rect 5166 25712 5172 25724
rect 5224 25712 5230 25764
rect 5261 25755 5319 25761
rect 5261 25721 5273 25755
rect 5307 25752 5319 25755
rect 7929 25755 7987 25761
rect 5307 25724 7880 25752
rect 5307 25721 5319 25724
rect 5261 25715 5319 25721
rect 2406 25684 2412 25696
rect 1872 25656 2412 25684
rect 2406 25644 2412 25656
rect 2464 25684 2470 25696
rect 3142 25684 3148 25696
rect 2464 25656 3148 25684
rect 2464 25644 2470 25656
rect 3142 25644 3148 25656
rect 3200 25644 3206 25696
rect 5905 25687 5963 25693
rect 5905 25653 5917 25687
rect 5951 25684 5963 25687
rect 6270 25684 6276 25696
rect 5951 25656 6276 25684
rect 5951 25653 5963 25656
rect 5905 25647 5963 25653
rect 6270 25644 6276 25656
rect 6328 25644 6334 25696
rect 7852 25684 7880 25724
rect 7929 25721 7941 25755
rect 7975 25752 7987 25755
rect 8662 25752 8668 25764
rect 7975 25724 8668 25752
rect 7975 25721 7987 25724
rect 7929 25715 7987 25721
rect 8662 25712 8668 25724
rect 8720 25712 8726 25764
rect 8202 25684 8208 25696
rect 7852 25656 8208 25684
rect 8202 25644 8208 25656
rect 8260 25644 8266 25696
rect 9140 25684 9168 25783
rect 9766 25780 9772 25792
rect 9824 25780 9830 25832
rect 9876 25792 13124 25820
rect 9214 25712 9220 25764
rect 9272 25752 9278 25764
rect 9876 25752 9904 25792
rect 9272 25724 9904 25752
rect 10321 25755 10379 25761
rect 9272 25712 9278 25724
rect 10321 25721 10333 25755
rect 10367 25752 10379 25755
rect 10594 25752 10600 25764
rect 10367 25724 10600 25752
rect 10367 25721 10379 25724
rect 10321 25715 10379 25721
rect 10594 25712 10600 25724
rect 10652 25712 10658 25764
rect 12434 25752 12440 25764
rect 10980 25724 12440 25752
rect 10980 25684 11008 25724
rect 12434 25712 12440 25724
rect 12492 25752 12498 25764
rect 12621 25755 12679 25761
rect 12621 25752 12633 25755
rect 12492 25724 12633 25752
rect 12492 25712 12498 25724
rect 12621 25721 12633 25724
rect 12667 25752 12679 25755
rect 12894 25752 12900 25764
rect 12667 25724 12900 25752
rect 12667 25721 12679 25724
rect 12621 25715 12679 25721
rect 12894 25712 12900 25724
rect 12952 25712 12958 25764
rect 13096 25752 13124 25792
rect 13538 25780 13544 25832
rect 13596 25820 13602 25832
rect 13906 25820 13912 25832
rect 13596 25792 13912 25820
rect 13596 25780 13602 25792
rect 13906 25780 13912 25792
rect 13964 25780 13970 25832
rect 14182 25820 14188 25832
rect 14143 25792 14188 25820
rect 14182 25780 14188 25792
rect 14240 25780 14246 25832
rect 17773 25823 17831 25829
rect 17773 25820 17785 25823
rect 14384 25792 17785 25820
rect 14384 25752 14412 25792
rect 17773 25789 17785 25792
rect 17819 25820 17831 25823
rect 18230 25820 18236 25832
rect 17819 25792 18236 25820
rect 17819 25789 17831 25792
rect 17773 25783 17831 25789
rect 18230 25780 18236 25792
rect 18288 25780 18294 25832
rect 13096 25724 14412 25752
rect 14458 25712 14464 25764
rect 14516 25752 14522 25764
rect 16209 25755 16267 25761
rect 16209 25752 16221 25755
rect 14516 25724 16221 25752
rect 14516 25712 14522 25724
rect 16209 25721 16221 25724
rect 16255 25721 16267 25755
rect 16209 25715 16267 25721
rect 17034 25712 17040 25764
rect 17092 25752 17098 25764
rect 18340 25752 18368 25860
rect 19245 25857 19257 25860
rect 19291 25888 19303 25891
rect 20990 25888 20996 25900
rect 19291 25860 20996 25888
rect 19291 25857 19303 25860
rect 19245 25851 19303 25857
rect 20990 25848 20996 25860
rect 21048 25848 21054 25900
rect 21192 25897 21220 25928
rect 22066 25928 22569 25956
rect 21177 25891 21235 25897
rect 21177 25857 21189 25891
rect 21223 25857 21235 25891
rect 21177 25851 21235 25857
rect 19886 25820 19892 25832
rect 19847 25792 19892 25820
rect 19886 25780 19892 25792
rect 19944 25780 19950 25832
rect 20073 25823 20131 25829
rect 20073 25789 20085 25823
rect 20119 25820 20131 25823
rect 21082 25820 21088 25832
rect 20119 25792 21088 25820
rect 20119 25789 20131 25792
rect 20073 25783 20131 25789
rect 21082 25780 21088 25792
rect 21140 25780 21146 25832
rect 17092 25724 18368 25752
rect 18417 25755 18475 25761
rect 17092 25712 17098 25724
rect 18417 25721 18429 25755
rect 18463 25752 18475 25755
rect 19242 25752 19248 25764
rect 18463 25724 19248 25752
rect 18463 25721 18475 25724
rect 18417 25715 18475 25721
rect 19242 25712 19248 25724
rect 19300 25752 19306 25764
rect 20257 25755 20315 25761
rect 20257 25752 20269 25755
rect 19300 25724 20269 25752
rect 19300 25712 19306 25724
rect 20257 25721 20269 25724
rect 20303 25721 20315 25755
rect 22066 25752 22094 25928
rect 22557 25925 22569 25928
rect 22603 25925 22615 25959
rect 22557 25919 22615 25925
rect 38013 25891 38071 25897
rect 38013 25857 38025 25891
rect 38059 25888 38071 25891
rect 38378 25888 38384 25900
rect 38059 25860 38384 25888
rect 38059 25857 38071 25860
rect 38013 25851 38071 25857
rect 38378 25848 38384 25860
rect 38436 25848 38442 25900
rect 20257 25715 20315 25721
rect 20364 25724 22094 25752
rect 9140 25656 11008 25684
rect 11057 25687 11115 25693
rect 11057 25653 11069 25687
rect 11103 25684 11115 25687
rect 11882 25684 11888 25696
rect 11103 25656 11888 25684
rect 11103 25653 11115 25656
rect 11057 25647 11115 25653
rect 11882 25644 11888 25656
rect 11940 25644 11946 25696
rect 11977 25687 12035 25693
rect 11977 25653 11989 25687
rect 12023 25684 12035 25687
rect 12526 25684 12532 25696
rect 12023 25656 12532 25684
rect 12023 25653 12035 25656
rect 11977 25647 12035 25653
rect 12526 25644 12532 25656
rect 12584 25644 12590 25696
rect 13170 25644 13176 25696
rect 13228 25684 13234 25696
rect 13722 25684 13728 25696
rect 13228 25656 13728 25684
rect 13228 25644 13234 25656
rect 13722 25644 13728 25656
rect 13780 25644 13786 25696
rect 13814 25644 13820 25696
rect 13872 25684 13878 25696
rect 14921 25687 14979 25693
rect 14921 25684 14933 25687
rect 13872 25656 14933 25684
rect 13872 25644 13878 25656
rect 14921 25653 14933 25656
rect 14967 25653 14979 25687
rect 15562 25684 15568 25696
rect 15523 25656 15568 25684
rect 14921 25647 14979 25653
rect 15562 25644 15568 25656
rect 15620 25644 15626 25696
rect 15654 25644 15660 25696
rect 15712 25684 15718 25696
rect 20364 25684 20392 25724
rect 15712 25656 20392 25684
rect 15712 25644 15718 25656
rect 20990 25644 20996 25696
rect 21048 25684 21054 25696
rect 22005 25687 22063 25693
rect 22005 25684 22017 25687
rect 21048 25656 22017 25684
rect 21048 25644 21054 25656
rect 22005 25653 22017 25656
rect 22051 25653 22063 25687
rect 22005 25647 22063 25653
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 1210 25440 1216 25492
rect 1268 25480 1274 25492
rect 2593 25483 2651 25489
rect 2593 25480 2605 25483
rect 1268 25452 2605 25480
rect 1268 25440 1274 25452
rect 2593 25449 2605 25452
rect 2639 25449 2651 25483
rect 2593 25443 2651 25449
rect 3237 25483 3295 25489
rect 3237 25449 3249 25483
rect 3283 25480 3295 25483
rect 3510 25480 3516 25492
rect 3283 25452 3516 25480
rect 3283 25449 3295 25452
rect 3237 25443 3295 25449
rect 3510 25440 3516 25452
rect 3568 25440 3574 25492
rect 3970 25440 3976 25492
rect 4028 25480 4034 25492
rect 4065 25483 4123 25489
rect 4065 25480 4077 25483
rect 4028 25452 4077 25480
rect 4028 25440 4034 25452
rect 4065 25449 4077 25452
rect 4111 25449 4123 25483
rect 5258 25480 5264 25492
rect 4065 25443 4123 25449
rect 4172 25452 5264 25480
rect 1949 25415 2007 25421
rect 1949 25381 1961 25415
rect 1995 25412 2007 25415
rect 4172 25412 4200 25452
rect 5258 25440 5264 25452
rect 5316 25440 5322 25492
rect 6178 25480 6184 25492
rect 6139 25452 6184 25480
rect 6178 25440 6184 25452
rect 6236 25440 6242 25492
rect 7926 25480 7932 25492
rect 7887 25452 7932 25480
rect 7926 25440 7932 25452
rect 7984 25440 7990 25492
rect 8018 25440 8024 25492
rect 8076 25480 8082 25492
rect 8076 25452 12434 25480
rect 8076 25440 8082 25452
rect 1995 25384 4200 25412
rect 4893 25415 4951 25421
rect 1995 25381 2007 25384
rect 1949 25375 2007 25381
rect 4893 25381 4905 25415
rect 4939 25412 4951 25415
rect 9030 25412 9036 25424
rect 4939 25384 9036 25412
rect 4939 25381 4951 25384
rect 4893 25375 4951 25381
rect 9030 25372 9036 25384
rect 9088 25372 9094 25424
rect 9306 25372 9312 25424
rect 9364 25412 9370 25424
rect 11698 25412 11704 25424
rect 9364 25384 11704 25412
rect 9364 25372 9370 25384
rect 11698 25372 11704 25384
rect 11756 25372 11762 25424
rect 12406 25412 12434 25452
rect 12618 25440 12624 25492
rect 12676 25480 12682 25492
rect 13725 25483 13783 25489
rect 13725 25480 13737 25483
rect 12676 25452 13737 25480
rect 12676 25440 12682 25452
rect 13725 25449 13737 25452
rect 13771 25480 13783 25483
rect 17497 25483 17555 25489
rect 13771 25452 16160 25480
rect 13771 25449 13783 25452
rect 13725 25443 13783 25449
rect 13538 25412 13544 25424
rect 12406 25384 13544 25412
rect 13538 25372 13544 25384
rect 13596 25372 13602 25424
rect 13630 25372 13636 25424
rect 13688 25412 13694 25424
rect 14918 25412 14924 25424
rect 13688 25384 14412 25412
rect 14879 25384 14924 25412
rect 13688 25372 13694 25384
rect 2958 25344 2964 25356
rect 1872 25316 2964 25344
rect 1872 25285 1900 25316
rect 2958 25304 2964 25316
rect 3016 25304 3022 25356
rect 3694 25304 3700 25356
rect 3752 25344 3758 25356
rect 5626 25344 5632 25356
rect 3752 25316 4936 25344
rect 5587 25316 5632 25344
rect 3752 25304 3758 25316
rect 1857 25279 1915 25285
rect 1857 25245 1869 25279
rect 1903 25245 1915 25279
rect 2498 25276 2504 25288
rect 2459 25248 2504 25276
rect 1857 25239 1915 25245
rect 2498 25236 2504 25248
rect 2556 25236 2562 25288
rect 2774 25236 2780 25288
rect 2832 25276 2838 25288
rect 3145 25279 3203 25285
rect 3145 25276 3157 25279
rect 2832 25248 3157 25276
rect 2832 25236 2838 25248
rect 3145 25245 3157 25248
rect 3191 25245 3203 25279
rect 4154 25276 4160 25288
rect 4067 25248 4160 25276
rect 3145 25239 3203 25245
rect 4154 25236 4160 25248
rect 4212 25276 4218 25288
rect 4798 25276 4804 25288
rect 4212 25248 4292 25276
rect 4759 25248 4804 25276
rect 4212 25236 4218 25248
rect 4264 25208 4292 25248
rect 4798 25236 4804 25248
rect 4856 25236 4862 25288
rect 4908 25276 4936 25316
rect 5626 25304 5632 25316
rect 5684 25304 5690 25356
rect 5994 25304 6000 25356
rect 6052 25344 6058 25356
rect 7561 25347 7619 25353
rect 7561 25344 7573 25347
rect 6052 25316 7573 25344
rect 6052 25304 6058 25316
rect 7561 25313 7573 25316
rect 7607 25313 7619 25347
rect 7561 25307 7619 25313
rect 8573 25347 8631 25353
rect 8573 25313 8585 25347
rect 8619 25344 8631 25347
rect 9490 25344 9496 25356
rect 8619 25316 9496 25344
rect 8619 25313 8631 25316
rect 8573 25307 8631 25313
rect 9490 25304 9496 25316
rect 9548 25304 9554 25356
rect 9858 25304 9864 25356
rect 9916 25344 9922 25356
rect 9953 25347 10011 25353
rect 9953 25344 9965 25347
rect 9916 25316 9965 25344
rect 9916 25304 9922 25316
rect 9953 25313 9965 25316
rect 9999 25313 10011 25347
rect 9953 25307 10011 25313
rect 11333 25347 11391 25353
rect 11333 25313 11345 25347
rect 11379 25344 11391 25347
rect 11422 25344 11428 25356
rect 11379 25316 11428 25344
rect 11379 25313 11391 25316
rect 11333 25307 11391 25313
rect 11422 25304 11428 25316
rect 11480 25304 11486 25356
rect 12434 25344 12440 25356
rect 12395 25316 12440 25344
rect 12434 25304 12440 25316
rect 12492 25304 12498 25356
rect 13078 25304 13084 25356
rect 13136 25344 13142 25356
rect 13814 25344 13820 25356
rect 13136 25316 13820 25344
rect 13136 25304 13142 25316
rect 13814 25304 13820 25316
rect 13872 25304 13878 25356
rect 14384 25353 14412 25384
rect 14918 25372 14924 25384
rect 14976 25372 14982 25424
rect 14369 25347 14427 25353
rect 14369 25313 14381 25347
rect 14415 25313 14427 25347
rect 14369 25307 14427 25313
rect 6089 25279 6147 25285
rect 6089 25276 6101 25279
rect 4908 25248 6101 25276
rect 6089 25245 6101 25248
rect 6135 25245 6147 25279
rect 6089 25239 6147 25245
rect 6733 25279 6791 25285
rect 6733 25245 6745 25279
rect 6779 25245 6791 25279
rect 6733 25239 6791 25245
rect 4982 25208 4988 25220
rect 4264 25180 4988 25208
rect 4982 25168 4988 25180
rect 5040 25168 5046 25220
rect 5166 25168 5172 25220
rect 5224 25208 5230 25220
rect 6362 25208 6368 25220
rect 5224 25180 6368 25208
rect 5224 25168 5230 25180
rect 6362 25168 6368 25180
rect 6420 25168 6426 25220
rect 5626 25100 5632 25152
rect 5684 25140 5690 25152
rect 6748 25140 6776 25239
rect 7282 25236 7288 25288
rect 7340 25276 7346 25288
rect 7377 25279 7435 25285
rect 7377 25276 7389 25279
rect 7340 25248 7389 25276
rect 7340 25236 7346 25248
rect 7377 25245 7389 25248
rect 7423 25245 7435 25279
rect 7377 25239 7435 25245
rect 11517 25279 11575 25285
rect 11517 25245 11529 25279
rect 11563 25245 11575 25279
rect 11517 25239 11575 25245
rect 6825 25211 6883 25217
rect 6825 25177 6837 25211
rect 6871 25208 6883 25211
rect 9122 25208 9128 25220
rect 6871 25180 9128 25208
rect 6871 25177 6883 25180
rect 6825 25171 6883 25177
rect 9122 25168 9128 25180
rect 9180 25208 9186 25220
rect 9677 25211 9735 25217
rect 9677 25208 9689 25211
rect 9180 25180 9689 25208
rect 9180 25168 9186 25180
rect 9677 25177 9689 25180
rect 9723 25177 9735 25211
rect 9677 25171 9735 25177
rect 9766 25168 9772 25220
rect 9824 25208 9830 25220
rect 11532 25208 11560 25239
rect 13630 25236 13636 25288
rect 13688 25236 13694 25288
rect 9824 25180 9869 25208
rect 9968 25180 11560 25208
rect 9824 25168 9830 25180
rect 8018 25140 8024 25152
rect 5684 25112 8024 25140
rect 5684 25100 5690 25112
rect 8018 25100 8024 25112
rect 8076 25100 8082 25152
rect 8294 25100 8300 25152
rect 8352 25140 8358 25152
rect 8478 25140 8484 25152
rect 8352 25112 8484 25140
rect 8352 25100 8358 25112
rect 8478 25100 8484 25112
rect 8536 25100 8542 25152
rect 8570 25100 8576 25152
rect 8628 25140 8634 25152
rect 9968 25140 9996 25180
rect 11698 25168 11704 25220
rect 11756 25208 11762 25220
rect 12989 25211 13047 25217
rect 12989 25208 13001 25211
rect 11756 25180 13001 25208
rect 11756 25168 11762 25180
rect 12989 25177 13001 25180
rect 13035 25177 13047 25211
rect 12989 25171 13047 25177
rect 13081 25211 13139 25217
rect 13081 25177 13093 25211
rect 13127 25208 13139 25211
rect 13648 25208 13676 25236
rect 14366 25208 14372 25220
rect 13127 25180 13676 25208
rect 13740 25180 14372 25208
rect 13127 25177 13139 25180
rect 13081 25171 13139 25177
rect 8628 25112 9996 25140
rect 8628 25100 8634 25112
rect 10226 25100 10232 25152
rect 10284 25140 10290 25152
rect 10781 25143 10839 25149
rect 10781 25140 10793 25143
rect 10284 25112 10793 25140
rect 10284 25100 10290 25112
rect 10781 25109 10793 25112
rect 10827 25140 10839 25143
rect 11422 25140 11428 25152
rect 10827 25112 11428 25140
rect 10827 25109 10839 25112
rect 10781 25103 10839 25109
rect 11422 25100 11428 25112
rect 11480 25100 11486 25152
rect 11977 25143 12035 25149
rect 11977 25109 11989 25143
rect 12023 25140 12035 25143
rect 13740 25140 13768 25180
rect 14366 25168 14372 25180
rect 14424 25168 14430 25220
rect 14458 25168 14464 25220
rect 14516 25208 14522 25220
rect 16132 25208 16160 25452
rect 17497 25449 17509 25483
rect 17543 25480 17555 25483
rect 17770 25480 17776 25492
rect 17543 25452 17776 25480
rect 17543 25449 17555 25452
rect 17497 25443 17555 25449
rect 17770 25440 17776 25452
rect 17828 25440 17834 25492
rect 21082 25480 21088 25492
rect 21043 25452 21088 25480
rect 21082 25440 21088 25452
rect 21140 25440 21146 25492
rect 18785 25415 18843 25421
rect 18785 25381 18797 25415
rect 18831 25412 18843 25415
rect 20438 25412 20444 25424
rect 18831 25384 20444 25412
rect 18831 25381 18843 25384
rect 18785 25375 18843 25381
rect 20438 25372 20444 25384
rect 20496 25372 20502 25424
rect 16209 25347 16267 25353
rect 16209 25313 16221 25347
rect 16255 25344 16267 25347
rect 17494 25344 17500 25356
rect 16255 25316 17500 25344
rect 16255 25313 16267 25316
rect 16209 25307 16267 25313
rect 17494 25304 17500 25316
rect 17552 25304 17558 25356
rect 18230 25344 18236 25356
rect 18191 25316 18236 25344
rect 18230 25304 18236 25316
rect 18288 25304 18294 25356
rect 26234 25304 26240 25356
rect 26292 25344 26298 25356
rect 26292 25316 29776 25344
rect 26292 25304 26298 25316
rect 16390 25276 16396 25288
rect 16351 25248 16396 25276
rect 16390 25236 16396 25248
rect 16448 25236 16454 25288
rect 17034 25276 17040 25288
rect 16947 25248 17040 25276
rect 17034 25236 17040 25248
rect 17092 25236 17098 25288
rect 17678 25276 17684 25288
rect 17639 25248 17684 25276
rect 17678 25236 17684 25248
rect 17736 25236 17742 25288
rect 20990 25236 20996 25288
rect 21048 25276 21054 25288
rect 29748 25285 29776 25316
rect 21177 25279 21235 25285
rect 21177 25276 21189 25279
rect 21048 25248 21189 25276
rect 21048 25236 21054 25248
rect 21177 25245 21189 25248
rect 21223 25276 21235 25279
rect 21637 25279 21695 25285
rect 21637 25276 21649 25279
rect 21223 25248 21649 25276
rect 21223 25245 21235 25248
rect 21177 25239 21235 25245
rect 21637 25245 21649 25248
rect 21683 25245 21695 25279
rect 28353 25279 28411 25285
rect 28353 25276 28365 25279
rect 21637 25239 21695 25245
rect 22112 25248 28365 25276
rect 17052 25208 17080 25236
rect 14516 25180 14561 25208
rect 16132 25180 17080 25208
rect 14516 25168 14522 25180
rect 18322 25168 18328 25220
rect 18380 25208 18386 25220
rect 18380 25180 18425 25208
rect 18380 25168 18386 25180
rect 19426 25168 19432 25220
rect 19484 25208 19490 25220
rect 19886 25208 19892 25220
rect 19484 25180 19892 25208
rect 19484 25168 19490 25180
rect 19886 25168 19892 25180
rect 19944 25168 19950 25220
rect 19978 25168 19984 25220
rect 20036 25208 20042 25220
rect 20036 25180 20081 25208
rect 20036 25168 20042 25180
rect 12023 25112 13768 25140
rect 12023 25109 12035 25112
rect 11977 25103 12035 25109
rect 13814 25100 13820 25152
rect 13872 25140 13878 25152
rect 15749 25143 15807 25149
rect 15749 25140 15761 25143
rect 13872 25112 15761 25140
rect 13872 25100 13878 25112
rect 15749 25109 15761 25112
rect 15795 25109 15807 25143
rect 15749 25103 15807 25109
rect 15838 25100 15844 25152
rect 15896 25140 15902 25152
rect 16945 25143 17003 25149
rect 16945 25140 16957 25143
rect 15896 25112 16957 25140
rect 15896 25100 15902 25112
rect 16945 25109 16957 25112
rect 16991 25109 17003 25143
rect 16945 25103 17003 25109
rect 17862 25100 17868 25152
rect 17920 25140 17926 25152
rect 22112 25140 22140 25248
rect 28353 25245 28365 25248
rect 28399 25245 28411 25279
rect 28353 25239 28411 25245
rect 29733 25279 29791 25285
rect 29733 25245 29745 25279
rect 29779 25245 29791 25279
rect 29733 25239 29791 25245
rect 37734 25236 37740 25288
rect 37792 25276 37798 25288
rect 37829 25279 37887 25285
rect 37829 25276 37841 25279
rect 37792 25248 37841 25276
rect 37792 25236 37798 25248
rect 37829 25245 37841 25248
rect 37875 25276 37887 25279
rect 38102 25276 38108 25288
rect 37875 25248 38108 25276
rect 37875 25245 37887 25248
rect 37829 25239 37887 25245
rect 38102 25236 38108 25248
rect 38160 25236 38166 25288
rect 28445 25211 28503 25217
rect 28445 25177 28457 25211
rect 28491 25208 28503 25211
rect 37274 25208 37280 25220
rect 28491 25180 37280 25208
rect 28491 25177 28503 25180
rect 28445 25171 28503 25177
rect 37274 25168 37280 25180
rect 37332 25168 37338 25220
rect 17920 25112 22140 25140
rect 29825 25143 29883 25149
rect 17920 25100 17926 25112
rect 29825 25109 29837 25143
rect 29871 25140 29883 25143
rect 36814 25140 36820 25152
rect 29871 25112 36820 25140
rect 29871 25109 29883 25112
rect 29825 25103 29883 25109
rect 36814 25100 36820 25112
rect 36872 25100 36878 25152
rect 38010 25140 38016 25152
rect 37971 25112 38016 25140
rect 38010 25100 38016 25112
rect 38068 25100 38074 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 7929 24939 7987 24945
rect 7929 24905 7941 24939
rect 7975 24936 7987 24939
rect 14182 24936 14188 24948
rect 7975 24908 14188 24936
rect 7975 24905 7987 24908
rect 7929 24899 7987 24905
rect 14182 24896 14188 24908
rect 14240 24896 14246 24948
rect 14826 24896 14832 24948
rect 14884 24936 14890 24948
rect 20070 24936 20076 24948
rect 14884 24908 20076 24936
rect 14884 24896 14890 24908
rect 20070 24896 20076 24908
rect 20128 24896 20134 24948
rect 2976 24840 3832 24868
rect 1857 24803 1915 24809
rect 1857 24769 1869 24803
rect 1903 24769 1915 24803
rect 1857 24763 1915 24769
rect 2317 24803 2375 24809
rect 2317 24769 2329 24803
rect 2363 24800 2375 24803
rect 2774 24800 2780 24812
rect 2363 24772 2780 24800
rect 2363 24769 2375 24772
rect 2317 24763 2375 24769
rect 1118 24624 1124 24676
rect 1176 24664 1182 24676
rect 1872 24664 1900 24763
rect 2774 24760 2780 24772
rect 2832 24800 2838 24812
rect 2976 24809 3004 24840
rect 2961 24803 3019 24809
rect 2961 24800 2973 24803
rect 2832 24772 2973 24800
rect 2832 24760 2838 24772
rect 2961 24769 2973 24772
rect 3007 24769 3019 24803
rect 3694 24800 3700 24812
rect 3655 24772 3700 24800
rect 2961 24763 3019 24769
rect 3694 24760 3700 24772
rect 3752 24760 3758 24812
rect 3804 24809 3832 24840
rect 8018 24828 8024 24880
rect 8076 24868 8082 24880
rect 9490 24868 9496 24880
rect 8076 24840 9496 24868
rect 8076 24828 8082 24840
rect 9490 24828 9496 24840
rect 9548 24868 9554 24880
rect 10594 24868 10600 24880
rect 9548 24840 9628 24868
rect 10555 24840 10600 24868
rect 9548 24828 9554 24840
rect 3789 24803 3847 24809
rect 3789 24769 3801 24803
rect 3835 24800 3847 24803
rect 3970 24800 3976 24812
rect 3835 24772 3976 24800
rect 3835 24769 3847 24772
rect 3789 24763 3847 24769
rect 3970 24760 3976 24772
rect 4028 24760 4034 24812
rect 4706 24760 4712 24812
rect 4764 24800 4770 24812
rect 4801 24803 4859 24809
rect 4801 24800 4813 24803
rect 4764 24772 4813 24800
rect 4764 24760 4770 24772
rect 4801 24769 4813 24772
rect 4847 24800 4859 24803
rect 5626 24800 5632 24812
rect 4847 24772 5632 24800
rect 4847 24769 4859 24772
rect 4801 24763 4859 24769
rect 5626 24760 5632 24772
rect 5684 24760 5690 24812
rect 5813 24803 5871 24809
rect 5813 24769 5825 24803
rect 5859 24769 5871 24803
rect 5813 24763 5871 24769
rect 5905 24803 5963 24809
rect 5905 24769 5917 24803
rect 5951 24800 5963 24803
rect 5994 24800 6000 24812
rect 5951 24772 6000 24800
rect 5951 24769 5963 24772
rect 5905 24763 5963 24769
rect 3053 24735 3111 24741
rect 3053 24701 3065 24735
rect 3099 24732 3111 24735
rect 4614 24732 4620 24744
rect 3099 24704 4620 24732
rect 3099 24701 3111 24704
rect 3053 24695 3111 24701
rect 4614 24692 4620 24704
rect 4672 24692 4678 24744
rect 5828 24732 5856 24763
rect 5994 24760 6000 24772
rect 6052 24760 6058 24812
rect 6733 24803 6791 24809
rect 6733 24769 6745 24803
rect 6779 24800 6791 24803
rect 7837 24803 7895 24809
rect 7837 24800 7849 24803
rect 6779 24772 7849 24800
rect 6779 24769 6791 24772
rect 6733 24763 6791 24769
rect 7837 24769 7849 24772
rect 7883 24800 7895 24803
rect 8294 24800 8300 24812
rect 7883 24772 8300 24800
rect 7883 24769 7895 24772
rect 7837 24763 7895 24769
rect 8294 24760 8300 24772
rect 8352 24760 8358 24812
rect 8478 24800 8484 24812
rect 8439 24772 8484 24800
rect 8478 24760 8484 24772
rect 8536 24760 8542 24812
rect 8573 24803 8631 24809
rect 8573 24769 8585 24803
rect 8619 24800 8631 24803
rect 8846 24800 8852 24812
rect 8619 24772 8852 24800
rect 8619 24769 8631 24772
rect 8573 24763 8631 24769
rect 8846 24760 8852 24772
rect 8904 24760 8910 24812
rect 9600 24800 9628 24840
rect 10594 24828 10600 24840
rect 10652 24828 10658 24880
rect 11882 24828 11888 24880
rect 11940 24868 11946 24880
rect 12345 24871 12403 24877
rect 12345 24868 12357 24871
rect 11940 24840 12357 24868
rect 11940 24828 11946 24840
rect 12345 24837 12357 24840
rect 12391 24837 12403 24871
rect 12345 24831 12403 24837
rect 12710 24828 12716 24880
rect 12768 24868 12774 24880
rect 15470 24868 15476 24880
rect 12768 24840 15476 24868
rect 12768 24828 12774 24840
rect 9769 24803 9827 24809
rect 9769 24800 9781 24803
rect 8956 24772 9444 24800
rect 9600 24772 9781 24800
rect 7006 24732 7012 24744
rect 5828 24704 7012 24732
rect 7006 24692 7012 24704
rect 7064 24692 7070 24744
rect 7377 24735 7435 24741
rect 7377 24701 7389 24735
rect 7423 24732 7435 24735
rect 8956 24732 8984 24772
rect 9122 24732 9128 24744
rect 7423 24704 8984 24732
rect 9083 24704 9128 24732
rect 7423 24701 7435 24704
rect 7377 24695 7435 24701
rect 9122 24692 9128 24704
rect 9180 24692 9186 24744
rect 9214 24692 9220 24744
rect 9272 24732 9278 24744
rect 9309 24735 9367 24741
rect 9309 24732 9321 24735
rect 9272 24704 9321 24732
rect 9272 24692 9278 24704
rect 9309 24701 9321 24704
rect 9355 24701 9367 24735
rect 9416 24732 9444 24772
rect 9769 24769 9781 24772
rect 9815 24769 9827 24803
rect 9769 24763 9827 24769
rect 12894 24760 12900 24812
rect 12952 24800 12958 24812
rect 13464 24809 13492 24840
rect 15470 24828 15476 24840
rect 15528 24828 15534 24880
rect 15749 24871 15807 24877
rect 15749 24837 15761 24871
rect 15795 24868 15807 24871
rect 15838 24868 15844 24880
rect 15795 24840 15844 24868
rect 15795 24837 15807 24840
rect 15749 24831 15807 24837
rect 15838 24828 15844 24840
rect 15896 24828 15902 24880
rect 19797 24871 19855 24877
rect 19797 24868 19809 24871
rect 19260 24840 19809 24868
rect 13449 24803 13507 24809
rect 12952 24772 12997 24800
rect 12952 24760 12958 24772
rect 13449 24769 13461 24803
rect 13495 24769 13507 24803
rect 14550 24800 14556 24812
rect 14511 24772 14556 24800
rect 13449 24763 13507 24769
rect 14550 24760 14556 24772
rect 14608 24760 14614 24812
rect 14734 24800 14740 24812
rect 14695 24772 14740 24800
rect 14734 24760 14740 24772
rect 14792 24760 14798 24812
rect 16316 24772 17356 24800
rect 10505 24735 10563 24741
rect 10505 24732 10517 24735
rect 9416 24704 10517 24732
rect 9309 24695 9367 24701
rect 10505 24701 10517 24704
rect 10551 24701 10563 24735
rect 10505 24695 10563 24701
rect 11514 24692 11520 24744
rect 11572 24732 11578 24744
rect 12253 24735 12311 24741
rect 12253 24732 12265 24735
rect 11572 24704 12265 24732
rect 11572 24692 11578 24704
rect 12253 24701 12265 24704
rect 12299 24732 12311 24735
rect 13078 24732 13084 24744
rect 12299 24704 13084 24732
rect 12299 24701 12311 24704
rect 12253 24695 12311 24701
rect 13078 24692 13084 24704
rect 13136 24692 13142 24744
rect 13262 24692 13268 24744
rect 13320 24732 13326 24744
rect 15654 24732 15660 24744
rect 13320 24704 15516 24732
rect 15615 24704 15660 24732
rect 13320 24692 13326 24704
rect 1176 24636 1808 24664
rect 1872 24636 9904 24664
rect 1176 24624 1182 24636
rect 1670 24596 1676 24608
rect 1631 24568 1676 24596
rect 1670 24556 1676 24568
rect 1728 24556 1734 24608
rect 1780 24596 1808 24636
rect 2409 24599 2467 24605
rect 2409 24596 2421 24599
rect 1780 24568 2421 24596
rect 2409 24565 2421 24568
rect 2455 24565 2467 24599
rect 2409 24559 2467 24565
rect 2498 24556 2504 24608
rect 2556 24596 2562 24608
rect 4154 24596 4160 24608
rect 2556 24568 4160 24596
rect 2556 24556 2562 24568
rect 4154 24556 4160 24568
rect 4212 24556 4218 24608
rect 5350 24596 5356 24608
rect 5311 24568 5356 24596
rect 5350 24556 5356 24568
rect 5408 24556 5414 24608
rect 6641 24599 6699 24605
rect 6641 24565 6653 24599
rect 6687 24596 6699 24599
rect 9674 24596 9680 24608
rect 6687 24568 9680 24596
rect 6687 24565 6699 24568
rect 6641 24559 6699 24565
rect 9674 24556 9680 24568
rect 9732 24556 9738 24608
rect 9876 24596 9904 24636
rect 9950 24624 9956 24676
rect 10008 24664 10014 24676
rect 11057 24667 11115 24673
rect 11057 24664 11069 24667
rect 10008 24636 11069 24664
rect 10008 24624 10014 24636
rect 11057 24633 11069 24636
rect 11103 24633 11115 24667
rect 12986 24664 12992 24676
rect 11057 24627 11115 24633
rect 11164 24636 12992 24664
rect 11164 24596 11192 24636
rect 12986 24624 12992 24636
rect 13044 24624 13050 24676
rect 13170 24624 13176 24676
rect 13228 24664 13234 24676
rect 14366 24664 14372 24676
rect 13228 24636 14228 24664
rect 14279 24636 14372 24664
rect 13228 24624 13234 24636
rect 9876 24568 11192 24596
rect 11422 24556 11428 24608
rect 11480 24596 11486 24608
rect 13354 24596 13360 24608
rect 11480 24568 13360 24596
rect 11480 24556 11486 24568
rect 13354 24556 13360 24568
rect 13412 24556 13418 24608
rect 13538 24596 13544 24608
rect 13499 24568 13544 24596
rect 13538 24556 13544 24568
rect 13596 24556 13602 24608
rect 13722 24556 13728 24608
rect 13780 24596 13786 24608
rect 13998 24596 14004 24608
rect 13780 24568 14004 24596
rect 13780 24556 13786 24568
rect 13998 24556 14004 24568
rect 14056 24556 14062 24608
rect 14200 24596 14228 24636
rect 14366 24624 14372 24636
rect 14424 24664 14430 24676
rect 15102 24664 15108 24676
rect 14424 24636 15108 24664
rect 14424 24624 14430 24636
rect 15102 24624 15108 24636
rect 15160 24624 15166 24676
rect 15488 24664 15516 24704
rect 15654 24692 15660 24704
rect 15712 24692 15718 24744
rect 16316 24732 16344 24772
rect 16850 24732 16856 24744
rect 16132 24704 16344 24732
rect 16811 24704 16856 24732
rect 16132 24664 16160 24704
rect 16850 24692 16856 24704
rect 16908 24692 16914 24744
rect 17328 24732 17356 24772
rect 17402 24760 17408 24812
rect 17460 24800 17466 24812
rect 17957 24803 18015 24809
rect 17957 24800 17969 24803
rect 17460 24772 17969 24800
rect 17460 24760 17466 24772
rect 17957 24769 17969 24772
rect 18003 24769 18015 24803
rect 17957 24763 18015 24769
rect 18601 24803 18659 24809
rect 18601 24769 18613 24803
rect 18647 24769 18659 24803
rect 18601 24763 18659 24769
rect 18693 24803 18751 24809
rect 18693 24769 18705 24803
rect 18739 24800 18751 24803
rect 19260 24800 19288 24840
rect 19797 24837 19809 24840
rect 19843 24837 19855 24871
rect 19797 24831 19855 24837
rect 38010 24800 38016 24812
rect 18739 24772 19288 24800
rect 37971 24772 38016 24800
rect 18739 24769 18751 24772
rect 18693 24763 18751 24769
rect 17862 24732 17868 24744
rect 17328 24704 17868 24732
rect 17862 24692 17868 24704
rect 17920 24732 17926 24744
rect 18616 24732 18644 24763
rect 38010 24760 38016 24772
rect 38068 24760 38074 24812
rect 19886 24732 19892 24744
rect 17920 24704 18644 24732
rect 19847 24704 19892 24732
rect 17920 24692 17926 24704
rect 19886 24692 19892 24704
rect 19944 24732 19950 24744
rect 20441 24735 20499 24741
rect 20441 24732 20453 24735
rect 19944 24704 20453 24732
rect 19944 24692 19950 24704
rect 20441 24701 20453 24704
rect 20487 24732 20499 24735
rect 20622 24732 20628 24744
rect 20487 24704 20628 24732
rect 20487 24701 20499 24704
rect 20441 24695 20499 24701
rect 20622 24692 20628 24704
rect 20680 24692 20686 24744
rect 15488 24636 16160 24664
rect 16209 24667 16267 24673
rect 16209 24633 16221 24667
rect 16255 24664 16267 24667
rect 18506 24664 18512 24676
rect 16255 24636 18512 24664
rect 16255 24633 16267 24636
rect 16209 24627 16267 24633
rect 18506 24624 18512 24636
rect 18564 24664 18570 24676
rect 18690 24664 18696 24676
rect 18564 24636 18696 24664
rect 18564 24624 18570 24636
rect 18690 24624 18696 24636
rect 18748 24624 18754 24676
rect 19334 24664 19340 24676
rect 19295 24636 19340 24664
rect 19334 24624 19340 24636
rect 19392 24624 19398 24676
rect 17678 24596 17684 24608
rect 14200 24568 17684 24596
rect 17678 24556 17684 24568
rect 17736 24556 17742 24608
rect 18049 24599 18107 24605
rect 18049 24565 18061 24599
rect 18095 24596 18107 24599
rect 18138 24596 18144 24608
rect 18095 24568 18144 24596
rect 18095 24565 18107 24568
rect 18049 24559 18107 24565
rect 18138 24556 18144 24568
rect 18196 24556 18202 24608
rect 38194 24596 38200 24608
rect 38155 24568 38200 24596
rect 38194 24556 38200 24568
rect 38252 24556 38258 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 1946 24392 1952 24404
rect 1907 24364 1952 24392
rect 1946 24352 1952 24364
rect 2004 24352 2010 24404
rect 2593 24395 2651 24401
rect 2593 24361 2605 24395
rect 2639 24392 2651 24395
rect 2682 24392 2688 24404
rect 2639 24364 2688 24392
rect 2639 24361 2651 24364
rect 2593 24355 2651 24361
rect 2682 24352 2688 24364
rect 2740 24352 2746 24404
rect 3970 24392 3976 24404
rect 3931 24364 3976 24392
rect 3970 24352 3976 24364
rect 4028 24352 4034 24404
rect 5445 24395 5503 24401
rect 5445 24361 5457 24395
rect 5491 24392 5503 24395
rect 5810 24392 5816 24404
rect 5491 24364 5816 24392
rect 5491 24361 5503 24364
rect 5445 24355 5503 24361
rect 5810 24352 5816 24364
rect 5868 24352 5874 24404
rect 7837 24395 7895 24401
rect 7837 24361 7849 24395
rect 7883 24392 7895 24395
rect 8570 24392 8576 24404
rect 7883 24364 8576 24392
rect 7883 24361 7895 24364
rect 7837 24355 7895 24361
rect 8570 24352 8576 24364
rect 8628 24352 8634 24404
rect 8662 24352 8668 24404
rect 8720 24392 8726 24404
rect 9674 24392 9680 24404
rect 8720 24364 9680 24392
rect 8720 24352 8726 24364
rect 9674 24352 9680 24364
rect 9732 24352 9738 24404
rect 12897 24395 12955 24401
rect 12897 24361 12909 24395
rect 12943 24392 12955 24395
rect 13814 24392 13820 24404
rect 12943 24364 13820 24392
rect 12943 24361 12955 24364
rect 12897 24355 12955 24361
rect 13814 24352 13820 24364
rect 13872 24352 13878 24404
rect 13998 24352 14004 24404
rect 14056 24392 14062 24404
rect 17034 24392 17040 24404
rect 14056 24364 17040 24392
rect 14056 24352 14062 24364
rect 17034 24352 17040 24364
rect 17092 24352 17098 24404
rect 17494 24392 17500 24404
rect 17455 24364 17500 24392
rect 17494 24352 17500 24364
rect 17552 24352 17558 24404
rect 18046 24392 18052 24404
rect 18007 24364 18052 24392
rect 18046 24352 18052 24364
rect 18104 24352 18110 24404
rect 18322 24352 18328 24404
rect 18380 24392 18386 24404
rect 18693 24395 18751 24401
rect 18693 24392 18705 24395
rect 18380 24364 18705 24392
rect 18380 24352 18386 24364
rect 18693 24361 18705 24364
rect 18739 24361 18751 24395
rect 18693 24355 18751 24361
rect 19613 24395 19671 24401
rect 19613 24361 19625 24395
rect 19659 24392 19671 24395
rect 19978 24392 19984 24404
rect 19659 24364 19984 24392
rect 19659 24361 19671 24364
rect 19613 24355 19671 24361
rect 19978 24352 19984 24364
rect 20036 24352 20042 24404
rect 20070 24352 20076 24404
rect 20128 24392 20134 24404
rect 20165 24395 20223 24401
rect 20165 24392 20177 24395
rect 20128 24364 20177 24392
rect 20128 24352 20134 24364
rect 20165 24361 20177 24364
rect 20211 24361 20223 24395
rect 20165 24355 20223 24361
rect 1762 24284 1768 24336
rect 1820 24324 1826 24336
rect 6457 24327 6515 24333
rect 6457 24324 6469 24327
rect 1820 24296 6469 24324
rect 1820 24284 1826 24296
rect 6457 24293 6469 24296
rect 6503 24293 6515 24327
rect 6457 24287 6515 24293
rect 8478 24284 8484 24336
rect 8536 24324 8542 24336
rect 13170 24324 13176 24336
rect 8536 24296 9444 24324
rect 8536 24284 8542 24296
rect 8294 24256 8300 24268
rect 7116 24228 8300 24256
rect 1857 24191 1915 24197
rect 1857 24157 1869 24191
rect 1903 24157 1915 24191
rect 2498 24188 2504 24200
rect 2459 24160 2504 24188
rect 1857 24151 1915 24157
rect 1872 24120 1900 24151
rect 2498 24148 2504 24160
rect 2556 24188 2562 24200
rect 7116 24197 7144 24228
rect 8294 24216 8300 24228
rect 8352 24216 8358 24268
rect 9306 24256 9312 24268
rect 8496 24228 9312 24256
rect 3145 24191 3203 24197
rect 3145 24188 3157 24191
rect 2556 24160 3157 24188
rect 2556 24148 2562 24160
rect 3145 24157 3157 24160
rect 3191 24157 3203 24191
rect 3145 24151 3203 24157
rect 6641 24191 6699 24197
rect 6641 24157 6653 24191
rect 6687 24157 6699 24191
rect 6641 24151 6699 24157
rect 7101 24191 7159 24197
rect 7101 24157 7113 24191
rect 7147 24157 7159 24191
rect 7742 24188 7748 24200
rect 7703 24160 7748 24188
rect 7101 24151 7159 24157
rect 2774 24120 2780 24132
rect 1872 24092 2780 24120
rect 2774 24080 2780 24092
rect 2832 24080 2838 24132
rect 5997 24123 6055 24129
rect 5997 24089 6009 24123
rect 6043 24120 6055 24123
rect 6656 24120 6684 24151
rect 7742 24148 7748 24160
rect 7800 24148 7806 24200
rect 7834 24148 7840 24200
rect 7892 24188 7898 24200
rect 8496 24197 8524 24228
rect 9306 24216 9312 24228
rect 9364 24216 9370 24268
rect 9416 24256 9444 24296
rect 9600 24296 13176 24324
rect 9600 24256 9628 24296
rect 13170 24284 13176 24296
rect 13228 24284 13234 24336
rect 15562 24324 15568 24336
rect 13280 24296 15568 24324
rect 9416 24228 9628 24256
rect 9674 24216 9680 24268
rect 9732 24256 9738 24268
rect 12437 24259 12495 24265
rect 9732 24228 9777 24256
rect 9732 24216 9738 24228
rect 12437 24225 12449 24259
rect 12483 24256 12495 24259
rect 12526 24256 12532 24268
rect 12483 24228 12532 24256
rect 12483 24225 12495 24228
rect 12437 24219 12495 24225
rect 12526 24216 12532 24228
rect 12584 24216 12590 24268
rect 8389 24191 8447 24197
rect 8389 24188 8401 24191
rect 7892 24160 8401 24188
rect 7892 24148 7898 24160
rect 8389 24157 8401 24160
rect 8435 24157 8447 24191
rect 8389 24151 8447 24157
rect 8481 24191 8539 24197
rect 8481 24157 8493 24191
rect 8527 24157 8539 24191
rect 10686 24188 10692 24200
rect 10647 24160 10692 24188
rect 8481 24151 8539 24157
rect 10686 24148 10692 24160
rect 10744 24148 10750 24200
rect 10870 24188 10876 24200
rect 10831 24160 10876 24188
rect 10870 24148 10876 24160
rect 10928 24148 10934 24200
rect 12250 24188 12256 24200
rect 12211 24160 12256 24188
rect 12250 24148 12256 24160
rect 12308 24188 12314 24200
rect 13280 24188 13308 24296
rect 15562 24284 15568 24296
rect 15620 24284 15626 24336
rect 20714 24324 20720 24336
rect 16960 24296 20720 24324
rect 13354 24216 13360 24268
rect 13412 24256 13418 24268
rect 15654 24256 15660 24268
rect 13412 24228 14412 24256
rect 13412 24216 13418 24228
rect 12308 24160 13308 24188
rect 13541 24191 13599 24197
rect 12308 24148 12314 24160
rect 13541 24157 13553 24191
rect 13587 24188 13599 24191
rect 13630 24188 13636 24200
rect 13587 24160 13636 24188
rect 13587 24157 13599 24160
rect 13541 24151 13599 24157
rect 13630 24148 13636 24160
rect 13688 24148 13694 24200
rect 14384 24197 14412 24228
rect 14476 24228 15660 24256
rect 14369 24191 14427 24197
rect 14369 24157 14381 24191
rect 14415 24157 14427 24191
rect 14369 24151 14427 24157
rect 8570 24120 8576 24132
rect 6043 24092 8576 24120
rect 6043 24089 6055 24092
rect 5997 24083 6055 24089
rect 8570 24080 8576 24092
rect 8628 24080 8634 24132
rect 8938 24080 8944 24132
rect 8996 24120 9002 24132
rect 9217 24123 9275 24129
rect 9217 24120 9229 24123
rect 8996 24092 9229 24120
rect 8996 24080 9002 24092
rect 9217 24089 9229 24092
rect 9263 24089 9275 24123
rect 9217 24083 9275 24089
rect 4798 24052 4804 24064
rect 4759 24024 4804 24052
rect 4798 24012 4804 24024
rect 4856 24012 4862 24064
rect 7190 24052 7196 24064
rect 7151 24024 7196 24052
rect 7190 24012 7196 24024
rect 7248 24012 7254 24064
rect 8294 24012 8300 24064
rect 8352 24052 8358 24064
rect 8754 24052 8760 24064
rect 8352 24024 8760 24052
rect 8352 24012 8358 24024
rect 8754 24012 8760 24024
rect 8812 24012 8818 24064
rect 9232 24052 9260 24083
rect 9306 24080 9312 24132
rect 9364 24120 9370 24132
rect 10704 24120 10732 24148
rect 14476 24120 14504 24228
rect 15654 24216 15660 24228
rect 15712 24216 15718 24268
rect 16301 24259 16359 24265
rect 16301 24225 16313 24259
rect 16347 24256 16359 24259
rect 16758 24256 16764 24268
rect 16347 24228 16764 24256
rect 16347 24225 16359 24228
rect 16301 24219 16359 24225
rect 16758 24216 16764 24228
rect 16816 24216 16822 24268
rect 14642 24148 14648 24200
rect 14700 24188 14706 24200
rect 16960 24197 16988 24296
rect 20714 24284 20720 24296
rect 20772 24284 20778 24336
rect 17862 24216 17868 24268
rect 17920 24256 17926 24268
rect 17920 24228 18644 24256
rect 17920 24216 17926 24228
rect 15013 24191 15071 24197
rect 15013 24188 15025 24191
rect 14700 24160 15025 24188
rect 14700 24148 14706 24160
rect 15013 24157 15025 24160
rect 15059 24157 15071 24191
rect 16945 24191 17003 24197
rect 16945 24188 16957 24191
rect 15013 24151 15071 24157
rect 16500 24160 16957 24188
rect 9364 24092 9409 24120
rect 10704 24092 14504 24120
rect 14553 24123 14611 24129
rect 9364 24080 9370 24092
rect 14553 24089 14565 24123
rect 14599 24120 14611 24123
rect 14918 24120 14924 24132
rect 14599 24092 14924 24120
rect 14599 24089 14611 24092
rect 14553 24083 14611 24089
rect 14918 24080 14924 24092
rect 14976 24080 14982 24132
rect 9582 24052 9588 24064
rect 9232 24024 9588 24052
rect 9582 24012 9588 24024
rect 9640 24012 9646 24064
rect 11333 24055 11391 24061
rect 11333 24021 11345 24055
rect 11379 24052 11391 24055
rect 11698 24052 11704 24064
rect 11379 24024 11704 24052
rect 11379 24021 11391 24024
rect 11333 24015 11391 24021
rect 11698 24012 11704 24024
rect 11756 24012 11762 24064
rect 13633 24055 13691 24061
rect 13633 24021 13645 24055
rect 13679 24052 13691 24055
rect 14734 24052 14740 24064
rect 13679 24024 14740 24052
rect 13679 24021 13691 24024
rect 13633 24015 13691 24021
rect 14734 24012 14740 24024
rect 14792 24012 14798 24064
rect 15028 24052 15056 24151
rect 15746 24080 15752 24132
rect 15804 24120 15810 24132
rect 15804 24092 15849 24120
rect 15804 24080 15810 24092
rect 16500 24052 16528 24160
rect 16945 24157 16957 24160
rect 16991 24157 17003 24191
rect 16945 24151 17003 24157
rect 17589 24191 17647 24197
rect 17589 24157 17601 24191
rect 17635 24188 17647 24191
rect 18046 24188 18052 24200
rect 17635 24160 18052 24188
rect 17635 24157 17647 24160
rect 17589 24151 17647 24157
rect 18046 24148 18052 24160
rect 18104 24148 18110 24200
rect 18616 24197 18644 24228
rect 18601 24191 18659 24197
rect 18601 24157 18613 24191
rect 18647 24157 18659 24191
rect 18601 24151 18659 24157
rect 19521 24191 19579 24197
rect 19521 24157 19533 24191
rect 19567 24157 19579 24191
rect 19521 24151 19579 24157
rect 18322 24080 18328 24132
rect 18380 24120 18386 24132
rect 19536 24120 19564 24151
rect 18380 24092 19564 24120
rect 18380 24080 18386 24092
rect 15028 24024 16528 24052
rect 16574 24012 16580 24064
rect 16632 24052 16638 24064
rect 16853 24055 16911 24061
rect 16853 24052 16865 24055
rect 16632 24024 16865 24052
rect 16632 24012 16638 24024
rect 16853 24021 16865 24024
rect 16899 24021 16911 24055
rect 16853 24015 16911 24021
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 934 23808 940 23860
rect 992 23848 998 23860
rect 1949 23851 2007 23857
rect 1949 23848 1961 23851
rect 992 23820 1961 23848
rect 992 23808 998 23820
rect 1949 23817 1961 23820
rect 1995 23817 2007 23851
rect 1949 23811 2007 23817
rect 2774 23808 2780 23860
rect 2832 23848 2838 23860
rect 3237 23851 3295 23857
rect 3237 23848 3249 23851
rect 2832 23820 3249 23848
rect 2832 23808 2838 23820
rect 3237 23817 3249 23820
rect 3283 23817 3295 23851
rect 3237 23811 3295 23817
rect 4062 23808 4068 23860
rect 4120 23848 4126 23860
rect 4249 23851 4307 23857
rect 4249 23848 4261 23851
rect 4120 23820 4261 23848
rect 4120 23808 4126 23820
rect 4249 23817 4261 23820
rect 4295 23817 4307 23851
rect 4249 23811 4307 23817
rect 4982 23808 4988 23860
rect 5040 23848 5046 23860
rect 5077 23851 5135 23857
rect 5077 23848 5089 23851
rect 5040 23820 5089 23848
rect 5040 23808 5046 23820
rect 5077 23817 5089 23820
rect 5123 23848 5135 23851
rect 5258 23848 5264 23860
rect 5123 23820 5264 23848
rect 5123 23817 5135 23820
rect 5077 23811 5135 23817
rect 5258 23808 5264 23820
rect 5316 23808 5322 23860
rect 7837 23851 7895 23857
rect 7837 23817 7849 23851
rect 7883 23848 7895 23851
rect 11698 23848 11704 23860
rect 7883 23820 10548 23848
rect 11659 23820 11704 23848
rect 7883 23817 7895 23820
rect 7837 23811 7895 23817
rect 2130 23740 2136 23792
rect 2188 23780 2194 23792
rect 5905 23783 5963 23789
rect 5905 23780 5917 23783
rect 2188 23752 5917 23780
rect 2188 23740 2194 23752
rect 5905 23749 5917 23752
rect 5951 23749 5963 23783
rect 5905 23743 5963 23749
rect 7190 23740 7196 23792
rect 7248 23780 7254 23792
rect 7248 23752 9260 23780
rect 7248 23740 7254 23752
rect 2041 23715 2099 23721
rect 2041 23681 2053 23715
rect 2087 23712 2099 23715
rect 2498 23712 2504 23724
rect 2087 23684 2504 23712
rect 2087 23681 2099 23684
rect 2041 23675 2099 23681
rect 2498 23672 2504 23684
rect 2556 23712 2562 23724
rect 7098 23712 7104 23724
rect 2556 23684 2636 23712
rect 7011 23684 7104 23712
rect 2556 23672 2562 23684
rect 2608 23576 2636 23684
rect 7098 23672 7104 23684
rect 7156 23672 7162 23724
rect 7742 23712 7748 23724
rect 7703 23684 7748 23712
rect 7742 23672 7748 23684
rect 7800 23672 7806 23724
rect 9232 23721 9260 23752
rect 9490 23740 9496 23792
rect 9548 23780 9554 23792
rect 10520 23789 10548 23820
rect 11698 23808 11704 23820
rect 11756 23808 11762 23860
rect 13354 23808 13360 23860
rect 13412 23848 13418 23860
rect 15562 23848 15568 23860
rect 13412 23820 15568 23848
rect 13412 23808 13418 23820
rect 15562 23808 15568 23820
rect 15620 23808 15626 23860
rect 15746 23808 15752 23860
rect 15804 23848 15810 23860
rect 16945 23851 17003 23857
rect 16945 23848 16957 23851
rect 15804 23820 16957 23848
rect 15804 23808 15810 23820
rect 16945 23817 16957 23820
rect 16991 23817 17003 23851
rect 16945 23811 17003 23817
rect 17034 23808 17040 23860
rect 17092 23848 17098 23860
rect 18322 23848 18328 23860
rect 17092 23820 18328 23848
rect 17092 23808 17098 23820
rect 18322 23808 18328 23820
rect 18380 23808 18386 23860
rect 27246 23848 27252 23860
rect 22066 23820 27252 23848
rect 9677 23783 9735 23789
rect 9677 23780 9689 23783
rect 9548 23752 9689 23780
rect 9548 23740 9554 23752
rect 9677 23749 9689 23752
rect 9723 23749 9735 23783
rect 9677 23743 9735 23749
rect 10505 23783 10563 23789
rect 10505 23749 10517 23783
rect 10551 23749 10563 23783
rect 10505 23743 10563 23749
rect 11057 23783 11115 23789
rect 11057 23749 11069 23783
rect 11103 23780 11115 23783
rect 11238 23780 11244 23792
rect 11103 23752 11244 23780
rect 11103 23749 11115 23752
rect 11057 23743 11115 23749
rect 11238 23740 11244 23752
rect 11296 23740 11302 23792
rect 11606 23740 11612 23792
rect 11664 23780 11670 23792
rect 13449 23783 13507 23789
rect 13449 23780 13461 23783
rect 11664 23752 13461 23780
rect 11664 23740 11670 23752
rect 13449 23749 13461 23752
rect 13495 23749 13507 23783
rect 13449 23743 13507 23749
rect 13538 23740 13544 23792
rect 13596 23780 13602 23792
rect 15657 23783 15715 23789
rect 15657 23780 15669 23783
rect 13596 23752 15669 23780
rect 13596 23740 13602 23752
rect 15657 23749 15669 23752
rect 15703 23749 15715 23783
rect 18138 23780 18144 23792
rect 18099 23752 18144 23780
rect 15657 23743 15715 23749
rect 18138 23740 18144 23752
rect 18196 23740 18202 23792
rect 18690 23780 18696 23792
rect 18651 23752 18696 23780
rect 18690 23740 18696 23752
rect 18748 23740 18754 23792
rect 8389 23715 8447 23721
rect 8389 23681 8401 23715
rect 8435 23681 8447 23715
rect 8389 23675 8447 23681
rect 8481 23715 8539 23721
rect 8481 23681 8493 23715
rect 8527 23712 8539 23715
rect 9217 23715 9275 23721
rect 8527 23684 9168 23712
rect 8527 23681 8539 23684
rect 8481 23675 8539 23681
rect 7116 23644 7144 23672
rect 7834 23644 7840 23656
rect 7116 23616 7840 23644
rect 7834 23604 7840 23616
rect 7892 23604 7898 23656
rect 8404 23644 8432 23675
rect 8846 23644 8852 23656
rect 8404 23616 8852 23644
rect 4614 23576 4620 23588
rect 2608 23548 4620 23576
rect 2608 23517 2636 23548
rect 4614 23536 4620 23548
rect 4672 23536 4678 23588
rect 7190 23576 7196 23588
rect 7151 23548 7196 23576
rect 7190 23536 7196 23548
rect 7248 23536 7254 23588
rect 2593 23511 2651 23517
rect 2593 23477 2605 23511
rect 2639 23508 2651 23511
rect 2682 23508 2688 23520
rect 2639 23480 2688 23508
rect 2639 23477 2651 23480
rect 2593 23471 2651 23477
rect 2682 23468 2688 23480
rect 2740 23468 2746 23520
rect 6641 23511 6699 23517
rect 6641 23477 6653 23511
rect 6687 23508 6699 23511
rect 8404 23508 8432 23616
rect 8846 23604 8852 23616
rect 8904 23604 8910 23656
rect 9030 23644 9036 23656
rect 8991 23616 9036 23644
rect 9030 23604 9036 23616
rect 9088 23604 9094 23656
rect 9140 23644 9168 23684
rect 9217 23681 9229 23715
rect 9263 23681 9275 23715
rect 9217 23675 9275 23681
rect 12250 23672 12256 23724
rect 12308 23712 12314 23724
rect 12345 23715 12403 23721
rect 12345 23712 12357 23715
rect 12308 23684 12357 23712
rect 12308 23672 12314 23684
rect 12345 23681 12357 23684
rect 12391 23681 12403 23715
rect 12345 23675 12403 23681
rect 13998 23672 14004 23724
rect 14056 23712 14062 23724
rect 14461 23715 14519 23721
rect 14461 23712 14473 23715
rect 14056 23684 14473 23712
rect 14056 23672 14062 23684
rect 14461 23681 14473 23684
rect 14507 23681 14519 23715
rect 17034 23712 17040 23724
rect 16995 23684 17040 23712
rect 14461 23675 14519 23681
rect 17034 23672 17040 23684
rect 17092 23672 17098 23724
rect 10042 23644 10048 23656
rect 9140 23616 10048 23644
rect 10042 23604 10048 23616
rect 10100 23604 10106 23656
rect 10413 23647 10471 23653
rect 10413 23613 10425 23647
rect 10459 23613 10471 23647
rect 10413 23607 10471 23613
rect 10318 23536 10324 23588
rect 10376 23576 10382 23588
rect 10428 23576 10456 23607
rect 11054 23604 11060 23656
rect 11112 23644 11118 23656
rect 12161 23647 12219 23653
rect 12161 23644 12173 23647
rect 11112 23616 12173 23644
rect 11112 23604 11118 23616
rect 12161 23613 12173 23616
rect 12207 23613 12219 23647
rect 12161 23607 12219 23613
rect 13357 23647 13415 23653
rect 13357 23613 13369 23647
rect 13403 23644 13415 23647
rect 13814 23644 13820 23656
rect 13403 23616 13820 23644
rect 13403 23613 13415 23616
rect 13357 23607 13415 23613
rect 13814 23604 13820 23616
rect 13872 23604 13878 23656
rect 15749 23647 15807 23653
rect 14476 23616 15700 23644
rect 10376 23548 10456 23576
rect 13909 23579 13967 23585
rect 10376 23536 10382 23548
rect 13909 23545 13921 23579
rect 13955 23576 13967 23579
rect 14366 23576 14372 23588
rect 13955 23548 14372 23576
rect 13955 23545 13967 23548
rect 13909 23539 13967 23545
rect 14366 23536 14372 23548
rect 14424 23536 14430 23588
rect 6687 23480 8432 23508
rect 6687 23477 6699 23480
rect 6641 23471 6699 23477
rect 8570 23468 8576 23520
rect 8628 23508 8634 23520
rect 13354 23508 13360 23520
rect 8628 23480 13360 23508
rect 8628 23468 8634 23480
rect 13354 23468 13360 23480
rect 13412 23468 13418 23520
rect 13630 23468 13636 23520
rect 13688 23508 13694 23520
rect 14476 23508 14504 23616
rect 15194 23576 15200 23588
rect 15107 23548 15200 23576
rect 15194 23536 15200 23548
rect 15252 23576 15258 23588
rect 15672 23576 15700 23616
rect 15749 23613 15761 23647
rect 15795 23644 15807 23647
rect 16850 23644 16856 23656
rect 15795 23616 16856 23644
rect 15795 23613 15807 23616
rect 15749 23607 15807 23613
rect 16850 23604 16856 23616
rect 16908 23604 16914 23656
rect 17770 23604 17776 23656
rect 17828 23644 17834 23656
rect 18049 23647 18107 23653
rect 18049 23644 18061 23647
rect 17828 23616 18061 23644
rect 17828 23604 17834 23616
rect 18049 23613 18061 23616
rect 18095 23644 18107 23647
rect 19153 23647 19211 23653
rect 19153 23644 19165 23647
rect 18095 23616 19165 23644
rect 18095 23613 18107 23616
rect 18049 23607 18107 23613
rect 19153 23613 19165 23616
rect 19199 23613 19211 23647
rect 19153 23607 19211 23613
rect 19705 23579 19763 23585
rect 19705 23576 19717 23579
rect 15252 23548 15608 23576
rect 15672 23548 19717 23576
rect 15252 23536 15258 23548
rect 13688 23480 14504 23508
rect 14553 23511 14611 23517
rect 13688 23468 13694 23480
rect 14553 23477 14565 23511
rect 14599 23508 14611 23511
rect 15378 23508 15384 23520
rect 14599 23480 15384 23508
rect 14599 23477 14611 23480
rect 14553 23471 14611 23477
rect 15378 23468 15384 23480
rect 15436 23468 15442 23520
rect 15580 23508 15608 23548
rect 19705 23545 19717 23548
rect 19751 23576 19763 23579
rect 22066 23576 22094 23820
rect 27246 23808 27252 23820
rect 27304 23808 27310 23860
rect 37274 23672 37280 23724
rect 37332 23712 37338 23724
rect 38013 23715 38071 23721
rect 38013 23712 38025 23715
rect 37332 23684 38025 23712
rect 37332 23672 37338 23684
rect 38013 23681 38025 23684
rect 38059 23681 38071 23715
rect 38013 23675 38071 23681
rect 19751 23548 22094 23576
rect 19751 23545 19763 23548
rect 19705 23539 19763 23545
rect 17586 23508 17592 23520
rect 15580 23480 17592 23508
rect 17586 23468 17592 23480
rect 17644 23468 17650 23520
rect 38194 23508 38200 23520
rect 38155 23480 38200 23508
rect 38194 23468 38200 23480
rect 38252 23468 38258 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 2774 23264 2780 23316
rect 2832 23304 2838 23316
rect 2961 23307 3019 23313
rect 2961 23304 2973 23307
rect 2832 23276 2973 23304
rect 2832 23264 2838 23276
rect 2961 23273 2973 23276
rect 3007 23304 3019 23307
rect 3973 23307 4031 23313
rect 3973 23304 3985 23307
rect 3007 23276 3985 23304
rect 3007 23273 3019 23276
rect 2961 23267 3019 23273
rect 3973 23273 3985 23276
rect 4019 23273 4031 23307
rect 4614 23304 4620 23316
rect 4575 23276 4620 23304
rect 3973 23267 4031 23273
rect 4614 23264 4620 23276
rect 4672 23264 4678 23316
rect 5169 23307 5227 23313
rect 5169 23273 5181 23307
rect 5215 23304 5227 23307
rect 5534 23304 5540 23316
rect 5215 23276 5540 23304
rect 5215 23273 5227 23276
rect 5169 23267 5227 23273
rect 5534 23264 5540 23276
rect 5592 23264 5598 23316
rect 5718 23304 5724 23316
rect 5679 23276 5724 23304
rect 5718 23264 5724 23276
rect 5776 23264 5782 23316
rect 6733 23307 6791 23313
rect 6733 23273 6745 23307
rect 6779 23304 6791 23307
rect 6822 23304 6828 23316
rect 6779 23276 6828 23304
rect 6779 23273 6791 23276
rect 6733 23267 6791 23273
rect 6822 23264 6828 23276
rect 6880 23264 6886 23316
rect 9677 23307 9735 23313
rect 9677 23273 9689 23307
rect 9723 23304 9735 23307
rect 11054 23304 11060 23316
rect 9723 23276 11060 23304
rect 9723 23273 9735 23276
rect 9677 23267 9735 23273
rect 11054 23264 11060 23276
rect 11112 23264 11118 23316
rect 11698 23264 11704 23316
rect 11756 23304 11762 23316
rect 12069 23307 12127 23313
rect 12069 23304 12081 23307
rect 11756 23276 12081 23304
rect 11756 23264 11762 23276
rect 12069 23273 12081 23276
rect 12115 23273 12127 23307
rect 12069 23267 12127 23273
rect 17678 23264 17684 23316
rect 17736 23304 17742 23316
rect 17773 23307 17831 23313
rect 17773 23304 17785 23307
rect 17736 23276 17785 23304
rect 17736 23264 17742 23276
rect 17773 23273 17785 23276
rect 17819 23304 17831 23307
rect 27246 23304 27252 23316
rect 17819 23276 22094 23304
rect 27207 23276 27252 23304
rect 17819 23273 17831 23276
rect 17773 23267 17831 23273
rect 8481 23239 8539 23245
rect 8481 23205 8493 23239
rect 8527 23236 8539 23239
rect 10686 23236 10692 23248
rect 8527 23208 10692 23236
rect 8527 23205 8539 23208
rect 8481 23199 8539 23205
rect 10686 23196 10692 23208
rect 10744 23196 10750 23248
rect 14366 23236 14372 23248
rect 14327 23208 14372 23236
rect 14366 23196 14372 23208
rect 14424 23196 14430 23248
rect 18417 23239 18475 23245
rect 18417 23205 18429 23239
rect 18463 23236 18475 23239
rect 18598 23236 18604 23248
rect 18463 23208 18604 23236
rect 18463 23205 18475 23208
rect 18417 23199 18475 23205
rect 18598 23196 18604 23208
rect 18656 23196 18662 23248
rect 7929 23171 7987 23177
rect 7929 23137 7941 23171
rect 7975 23168 7987 23171
rect 9030 23168 9036 23180
rect 7975 23140 9036 23168
rect 7975 23137 7987 23140
rect 7929 23131 7987 23137
rect 9030 23128 9036 23140
rect 9088 23128 9094 23180
rect 10502 23168 10508 23180
rect 9600 23140 10508 23168
rect 1762 23060 1768 23112
rect 1820 23100 1826 23112
rect 9600 23109 9628 23140
rect 10502 23128 10508 23140
rect 10560 23128 10566 23180
rect 10778 23168 10784 23180
rect 10739 23140 10784 23168
rect 10778 23128 10784 23140
rect 10836 23128 10842 23180
rect 11790 23128 11796 23180
rect 11848 23168 11854 23180
rect 16669 23171 16727 23177
rect 11848 23140 13492 23168
rect 11848 23128 11854 23140
rect 1949 23103 2007 23109
rect 1949 23100 1961 23103
rect 1820 23072 1961 23100
rect 1820 23060 1826 23072
rect 1949 23069 1961 23072
rect 1995 23100 2007 23103
rect 2409 23103 2467 23109
rect 2409 23100 2421 23103
rect 1995 23072 2421 23100
rect 1995 23069 2007 23072
rect 1949 23063 2007 23069
rect 2409 23069 2421 23072
rect 2455 23100 2467 23103
rect 7193 23103 7251 23109
rect 7193 23100 7205 23103
rect 2455 23072 7205 23100
rect 2455 23069 2467 23072
rect 2409 23063 2467 23069
rect 7193 23069 7205 23072
rect 7239 23100 7251 23103
rect 8389 23103 8447 23109
rect 8389 23100 8401 23103
rect 7239 23072 8401 23100
rect 7239 23069 7251 23072
rect 7193 23063 7251 23069
rect 8389 23069 8401 23072
rect 8435 23069 8447 23103
rect 8389 23063 8447 23069
rect 9585 23103 9643 23109
rect 9585 23069 9597 23103
rect 9631 23069 9643 23103
rect 9585 23063 9643 23069
rect 10962 23060 10968 23112
rect 11020 23100 11026 23112
rect 11425 23103 11483 23109
rect 11425 23100 11437 23103
rect 11020 23072 11437 23100
rect 11020 23060 11026 23072
rect 11425 23069 11437 23072
rect 11471 23069 11483 23103
rect 12526 23100 12532 23112
rect 12487 23072 12532 23100
rect 11425 23063 11483 23069
rect 12526 23060 12532 23072
rect 12584 23060 12590 23112
rect 13464 23109 13492 23140
rect 16669 23137 16681 23171
rect 16715 23168 16727 23171
rect 16758 23168 16764 23180
rect 16715 23140 16764 23168
rect 16715 23137 16727 23140
rect 16669 23131 16727 23137
rect 16758 23128 16764 23140
rect 16816 23128 16822 23180
rect 22066 23168 22094 23276
rect 27246 23264 27252 23276
rect 27304 23264 27310 23316
rect 27982 23304 27988 23316
rect 27943 23276 27988 23304
rect 27982 23264 27988 23276
rect 28040 23264 28046 23316
rect 33686 23168 33692 23180
rect 22066 23140 33692 23168
rect 33686 23128 33692 23140
rect 33744 23128 33750 23180
rect 12713 23103 12771 23109
rect 12713 23069 12725 23103
rect 12759 23069 12771 23103
rect 12713 23063 12771 23069
rect 13449 23103 13507 23109
rect 13449 23069 13461 23103
rect 13495 23100 13507 23103
rect 13998 23100 14004 23112
rect 13495 23072 14004 23100
rect 13495 23069 13507 23072
rect 13449 23063 13507 23069
rect 10318 23032 10324 23044
rect 10279 23004 10324 23032
rect 10318 22992 10324 23004
rect 10376 22992 10382 23044
rect 10410 22992 10416 23044
rect 10468 23032 10474 23044
rect 10468 23004 10513 23032
rect 10468 22992 10474 23004
rect 11146 22992 11152 23044
rect 11204 23032 11210 23044
rect 12342 23032 12348 23044
rect 11204 23004 12348 23032
rect 11204 22992 11210 23004
rect 12342 22992 12348 23004
rect 12400 23032 12406 23044
rect 12728 23032 12756 23063
rect 13998 23060 14004 23072
rect 14056 23060 14062 23112
rect 17313 23103 17371 23109
rect 17313 23069 17325 23103
rect 17359 23100 17371 23103
rect 17862 23100 17868 23112
rect 17359 23072 17868 23100
rect 17359 23069 17371 23072
rect 17313 23063 17371 23069
rect 17862 23060 17868 23072
rect 17920 23060 17926 23112
rect 27246 23060 27252 23112
rect 27304 23100 27310 23112
rect 27893 23103 27951 23109
rect 27893 23100 27905 23103
rect 27304 23072 27905 23100
rect 27304 23060 27310 23072
rect 27893 23069 27905 23072
rect 27939 23069 27951 23103
rect 27893 23063 27951 23069
rect 12400 23004 12756 23032
rect 12400 22992 12406 23004
rect 14090 22992 14096 23044
rect 14148 23032 14154 23044
rect 14829 23035 14887 23041
rect 14829 23032 14841 23035
rect 14148 23004 14841 23032
rect 14148 22992 14154 23004
rect 14829 23001 14841 23004
rect 14875 23001 14887 23035
rect 14829 22995 14887 23001
rect 14921 23035 14979 23041
rect 14921 23001 14933 23035
rect 14967 23032 14979 23035
rect 15562 23032 15568 23044
rect 14967 23004 15568 23032
rect 14967 23001 14979 23004
rect 14921 22995 14979 23001
rect 15562 22992 15568 23004
rect 15620 22992 15626 23044
rect 16022 23032 16028 23044
rect 15983 23004 16028 23032
rect 16022 22992 16028 23004
rect 16080 22992 16086 23044
rect 16117 23035 16175 23041
rect 16117 23001 16129 23035
rect 16163 23032 16175 23035
rect 16482 23032 16488 23044
rect 16163 23004 16488 23032
rect 16163 23001 16175 23004
rect 16117 22995 16175 23001
rect 16482 22992 16488 23004
rect 16540 22992 16546 23044
rect 1765 22967 1823 22973
rect 1765 22933 1777 22967
rect 1811 22964 1823 22967
rect 1854 22964 1860 22976
rect 1811 22936 1860 22964
rect 1811 22933 1823 22936
rect 1765 22927 1823 22933
rect 1854 22924 1860 22936
rect 1912 22924 1918 22976
rect 11514 22964 11520 22976
rect 11475 22936 11520 22964
rect 11514 22924 11520 22936
rect 11572 22924 11578 22976
rect 13354 22964 13360 22976
rect 13315 22936 13360 22964
rect 13354 22924 13360 22936
rect 13412 22924 13418 22976
rect 17126 22924 17132 22976
rect 17184 22964 17190 22976
rect 17221 22967 17279 22973
rect 17221 22964 17233 22967
rect 17184 22936 17233 22964
rect 17184 22924 17190 22936
rect 17221 22933 17233 22936
rect 17267 22933 17279 22967
rect 17221 22927 17279 22933
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 3142 22720 3148 22772
rect 3200 22760 3206 22772
rect 3421 22763 3479 22769
rect 3421 22760 3433 22763
rect 3200 22732 3433 22760
rect 3200 22720 3206 22732
rect 3421 22729 3433 22732
rect 3467 22760 3479 22763
rect 3510 22760 3516 22772
rect 3467 22732 3516 22760
rect 3467 22729 3479 22732
rect 3421 22723 3479 22729
rect 3510 22720 3516 22732
rect 3568 22720 3574 22772
rect 3878 22720 3884 22772
rect 3936 22760 3942 22772
rect 3973 22763 4031 22769
rect 3973 22760 3985 22763
rect 3936 22732 3985 22760
rect 3936 22720 3942 22732
rect 3973 22729 3985 22732
rect 4019 22729 4031 22763
rect 3973 22723 4031 22729
rect 4893 22763 4951 22769
rect 4893 22729 4905 22763
rect 4939 22760 4951 22763
rect 5166 22760 5172 22772
rect 4939 22732 5172 22760
rect 4939 22729 4951 22732
rect 4893 22723 4951 22729
rect 5166 22720 5172 22732
rect 5224 22760 5230 22772
rect 5442 22760 5448 22772
rect 5224 22732 5448 22760
rect 5224 22720 5230 22732
rect 5442 22720 5448 22732
rect 5500 22720 5506 22772
rect 5534 22720 5540 22772
rect 5592 22760 5598 22772
rect 6549 22763 6607 22769
rect 6549 22760 6561 22763
rect 5592 22732 6561 22760
rect 5592 22720 5598 22732
rect 6549 22729 6561 22732
rect 6595 22729 6607 22763
rect 6549 22723 6607 22729
rect 7285 22763 7343 22769
rect 7285 22729 7297 22763
rect 7331 22760 7343 22763
rect 7742 22760 7748 22772
rect 7331 22732 7748 22760
rect 7331 22729 7343 22732
rect 7285 22723 7343 22729
rect 7742 22720 7748 22732
rect 7800 22720 7806 22772
rect 9033 22763 9091 22769
rect 9033 22729 9045 22763
rect 9079 22760 9091 22763
rect 10410 22760 10416 22772
rect 9079 22732 10416 22760
rect 9079 22729 9091 22732
rect 9033 22723 9091 22729
rect 10410 22720 10416 22732
rect 10468 22720 10474 22772
rect 11514 22720 11520 22772
rect 11572 22760 11578 22772
rect 11572 22732 14228 22760
rect 11572 22720 11578 22732
rect 5258 22652 5264 22704
rect 5316 22692 5322 22704
rect 5353 22695 5411 22701
rect 5353 22692 5365 22695
rect 5316 22664 5365 22692
rect 5316 22652 5322 22664
rect 5353 22661 5365 22664
rect 5399 22661 5411 22695
rect 5353 22655 5411 22661
rect 8389 22695 8447 22701
rect 8389 22661 8401 22695
rect 8435 22692 8447 22695
rect 9306 22692 9312 22704
rect 8435 22664 9312 22692
rect 8435 22661 8447 22664
rect 8389 22655 8447 22661
rect 9306 22652 9312 22664
rect 9364 22652 9370 22704
rect 9677 22695 9735 22701
rect 9677 22661 9689 22695
rect 9723 22692 9735 22695
rect 10594 22692 10600 22704
rect 9723 22664 10600 22692
rect 9723 22661 9735 22664
rect 9677 22655 9735 22661
rect 10594 22652 10600 22664
rect 10652 22652 10658 22704
rect 14200 22701 14228 22732
rect 12989 22695 13047 22701
rect 12989 22692 13001 22695
rect 10704 22664 13001 22692
rect 1854 22624 1860 22636
rect 1815 22596 1860 22624
rect 1854 22584 1860 22596
rect 1912 22584 1918 22636
rect 3418 22584 3424 22636
rect 3476 22624 3482 22636
rect 8297 22627 8355 22633
rect 8297 22624 8309 22627
rect 3476 22596 8309 22624
rect 3476 22584 3482 22596
rect 8297 22593 8309 22596
rect 8343 22624 8355 22627
rect 8941 22627 8999 22633
rect 8941 22624 8953 22627
rect 8343 22596 8953 22624
rect 8343 22593 8355 22596
rect 8297 22587 8355 22593
rect 8941 22593 8953 22596
rect 8987 22593 8999 22627
rect 9582 22624 9588 22636
rect 9543 22596 9588 22624
rect 8941 22587 8999 22593
rect 9582 22584 9588 22596
rect 9640 22584 9646 22636
rect 10226 22624 10232 22636
rect 10139 22596 10232 22624
rect 10226 22584 10232 22596
rect 10284 22624 10290 22636
rect 10502 22624 10508 22636
rect 10284 22596 10508 22624
rect 10284 22584 10290 22596
rect 10502 22584 10508 22596
rect 10560 22584 10566 22636
rect 5994 22556 6000 22568
rect 5907 22528 6000 22556
rect 5994 22516 6000 22528
rect 6052 22556 6058 22568
rect 6546 22556 6552 22568
rect 6052 22528 6552 22556
rect 6052 22516 6058 22528
rect 6546 22516 6552 22528
rect 6604 22516 6610 22568
rect 7837 22559 7895 22565
rect 7837 22525 7849 22559
rect 7883 22556 7895 22559
rect 10244 22556 10272 22584
rect 7883 22528 10272 22556
rect 7883 22525 7895 22528
rect 7837 22519 7895 22525
rect 1670 22488 1676 22500
rect 1631 22460 1676 22488
rect 1670 22448 1676 22460
rect 1728 22448 1734 22500
rect 7926 22448 7932 22500
rect 7984 22488 7990 22500
rect 10704 22488 10732 22664
rect 12989 22661 13001 22664
rect 13035 22661 13047 22695
rect 12989 22655 13047 22661
rect 14185 22695 14243 22701
rect 14185 22661 14197 22695
rect 14231 22661 14243 22695
rect 17126 22692 17132 22704
rect 17087 22664 17132 22692
rect 14185 22655 14243 22661
rect 17126 22652 17132 22664
rect 17184 22652 17190 22704
rect 18417 22695 18475 22701
rect 18417 22661 18429 22695
rect 18463 22692 18475 22695
rect 19153 22695 19211 22701
rect 19153 22692 19165 22695
rect 18463 22664 19165 22692
rect 18463 22661 18475 22664
rect 18417 22655 18475 22661
rect 19153 22661 19165 22664
rect 19199 22661 19211 22695
rect 19153 22655 19211 22661
rect 11057 22627 11115 22633
rect 11057 22593 11069 22627
rect 11103 22624 11115 22627
rect 11238 22624 11244 22636
rect 11103 22596 11244 22624
rect 11103 22593 11115 22596
rect 11057 22587 11115 22593
rect 11238 22584 11244 22596
rect 11296 22584 11302 22636
rect 11701 22627 11759 22633
rect 11701 22593 11713 22627
rect 11747 22624 11759 22627
rect 12618 22624 12624 22636
rect 11747 22596 12624 22624
rect 11747 22593 11759 22596
rect 11701 22587 11759 22593
rect 12618 22584 12624 22596
rect 12676 22584 12682 22636
rect 14734 22584 14740 22636
rect 14792 22624 14798 22636
rect 15197 22627 15255 22633
rect 15197 22624 15209 22627
rect 14792 22596 15209 22624
rect 14792 22584 14798 22596
rect 15197 22593 15209 22596
rect 15243 22593 15255 22627
rect 15378 22624 15384 22636
rect 15339 22596 15384 22624
rect 15197 22587 15255 22593
rect 15378 22584 15384 22596
rect 15436 22584 15442 22636
rect 18322 22624 18328 22636
rect 18283 22596 18328 22624
rect 18322 22584 18328 22596
rect 18380 22584 18386 22636
rect 11885 22559 11943 22565
rect 11885 22556 11897 22559
rect 7984 22460 10732 22488
rect 10796 22528 11897 22556
rect 7984 22448 7990 22460
rect 2685 22423 2743 22429
rect 2685 22389 2697 22423
rect 2731 22420 2743 22423
rect 2774 22420 2780 22432
rect 2731 22392 2780 22420
rect 2731 22389 2743 22392
rect 2685 22383 2743 22389
rect 2774 22380 2780 22392
rect 2832 22420 2838 22432
rect 2958 22420 2964 22432
rect 2832 22392 2964 22420
rect 2832 22380 2838 22392
rect 2958 22380 2964 22392
rect 3016 22380 3022 22432
rect 10321 22423 10379 22429
rect 10321 22389 10333 22423
rect 10367 22420 10379 22423
rect 10796 22420 10824 22528
rect 11885 22525 11897 22528
rect 11931 22525 11943 22559
rect 11885 22519 11943 22525
rect 12897 22559 12955 22565
rect 12897 22525 12909 22559
rect 12943 22556 12955 22559
rect 13538 22556 13544 22568
rect 12943 22528 13544 22556
rect 12943 22525 12955 22528
rect 12897 22519 12955 22525
rect 13538 22516 13544 22528
rect 13596 22516 13602 22568
rect 14090 22556 14096 22568
rect 14051 22528 14096 22556
rect 14090 22516 14096 22528
rect 14148 22516 14154 22568
rect 17037 22559 17095 22565
rect 17037 22525 17049 22559
rect 17083 22556 17095 22559
rect 17126 22556 17132 22568
rect 17083 22528 17132 22556
rect 17083 22525 17095 22528
rect 17037 22519 17095 22525
rect 17126 22516 17132 22528
rect 17184 22516 17190 22568
rect 17313 22559 17371 22565
rect 17313 22525 17325 22559
rect 17359 22525 17371 22559
rect 17313 22519 17371 22525
rect 13449 22491 13507 22497
rect 13449 22457 13461 22491
rect 13495 22488 13507 22491
rect 14366 22488 14372 22500
rect 13495 22460 14372 22488
rect 13495 22457 13507 22460
rect 13449 22451 13507 22457
rect 14366 22448 14372 22460
rect 14424 22448 14430 22500
rect 14645 22491 14703 22497
rect 14645 22457 14657 22491
rect 14691 22488 14703 22491
rect 15194 22488 15200 22500
rect 14691 22460 15200 22488
rect 14691 22457 14703 22460
rect 14645 22451 14703 22457
rect 15194 22448 15200 22460
rect 15252 22448 15258 22500
rect 15562 22488 15568 22500
rect 15523 22460 15568 22488
rect 15562 22448 15568 22460
rect 15620 22448 15626 22500
rect 16758 22448 16764 22500
rect 16816 22488 16822 22500
rect 17328 22488 17356 22519
rect 17862 22516 17868 22568
rect 17920 22556 17926 22568
rect 19061 22559 19119 22565
rect 19061 22556 19073 22559
rect 17920 22528 19073 22556
rect 17920 22516 17926 22528
rect 19061 22525 19073 22528
rect 19107 22525 19119 22559
rect 19334 22556 19340 22568
rect 19295 22528 19340 22556
rect 19061 22519 19119 22525
rect 19334 22516 19340 22528
rect 19392 22516 19398 22568
rect 16816 22460 17356 22488
rect 16816 22448 16822 22460
rect 10962 22420 10968 22432
rect 10367 22392 10824 22420
rect 10923 22392 10968 22420
rect 10367 22389 10379 22392
rect 10321 22383 10379 22389
rect 10962 22380 10968 22392
rect 11020 22380 11026 22432
rect 12158 22420 12164 22432
rect 12119 22392 12164 22420
rect 12158 22380 12164 22392
rect 12216 22380 12222 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 5169 22219 5227 22225
rect 5169 22185 5181 22219
rect 5215 22216 5227 22219
rect 5258 22216 5264 22228
rect 5215 22188 5264 22216
rect 5215 22185 5227 22188
rect 5169 22179 5227 22185
rect 5258 22176 5264 22188
rect 5316 22216 5322 22228
rect 5994 22216 6000 22228
rect 5316 22188 6000 22216
rect 5316 22176 5322 22188
rect 5994 22176 6000 22188
rect 6052 22216 6058 22228
rect 6457 22219 6515 22225
rect 6457 22216 6469 22219
rect 6052 22188 6469 22216
rect 6052 22176 6058 22188
rect 6457 22185 6469 22188
rect 6503 22185 6515 22219
rect 6457 22179 6515 22185
rect 8573 22219 8631 22225
rect 8573 22185 8585 22219
rect 8619 22216 8631 22219
rect 8846 22216 8852 22228
rect 8619 22188 8852 22216
rect 8619 22185 8631 22188
rect 8573 22179 8631 22185
rect 8846 22176 8852 22188
rect 8904 22216 8910 22228
rect 9582 22216 9588 22228
rect 8904 22188 9588 22216
rect 8904 22176 8910 22188
rect 9582 22176 9588 22188
rect 9640 22176 9646 22228
rect 10244 22120 11192 22148
rect 2225 22083 2283 22089
rect 2225 22049 2237 22083
rect 2271 22080 2283 22083
rect 2774 22080 2780 22092
rect 2271 22052 2780 22080
rect 2271 22049 2283 22052
rect 2225 22043 2283 22049
rect 2774 22040 2780 22052
rect 2832 22080 2838 22092
rect 4062 22080 4068 22092
rect 2832 22052 4068 22080
rect 2832 22040 2838 22052
rect 4062 22040 4068 22052
rect 4120 22040 4126 22092
rect 4617 22083 4675 22089
rect 4617 22049 4629 22083
rect 4663 22080 4675 22083
rect 5074 22080 5080 22092
rect 4663 22052 5080 22080
rect 4663 22049 4675 22052
rect 4617 22043 4675 22049
rect 5074 22040 5080 22052
rect 5132 22040 5138 22092
rect 7101 22083 7159 22089
rect 7101 22049 7113 22083
rect 7147 22080 7159 22083
rect 7374 22080 7380 22092
rect 7147 22052 7380 22080
rect 7147 22049 7159 22052
rect 7101 22043 7159 22049
rect 7374 22040 7380 22052
rect 7432 22040 7438 22092
rect 8202 22040 8208 22092
rect 8260 22080 8266 22092
rect 10244 22080 10272 22120
rect 10410 22080 10416 22092
rect 8260 22052 10272 22080
rect 10371 22052 10416 22080
rect 8260 22040 8266 22052
rect 10410 22040 10416 22052
rect 10468 22080 10474 22092
rect 10468 22052 11100 22080
rect 10468 22040 10474 22052
rect 1673 22015 1731 22021
rect 1673 21981 1685 22015
rect 1719 22012 1731 22015
rect 3421 22015 3479 22021
rect 3421 22012 3433 22015
rect 1719 21984 3433 22012
rect 1719 21981 1731 21984
rect 1673 21975 1731 21981
rect 3421 21981 3433 21984
rect 3467 22012 3479 22015
rect 3510 22012 3516 22024
rect 3467 21984 3516 22012
rect 3467 21981 3479 21984
rect 3421 21975 3479 21981
rect 3510 21972 3516 21984
rect 3568 22012 3574 22024
rect 4890 22012 4896 22024
rect 3568 21984 4896 22012
rect 3568 21972 3574 21984
rect 4890 21972 4896 21984
rect 4948 22012 4954 22024
rect 7561 22015 7619 22021
rect 7561 22012 7573 22015
rect 4948 21984 7573 22012
rect 4948 21972 4954 21984
rect 7561 21981 7573 21984
rect 7607 21981 7619 22015
rect 7561 21975 7619 21981
rect 10594 21944 10600 21956
rect 10555 21916 10600 21944
rect 10594 21904 10600 21916
rect 10652 21904 10658 21956
rect 10686 21904 10692 21956
rect 10744 21944 10750 21956
rect 10744 21916 10789 21944
rect 10744 21904 10750 21916
rect 2869 21879 2927 21885
rect 2869 21845 2881 21879
rect 2915 21876 2927 21879
rect 2958 21876 2964 21888
rect 2915 21848 2964 21876
rect 2915 21845 2927 21848
rect 2869 21839 2927 21845
rect 2958 21836 2964 21848
rect 3016 21876 3022 21888
rect 4065 21879 4123 21885
rect 4065 21876 4077 21879
rect 3016 21848 4077 21876
rect 3016 21836 3022 21848
rect 4065 21845 4077 21848
rect 4111 21845 4123 21879
rect 4065 21839 4123 21845
rect 9585 21879 9643 21885
rect 9585 21845 9597 21879
rect 9631 21876 9643 21879
rect 10502 21876 10508 21888
rect 9631 21848 10508 21876
rect 9631 21845 9643 21848
rect 9585 21839 9643 21845
rect 10502 21836 10508 21848
rect 10560 21836 10566 21888
rect 11072 21876 11100 22052
rect 11164 21944 11192 22120
rect 12342 22108 12348 22160
rect 12400 22148 12406 22160
rect 12400 22120 14964 22148
rect 12400 22108 12406 22120
rect 11333 22083 11391 22089
rect 11333 22049 11345 22083
rect 11379 22080 11391 22083
rect 11698 22080 11704 22092
rect 11379 22052 11704 22080
rect 11379 22049 11391 22052
rect 11333 22043 11391 22049
rect 11698 22040 11704 22052
rect 11756 22040 11762 22092
rect 12805 22083 12863 22089
rect 12805 22049 12817 22083
rect 12851 22080 12863 22083
rect 13354 22080 13360 22092
rect 12851 22052 13360 22080
rect 12851 22049 12863 22052
rect 12805 22043 12863 22049
rect 13354 22040 13360 22052
rect 13412 22040 13418 22092
rect 13814 22040 13820 22092
rect 13872 22080 13878 22092
rect 14553 22083 14611 22089
rect 14553 22080 14565 22083
rect 13872 22052 14565 22080
rect 13872 22040 13878 22052
rect 14553 22049 14565 22052
rect 14599 22049 14611 22083
rect 14553 22043 14611 22049
rect 12618 22012 12624 22024
rect 12579 21984 12624 22012
rect 12618 21972 12624 21984
rect 12676 21972 12682 22024
rect 14936 22012 14964 22120
rect 15013 22083 15071 22089
rect 15013 22049 15025 22083
rect 15059 22080 15071 22083
rect 15749 22083 15807 22089
rect 15749 22080 15761 22083
rect 15059 22052 15761 22080
rect 15059 22049 15071 22052
rect 15013 22043 15071 22049
rect 15749 22049 15761 22052
rect 15795 22049 15807 22083
rect 15749 22043 15807 22049
rect 15197 22015 15255 22021
rect 15197 22012 15209 22015
rect 14936 21984 15209 22012
rect 15197 21981 15209 21984
rect 15243 22012 15255 22015
rect 15286 22012 15292 22024
rect 15243 21984 15292 22012
rect 15243 21981 15255 21984
rect 15197 21975 15255 21981
rect 15286 21972 15292 21984
rect 15344 21972 15350 22024
rect 15841 22015 15899 22021
rect 15841 21981 15853 22015
rect 15887 22012 15899 22015
rect 16485 22015 16543 22021
rect 16485 22012 16497 22015
rect 15887 21984 16497 22012
rect 15887 21981 15899 21984
rect 15841 21975 15899 21981
rect 16485 21981 16497 21984
rect 16531 22012 16543 22015
rect 16531 21984 17080 22012
rect 16531 21981 16543 21984
rect 16485 21975 16543 21981
rect 11425 21947 11483 21953
rect 11425 21944 11437 21947
rect 11164 21916 11437 21944
rect 11425 21913 11437 21916
rect 11471 21913 11483 21947
rect 11425 21907 11483 21913
rect 11977 21947 12035 21953
rect 11977 21913 11989 21947
rect 12023 21913 12035 21947
rect 11977 21907 12035 21913
rect 11992 21876 12020 21907
rect 12066 21904 12072 21956
rect 12124 21944 12130 21956
rect 15856 21944 15884 21975
rect 17052 21953 17080 21984
rect 12124 21916 15884 21944
rect 17037 21947 17095 21953
rect 12124 21904 12130 21916
rect 17037 21913 17049 21947
rect 17083 21944 17095 21947
rect 18325 21947 18383 21953
rect 18325 21944 18337 21947
rect 17083 21916 18337 21944
rect 17083 21913 17095 21916
rect 17037 21907 17095 21913
rect 18325 21913 18337 21916
rect 18371 21913 18383 21947
rect 18325 21907 18383 21913
rect 11072 21848 12020 21876
rect 13265 21879 13323 21885
rect 13265 21845 13277 21879
rect 13311 21876 13323 21879
rect 13538 21876 13544 21888
rect 13311 21848 13544 21876
rect 13311 21845 13323 21848
rect 13265 21839 13323 21845
rect 13538 21836 13544 21848
rect 13596 21836 13602 21888
rect 15654 21836 15660 21888
rect 15712 21876 15718 21888
rect 16393 21879 16451 21885
rect 16393 21876 16405 21879
rect 15712 21848 16405 21876
rect 15712 21836 15718 21848
rect 16393 21845 16405 21848
rect 16439 21845 16451 21879
rect 16393 21839 16451 21845
rect 17126 21836 17132 21888
rect 17184 21876 17190 21888
rect 17770 21876 17776 21888
rect 17184 21848 17776 21876
rect 17184 21836 17190 21848
rect 17770 21836 17776 21848
rect 17828 21836 17834 21888
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 2409 21675 2467 21681
rect 2409 21641 2421 21675
rect 2455 21672 2467 21675
rect 2774 21672 2780 21684
rect 2455 21644 2780 21672
rect 2455 21641 2467 21644
rect 2409 21635 2467 21641
rect 2774 21632 2780 21644
rect 2832 21632 2838 21684
rect 2866 21632 2872 21684
rect 2924 21672 2930 21684
rect 3789 21675 3847 21681
rect 3789 21672 3801 21675
rect 2924 21644 3801 21672
rect 2924 21632 2930 21644
rect 3789 21641 3801 21644
rect 3835 21641 3847 21675
rect 4982 21672 4988 21684
rect 4943 21644 4988 21672
rect 3789 21635 3847 21641
rect 4982 21632 4988 21644
rect 5040 21632 5046 21684
rect 5813 21675 5871 21681
rect 5813 21641 5825 21675
rect 5859 21672 5871 21675
rect 6178 21672 6184 21684
rect 5859 21644 6184 21672
rect 5859 21641 5871 21644
rect 5813 21635 5871 21641
rect 6178 21632 6184 21644
rect 6236 21632 6242 21684
rect 6546 21672 6552 21684
rect 6507 21644 6552 21672
rect 6546 21632 6552 21644
rect 6604 21632 6610 21684
rect 11149 21675 11207 21681
rect 11149 21641 11161 21675
rect 11195 21672 11207 21675
rect 12158 21672 12164 21684
rect 11195 21644 12164 21672
rect 11195 21641 11207 21644
rect 11149 21635 11207 21641
rect 12158 21632 12164 21644
rect 12216 21632 12222 21684
rect 2792 21604 2820 21632
rect 3237 21607 3295 21613
rect 3237 21604 3249 21607
rect 2792 21576 3249 21604
rect 3237 21573 3249 21576
rect 3283 21573 3295 21607
rect 3237 21567 3295 21573
rect 6454 21564 6460 21616
rect 6512 21604 6518 21616
rect 10594 21604 10600 21616
rect 6512 21576 10600 21604
rect 6512 21564 6518 21576
rect 10594 21564 10600 21576
rect 10652 21564 10658 21616
rect 10686 21564 10692 21616
rect 10744 21604 10750 21616
rect 13906 21604 13912 21616
rect 10744 21576 13912 21604
rect 10744 21564 10750 21576
rect 13906 21564 13912 21576
rect 13964 21564 13970 21616
rect 14090 21604 14096 21616
rect 14051 21576 14096 21604
rect 14090 21564 14096 21576
rect 14148 21564 14154 21616
rect 1578 21496 1584 21548
rect 1636 21536 1642 21548
rect 1673 21539 1731 21545
rect 1673 21536 1685 21539
rect 1636 21508 1685 21536
rect 1636 21496 1642 21508
rect 1673 21505 1685 21508
rect 1719 21505 1731 21539
rect 1673 21499 1731 21505
rect 1857 21539 1915 21545
rect 1857 21505 1869 21539
rect 1903 21536 1915 21539
rect 5718 21536 5724 21548
rect 1903 21508 5724 21536
rect 1903 21505 1915 21508
rect 1857 21499 1915 21505
rect 5718 21496 5724 21508
rect 5776 21496 5782 21548
rect 10502 21536 10508 21548
rect 10463 21508 10508 21536
rect 10502 21496 10508 21508
rect 10560 21496 10566 21548
rect 13262 21536 13268 21548
rect 10612 21508 13268 21536
rect 9493 21471 9551 21477
rect 9493 21437 9505 21471
rect 9539 21468 9551 21471
rect 10226 21468 10232 21480
rect 9539 21440 10232 21468
rect 9539 21437 9551 21440
rect 9493 21431 9551 21437
rect 10226 21428 10232 21440
rect 10284 21468 10290 21480
rect 10612 21468 10640 21508
rect 13262 21496 13268 21508
rect 13320 21536 13326 21548
rect 13449 21539 13507 21545
rect 13449 21536 13461 21539
rect 13320 21508 13461 21536
rect 13320 21496 13326 21508
rect 13449 21505 13461 21508
rect 13495 21505 13507 21539
rect 13449 21499 13507 21505
rect 14369 21539 14427 21545
rect 14369 21505 14381 21539
rect 14415 21536 14427 21539
rect 15286 21536 15292 21548
rect 14415 21508 15292 21536
rect 14415 21505 14427 21508
rect 14369 21499 14427 21505
rect 15286 21496 15292 21508
rect 15344 21496 15350 21548
rect 15654 21536 15660 21548
rect 15615 21508 15660 21536
rect 15654 21496 15660 21508
rect 15712 21496 15718 21548
rect 36814 21496 36820 21548
rect 36872 21536 36878 21548
rect 38013 21539 38071 21545
rect 38013 21536 38025 21539
rect 36872 21508 38025 21536
rect 36872 21496 36878 21508
rect 38013 21505 38025 21508
rect 38059 21505 38071 21539
rect 38013 21499 38071 21505
rect 10284 21440 10640 21468
rect 10689 21471 10747 21477
rect 10284 21428 10290 21440
rect 10689 21437 10701 21471
rect 10735 21468 10747 21471
rect 11054 21468 11060 21480
rect 10735 21440 11060 21468
rect 10735 21437 10747 21440
rect 10689 21431 10747 21437
rect 11054 21428 11060 21440
rect 11112 21428 11118 21480
rect 11606 21428 11612 21480
rect 11664 21468 11670 21480
rect 12621 21471 12679 21477
rect 12621 21468 12633 21471
rect 11664 21440 12633 21468
rect 11664 21428 11670 21440
rect 12621 21437 12633 21440
rect 12667 21437 12679 21471
rect 12802 21468 12808 21480
rect 12763 21440 12808 21468
rect 12621 21431 12679 21437
rect 12802 21428 12808 21440
rect 12860 21428 12866 21480
rect 15378 21428 15384 21480
rect 15436 21468 15442 21480
rect 15841 21471 15899 21477
rect 15841 21468 15853 21471
rect 15436 21440 15853 21468
rect 15436 21428 15442 21440
rect 15841 21437 15853 21440
rect 15887 21468 15899 21471
rect 16022 21468 16028 21480
rect 15887 21440 16028 21468
rect 15887 21437 15899 21440
rect 15841 21431 15899 21437
rect 16022 21428 16028 21440
rect 16080 21428 16086 21480
rect 16666 21428 16672 21480
rect 16724 21468 16730 21480
rect 17313 21471 17371 21477
rect 17313 21468 17325 21471
rect 16724 21440 17325 21468
rect 16724 21428 16730 21440
rect 17313 21437 17325 21440
rect 17359 21437 17371 21471
rect 17313 21431 17371 21437
rect 17497 21471 17555 21477
rect 17497 21437 17509 21471
rect 17543 21468 17555 21471
rect 17862 21468 17868 21480
rect 17543 21440 17868 21468
rect 17543 21437 17555 21440
rect 17497 21431 17555 21437
rect 17862 21428 17868 21440
rect 17920 21428 17926 21480
rect 15473 21403 15531 21409
rect 15473 21369 15485 21403
rect 15519 21400 15531 21403
rect 15562 21400 15568 21412
rect 15519 21372 15568 21400
rect 15519 21369 15531 21372
rect 15473 21363 15531 21369
rect 15562 21360 15568 21372
rect 15620 21400 15626 21412
rect 15620 21372 16574 21400
rect 15620 21360 15626 21372
rect 4433 21335 4491 21341
rect 4433 21301 4445 21335
rect 4479 21332 4491 21335
rect 4614 21332 4620 21344
rect 4479 21304 4620 21332
rect 4479 21301 4491 21304
rect 4433 21295 4491 21301
rect 4614 21292 4620 21304
rect 4672 21292 4678 21344
rect 10045 21335 10103 21341
rect 10045 21301 10057 21335
rect 10091 21332 10103 21335
rect 11238 21332 11244 21344
rect 10091 21304 11244 21332
rect 10091 21301 10103 21304
rect 10045 21295 10103 21301
rect 11238 21292 11244 21304
rect 11296 21292 11302 21344
rect 13541 21335 13599 21341
rect 13541 21301 13553 21335
rect 13587 21332 13599 21335
rect 15102 21332 15108 21344
rect 13587 21304 15108 21332
rect 13587 21301 13599 21304
rect 13541 21295 13599 21301
rect 15102 21292 15108 21304
rect 15160 21292 15166 21344
rect 16546 21332 16574 21372
rect 16853 21335 16911 21341
rect 16853 21332 16865 21335
rect 16546 21304 16865 21332
rect 16853 21301 16865 21304
rect 16899 21301 16911 21335
rect 38194 21332 38200 21344
rect 38155 21304 38200 21332
rect 16853 21295 16911 21301
rect 38194 21292 38200 21304
rect 38252 21292 38258 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 1578 21128 1584 21140
rect 1539 21100 1584 21128
rect 1578 21088 1584 21100
rect 1636 21088 1642 21140
rect 2590 21088 2596 21140
rect 2648 21128 2654 21140
rect 2866 21128 2872 21140
rect 2648 21100 2872 21128
rect 2648 21088 2654 21100
rect 2866 21088 2872 21100
rect 2924 21128 2930 21140
rect 3145 21131 3203 21137
rect 3145 21128 3157 21131
rect 2924 21100 3157 21128
rect 2924 21088 2930 21100
rect 3145 21097 3157 21100
rect 3191 21097 3203 21131
rect 3145 21091 3203 21097
rect 4065 21131 4123 21137
rect 4065 21097 4077 21131
rect 4111 21128 4123 21131
rect 4614 21128 4620 21140
rect 4111 21100 4620 21128
rect 4111 21097 4123 21100
rect 4065 21091 4123 21097
rect 4614 21088 4620 21100
rect 4672 21128 4678 21140
rect 5169 21131 5227 21137
rect 5169 21128 5181 21131
rect 4672 21100 5181 21128
rect 4672 21088 4678 21100
rect 5169 21097 5181 21100
rect 5215 21128 5227 21131
rect 5258 21128 5264 21140
rect 5215 21100 5264 21128
rect 5215 21097 5227 21100
rect 5169 21091 5227 21097
rect 5258 21088 5264 21100
rect 5316 21088 5322 21140
rect 11606 21128 11612 21140
rect 11567 21100 11612 21128
rect 11606 21088 11612 21100
rect 11664 21088 11670 21140
rect 16666 21128 16672 21140
rect 16627 21100 16672 21128
rect 16666 21088 16672 21100
rect 16724 21088 16730 21140
rect 17957 21131 18015 21137
rect 17957 21097 17969 21131
rect 18003 21128 18015 21131
rect 18046 21128 18052 21140
rect 18003 21100 18052 21128
rect 18003 21097 18015 21100
rect 17957 21091 18015 21097
rect 18046 21088 18052 21100
rect 18104 21088 18110 21140
rect 2682 21060 2688 21072
rect 2643 21032 2688 21060
rect 2682 21020 2688 21032
rect 2740 21020 2746 21072
rect 12437 21063 12495 21069
rect 12437 21029 12449 21063
rect 12483 21060 12495 21063
rect 26510 21060 26516 21072
rect 12483 21032 26516 21060
rect 12483 21029 12495 21032
rect 12437 21023 12495 21029
rect 26510 21020 26516 21032
rect 26568 21020 26574 21072
rect 10965 20995 11023 21001
rect 10965 20961 10977 20995
rect 11011 20992 11023 20995
rect 12802 20992 12808 21004
rect 11011 20964 12808 20992
rect 11011 20961 11023 20964
rect 10965 20955 11023 20961
rect 12802 20952 12808 20964
rect 12860 20992 12866 21004
rect 12897 20995 12955 21001
rect 12897 20992 12909 20995
rect 12860 20964 12909 20992
rect 12860 20952 12866 20964
rect 12897 20961 12909 20964
rect 12943 20961 12955 20995
rect 12897 20955 12955 20961
rect 13906 20952 13912 21004
rect 13964 20992 13970 21004
rect 14277 20995 14335 21001
rect 14277 20992 14289 20995
rect 13964 20964 14289 20992
rect 13964 20952 13970 20964
rect 14277 20961 14289 20964
rect 14323 20961 14335 20995
rect 14277 20955 14335 20961
rect 15470 20952 15476 21004
rect 15528 20992 15534 21004
rect 17313 20995 17371 21001
rect 17313 20992 17325 20995
rect 15528 20964 17325 20992
rect 15528 20952 15534 20964
rect 17313 20961 17325 20964
rect 17359 20961 17371 20995
rect 17313 20955 17371 20961
rect 10873 20927 10931 20933
rect 10873 20893 10885 20927
rect 10919 20924 10931 20927
rect 11238 20924 11244 20936
rect 10919 20896 11244 20924
rect 10919 20893 10931 20896
rect 10873 20887 10931 20893
rect 11238 20884 11244 20896
rect 11296 20884 11302 20936
rect 11514 20924 11520 20936
rect 11475 20896 11520 20924
rect 11514 20884 11520 20896
rect 11572 20884 11578 20936
rect 13078 20924 13084 20936
rect 13039 20896 13084 20924
rect 13078 20884 13084 20896
rect 13136 20884 13142 20936
rect 16577 20927 16635 20933
rect 16577 20893 16589 20927
rect 16623 20924 16635 20927
rect 16942 20924 16948 20936
rect 16623 20896 16948 20924
rect 16623 20893 16635 20896
rect 16577 20887 16635 20893
rect 16942 20884 16948 20896
rect 17000 20924 17006 20936
rect 17405 20927 17463 20933
rect 17405 20924 17417 20927
rect 17000 20896 17417 20924
rect 17000 20884 17006 20896
rect 17405 20893 17417 20896
rect 17451 20924 17463 20927
rect 18046 20924 18052 20936
rect 17451 20896 18052 20924
rect 17451 20893 17463 20896
rect 17405 20887 17463 20893
rect 18046 20884 18052 20896
rect 18104 20884 18110 20936
rect 12253 20859 12311 20865
rect 12253 20856 12265 20859
rect 10520 20828 12265 20856
rect 10520 20800 10548 20828
rect 12253 20825 12265 20828
rect 12299 20825 12311 20859
rect 14826 20856 14832 20868
rect 14787 20828 14832 20856
rect 12253 20819 12311 20825
rect 14826 20816 14832 20828
rect 14884 20816 14890 20868
rect 14921 20859 14979 20865
rect 14921 20825 14933 20859
rect 14967 20856 14979 20859
rect 15378 20856 15384 20868
rect 14967 20828 15384 20856
rect 14967 20825 14979 20828
rect 14921 20819 14979 20825
rect 15378 20816 15384 20828
rect 15436 20816 15442 20868
rect 15657 20859 15715 20865
rect 15657 20825 15669 20859
rect 15703 20856 15715 20859
rect 16666 20856 16672 20868
rect 15703 20828 16672 20856
rect 15703 20825 15715 20828
rect 15657 20819 15715 20825
rect 16666 20816 16672 20828
rect 16724 20856 16730 20868
rect 20806 20856 20812 20868
rect 16724 20828 20812 20856
rect 16724 20816 16730 20828
rect 20806 20816 20812 20828
rect 20864 20816 20870 20868
rect 4890 20748 4896 20800
rect 4948 20788 4954 20800
rect 5629 20791 5687 20797
rect 5629 20788 5641 20791
rect 4948 20760 5641 20788
rect 4948 20748 4954 20760
rect 5629 20757 5641 20760
rect 5675 20757 5687 20791
rect 5629 20751 5687 20757
rect 10413 20791 10471 20797
rect 10413 20757 10425 20791
rect 10459 20788 10471 20791
rect 10502 20788 10508 20800
rect 10459 20760 10508 20788
rect 10459 20757 10471 20760
rect 10413 20751 10471 20757
rect 10502 20748 10508 20760
rect 10560 20748 10566 20800
rect 12066 20748 12072 20800
rect 12124 20788 12130 20800
rect 12710 20788 12716 20800
rect 12124 20760 12716 20788
rect 12124 20748 12130 20760
rect 12710 20748 12716 20760
rect 12768 20748 12774 20800
rect 13538 20788 13544 20800
rect 13499 20760 13544 20788
rect 13538 20748 13544 20760
rect 13596 20748 13602 20800
rect 15562 20788 15568 20800
rect 15523 20760 15568 20788
rect 15562 20748 15568 20760
rect 15620 20748 15626 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 1578 20584 1584 20596
rect 1539 20556 1584 20584
rect 1578 20544 1584 20556
rect 1636 20544 1642 20596
rect 2225 20587 2283 20593
rect 2225 20553 2237 20587
rect 2271 20584 2283 20587
rect 2958 20584 2964 20596
rect 2271 20556 2964 20584
rect 2271 20553 2283 20556
rect 2225 20547 2283 20553
rect 2958 20544 2964 20556
rect 3016 20544 3022 20596
rect 3605 20587 3663 20593
rect 3605 20553 3617 20587
rect 3651 20584 3663 20587
rect 4062 20584 4068 20596
rect 3651 20556 4068 20584
rect 3651 20553 3663 20556
rect 3605 20547 3663 20553
rect 4062 20544 4068 20556
rect 4120 20584 4126 20596
rect 4157 20587 4215 20593
rect 4157 20584 4169 20587
rect 4120 20556 4169 20584
rect 4120 20544 4126 20556
rect 4157 20553 4169 20556
rect 4203 20584 4215 20587
rect 5258 20584 5264 20596
rect 4203 20556 5264 20584
rect 4203 20553 4215 20556
rect 4157 20547 4215 20553
rect 5258 20544 5264 20556
rect 5316 20544 5322 20596
rect 10318 20544 10324 20596
rect 10376 20584 10382 20596
rect 10413 20587 10471 20593
rect 10413 20584 10425 20587
rect 10376 20556 10425 20584
rect 10376 20544 10382 20556
rect 10413 20553 10425 20556
rect 10459 20553 10471 20587
rect 11054 20584 11060 20596
rect 11015 20556 11060 20584
rect 10413 20547 10471 20553
rect 11054 20544 11060 20556
rect 11112 20544 11118 20596
rect 11514 20544 11520 20596
rect 11572 20584 11578 20596
rect 12342 20584 12348 20596
rect 11572 20556 12348 20584
rect 11572 20544 11578 20556
rect 12342 20544 12348 20556
rect 12400 20584 12406 20596
rect 13173 20587 13231 20593
rect 12400 20556 13124 20584
rect 12400 20544 12406 20556
rect 2774 20516 2780 20528
rect 2687 20488 2780 20516
rect 2774 20476 2780 20488
rect 2832 20516 2838 20528
rect 3878 20516 3884 20528
rect 2832 20488 3884 20516
rect 2832 20476 2838 20488
rect 3878 20476 3884 20488
rect 3936 20476 3942 20528
rect 4709 20519 4767 20525
rect 4709 20485 4721 20519
rect 4755 20516 4767 20519
rect 4890 20516 4896 20528
rect 4755 20488 4896 20516
rect 4755 20485 4767 20488
rect 4709 20479 4767 20485
rect 4890 20476 4896 20488
rect 4948 20476 4954 20528
rect 6270 20476 6276 20528
rect 6328 20516 6334 20528
rect 12253 20519 12311 20525
rect 12253 20516 12265 20519
rect 6328 20488 12265 20516
rect 6328 20476 6334 20488
rect 12253 20485 12265 20488
rect 12299 20485 12311 20519
rect 12253 20479 12311 20485
rect 9861 20451 9919 20457
rect 9861 20417 9873 20451
rect 9907 20448 9919 20451
rect 10502 20448 10508 20460
rect 9907 20420 10508 20448
rect 9907 20417 9919 20420
rect 9861 20411 9919 20417
rect 10502 20408 10508 20420
rect 10560 20408 10566 20460
rect 10594 20408 10600 20460
rect 10652 20448 10658 20460
rect 13096 20457 13124 20556
rect 13173 20553 13185 20587
rect 13219 20584 13231 20587
rect 14826 20584 14832 20596
rect 13219 20556 14832 20584
rect 13219 20553 13231 20556
rect 13173 20547 13231 20553
rect 14826 20544 14832 20556
rect 14884 20544 14890 20596
rect 16942 20584 16948 20596
rect 16903 20556 16948 20584
rect 16942 20544 16948 20556
rect 17000 20544 17006 20596
rect 13817 20519 13875 20525
rect 13817 20485 13829 20519
rect 13863 20516 13875 20519
rect 16025 20519 16083 20525
rect 16025 20516 16037 20519
rect 13863 20488 16037 20516
rect 13863 20485 13875 20488
rect 13817 20479 13875 20485
rect 16025 20485 16037 20488
rect 16071 20485 16083 20519
rect 16025 20479 16083 20485
rect 16117 20519 16175 20525
rect 16117 20485 16129 20519
rect 16163 20516 16175 20519
rect 17862 20516 17868 20528
rect 16163 20488 17868 20516
rect 16163 20485 16175 20488
rect 16117 20479 16175 20485
rect 17862 20476 17868 20488
rect 17920 20476 17926 20528
rect 11149 20451 11207 20457
rect 11149 20448 11161 20451
rect 10652 20420 11161 20448
rect 10652 20408 10658 20420
rect 11149 20417 11161 20420
rect 11195 20417 11207 20451
rect 11149 20411 11207 20417
rect 13081 20451 13139 20457
rect 13081 20417 13093 20451
rect 13127 20417 13139 20451
rect 13725 20451 13783 20457
rect 13725 20448 13737 20451
rect 13081 20411 13139 20417
rect 13188 20420 13737 20448
rect 10318 20340 10324 20392
rect 10376 20380 10382 20392
rect 11701 20383 11759 20389
rect 11701 20380 11713 20383
rect 10376 20352 11713 20380
rect 10376 20340 10382 20352
rect 11701 20349 11713 20352
rect 11747 20349 11759 20383
rect 11701 20343 11759 20349
rect 12158 20340 12164 20392
rect 12216 20380 12222 20392
rect 12345 20383 12403 20389
rect 12345 20380 12357 20383
rect 12216 20352 12357 20380
rect 12216 20340 12222 20352
rect 12345 20349 12357 20352
rect 12391 20349 12403 20383
rect 13188 20380 13216 20420
rect 13725 20417 13737 20420
rect 13771 20417 13783 20451
rect 13725 20411 13783 20417
rect 14829 20451 14887 20457
rect 14829 20417 14841 20451
rect 14875 20448 14887 20451
rect 15470 20448 15476 20460
rect 14875 20420 15476 20448
rect 14875 20417 14887 20420
rect 14829 20411 14887 20417
rect 15470 20408 15476 20420
rect 15528 20408 15534 20460
rect 12345 20343 12403 20349
rect 12452 20352 13216 20380
rect 12452 20324 12480 20352
rect 13538 20340 13544 20392
rect 13596 20380 13602 20392
rect 14369 20383 14427 20389
rect 14369 20380 14381 20383
rect 13596 20352 14381 20380
rect 13596 20340 13602 20352
rect 14369 20349 14381 20352
rect 14415 20349 14427 20383
rect 15010 20380 15016 20392
rect 14971 20352 15016 20380
rect 14369 20343 14427 20349
rect 15010 20340 15016 20352
rect 15068 20340 15074 20392
rect 12434 20272 12440 20324
rect 12492 20272 12498 20324
rect 13906 20272 13912 20324
rect 13964 20312 13970 20324
rect 14826 20312 14832 20324
rect 13964 20284 14832 20312
rect 13964 20272 13970 20284
rect 14826 20272 14832 20284
rect 14884 20312 14890 20324
rect 15565 20315 15623 20321
rect 15565 20312 15577 20315
rect 14884 20284 15577 20312
rect 14884 20272 14890 20284
rect 15565 20281 15577 20284
rect 15611 20281 15623 20315
rect 15565 20275 15623 20281
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 1670 20040 1676 20052
rect 1631 20012 1676 20040
rect 1670 20000 1676 20012
rect 1728 20000 1734 20052
rect 2130 20000 2136 20052
rect 2188 20040 2194 20052
rect 2225 20043 2283 20049
rect 2225 20040 2237 20043
rect 2188 20012 2237 20040
rect 2188 20000 2194 20012
rect 2225 20009 2237 20012
rect 2271 20009 2283 20043
rect 2866 20040 2872 20052
rect 2827 20012 2872 20040
rect 2225 20003 2283 20009
rect 2866 20000 2872 20012
rect 2924 20040 2930 20052
rect 3142 20040 3148 20052
rect 2924 20012 3148 20040
rect 2924 20000 2930 20012
rect 3142 20000 3148 20012
rect 3200 20000 3206 20052
rect 3326 20040 3332 20052
rect 3287 20012 3332 20040
rect 3326 20000 3332 20012
rect 3384 20000 3390 20052
rect 4062 20040 4068 20052
rect 4023 20012 4068 20040
rect 4062 20000 4068 20012
rect 4120 20000 4126 20052
rect 10870 20000 10876 20052
rect 10928 20040 10934 20052
rect 12253 20043 12311 20049
rect 12253 20040 12265 20043
rect 10928 20012 12265 20040
rect 10928 20000 10934 20012
rect 12253 20009 12265 20012
rect 12299 20009 12311 20043
rect 12253 20003 12311 20009
rect 12526 20000 12532 20052
rect 12584 20040 12590 20052
rect 12989 20043 13047 20049
rect 12989 20040 13001 20043
rect 12584 20012 13001 20040
rect 12584 20000 12590 20012
rect 12989 20009 13001 20012
rect 13035 20009 13047 20043
rect 12989 20003 13047 20009
rect 13078 20000 13084 20052
rect 13136 20040 13142 20052
rect 13633 20043 13691 20049
rect 13633 20040 13645 20043
rect 13136 20012 13645 20040
rect 13136 20000 13142 20012
rect 13633 20009 13645 20012
rect 13679 20009 13691 20043
rect 16666 20040 16672 20052
rect 16627 20012 16672 20040
rect 13633 20003 13691 20009
rect 16666 20000 16672 20012
rect 16724 20000 16730 20052
rect 12342 19932 12348 19984
rect 12400 19932 12406 19984
rect 12360 19904 12388 19932
rect 12360 19876 13124 19904
rect 12345 19839 12403 19845
rect 12345 19805 12357 19839
rect 12391 19836 12403 19839
rect 12434 19836 12440 19848
rect 12391 19808 12440 19836
rect 12391 19805 12403 19808
rect 12345 19799 12403 19805
rect 12434 19796 12440 19808
rect 12492 19796 12498 19848
rect 13096 19845 13124 19876
rect 14826 19864 14832 19916
rect 14884 19904 14890 19916
rect 15381 19907 15439 19913
rect 15381 19904 15393 19907
rect 14884 19876 15393 19904
rect 14884 19864 14890 19876
rect 15381 19873 15393 19876
rect 15427 19873 15439 19907
rect 15381 19867 15439 19873
rect 16025 19907 16083 19913
rect 16025 19873 16037 19907
rect 16071 19904 16083 19907
rect 16574 19904 16580 19916
rect 16071 19876 16580 19904
rect 16071 19873 16083 19876
rect 16025 19867 16083 19873
rect 16574 19864 16580 19876
rect 16632 19864 16638 19916
rect 38013 19907 38071 19913
rect 38013 19873 38025 19907
rect 38059 19904 38071 19907
rect 38102 19904 38108 19916
rect 38059 19876 38108 19904
rect 38059 19873 38071 19876
rect 38013 19867 38071 19873
rect 38102 19864 38108 19876
rect 38160 19864 38166 19916
rect 13081 19839 13139 19845
rect 13081 19805 13093 19839
rect 13127 19805 13139 19839
rect 13081 19799 13139 19805
rect 13725 19839 13783 19845
rect 13725 19805 13737 19839
rect 13771 19805 13783 19839
rect 13725 19799 13783 19805
rect 14461 19839 14519 19845
rect 14461 19805 14473 19839
rect 14507 19836 14519 19839
rect 14734 19836 14740 19848
rect 14507 19808 14740 19836
rect 14507 19805 14519 19808
rect 14461 19799 14519 19805
rect 3326 19728 3332 19780
rect 3384 19768 3390 19780
rect 10962 19768 10968 19780
rect 3384 19740 10968 19768
rect 3384 19728 3390 19740
rect 10962 19728 10968 19740
rect 11020 19728 11026 19780
rect 12710 19728 12716 19780
rect 12768 19768 12774 19780
rect 13740 19768 13768 19799
rect 14734 19796 14740 19808
rect 14792 19796 14798 19848
rect 38286 19836 38292 19848
rect 38247 19808 38292 19836
rect 38286 19796 38292 19808
rect 38344 19796 38350 19848
rect 12768 19740 13768 19768
rect 15933 19771 15991 19777
rect 12768 19728 12774 19740
rect 15933 19737 15945 19771
rect 15979 19737 15991 19771
rect 15933 19731 15991 19737
rect 6178 19660 6184 19712
rect 6236 19700 6242 19712
rect 10594 19700 10600 19712
rect 6236 19672 10600 19700
rect 6236 19660 6242 19672
rect 10594 19660 10600 19672
rect 10652 19660 10658 19712
rect 11238 19700 11244 19712
rect 11199 19672 11244 19700
rect 11238 19660 11244 19672
rect 11296 19660 11302 19712
rect 14274 19700 14280 19712
rect 14235 19672 14280 19700
rect 14274 19660 14280 19672
rect 14332 19660 14338 19712
rect 15102 19660 15108 19712
rect 15160 19700 15166 19712
rect 15948 19700 15976 19731
rect 15160 19672 15976 19700
rect 15160 19660 15166 19672
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 10594 19456 10600 19508
rect 10652 19496 10658 19508
rect 11977 19499 12035 19505
rect 11977 19496 11989 19499
rect 10652 19468 11989 19496
rect 10652 19456 10658 19468
rect 11977 19465 11989 19468
rect 12023 19496 12035 19499
rect 12434 19496 12440 19508
rect 12023 19468 12440 19496
rect 12023 19465 12035 19468
rect 11977 19459 12035 19465
rect 12434 19456 12440 19468
rect 12492 19456 12498 19508
rect 12710 19496 12716 19508
rect 12671 19468 12716 19496
rect 12710 19456 12716 19468
rect 12768 19456 12774 19508
rect 14737 19499 14795 19505
rect 14737 19465 14749 19499
rect 14783 19496 14795 19499
rect 15010 19496 15016 19508
rect 14783 19468 15016 19496
rect 14783 19465 14795 19468
rect 14737 19459 14795 19465
rect 15010 19456 15016 19468
rect 15068 19456 15074 19508
rect 28534 19496 28540 19508
rect 16546 19468 28540 19496
rect 11238 19388 11244 19440
rect 11296 19428 11302 19440
rect 16546 19428 16574 19468
rect 28534 19456 28540 19468
rect 28592 19456 28598 19508
rect 38286 19496 38292 19508
rect 38247 19468 38292 19496
rect 38286 19456 38292 19468
rect 38344 19456 38350 19508
rect 11296 19400 16574 19428
rect 11296 19388 11302 19400
rect 1578 19320 1584 19372
rect 1636 19360 1642 19372
rect 1673 19363 1731 19369
rect 1673 19360 1685 19363
rect 1636 19332 1685 19360
rect 1636 19320 1642 19332
rect 1673 19329 1685 19332
rect 1719 19329 1731 19363
rect 1673 19323 1731 19329
rect 14734 19320 14740 19372
rect 14792 19360 14798 19372
rect 14792 19332 15240 19360
rect 14792 19320 14798 19332
rect 15212 19304 15240 19332
rect 2314 19292 2320 19304
rect 2275 19264 2320 19292
rect 2314 19252 2320 19264
rect 2372 19252 2378 19304
rect 13262 19292 13268 19304
rect 13223 19264 13268 19292
rect 13262 19252 13268 19264
rect 13320 19252 13326 19304
rect 15194 19292 15200 19304
rect 15107 19264 15200 19292
rect 15194 19252 15200 19264
rect 15252 19252 15258 19304
rect 1857 19227 1915 19233
rect 1857 19193 1869 19227
rect 1903 19224 1915 19227
rect 14001 19227 14059 19233
rect 14001 19224 14013 19227
rect 1903 19196 14013 19224
rect 1903 19193 1915 19196
rect 1857 19187 1915 19193
rect 14001 19193 14013 19196
rect 14047 19224 14059 19227
rect 15286 19224 15292 19236
rect 14047 19196 15292 19224
rect 14047 19193 14059 19196
rect 14001 19187 14059 19193
rect 15286 19184 15292 19196
rect 15344 19224 15350 19236
rect 16022 19224 16028 19236
rect 15344 19196 16028 19224
rect 15344 19184 15350 19196
rect 16022 19184 16028 19196
rect 16080 19184 16086 19236
rect 1026 19116 1032 19168
rect 1084 19156 1090 19168
rect 2869 19159 2927 19165
rect 2869 19156 2881 19159
rect 1084 19128 2881 19156
rect 1084 19116 1090 19128
rect 2869 19125 2881 19128
rect 2915 19125 2927 19159
rect 2869 19119 2927 19125
rect 16301 19159 16359 19165
rect 16301 19125 16313 19159
rect 16347 19156 16359 19159
rect 16574 19156 16580 19168
rect 16347 19128 16580 19156
rect 16347 19125 16359 19128
rect 16301 19119 16359 19125
rect 16574 19116 16580 19128
rect 16632 19156 16638 19168
rect 17770 19156 17776 19168
rect 16632 19128 17776 19156
rect 16632 19116 16638 19128
rect 17770 19116 17776 19128
rect 17828 19116 17834 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 1578 18952 1584 18964
rect 1539 18924 1584 18952
rect 1578 18912 1584 18924
rect 1636 18912 1642 18964
rect 2222 18952 2228 18964
rect 2183 18924 2228 18952
rect 2222 18912 2228 18924
rect 2280 18912 2286 18964
rect 4985 18955 5043 18961
rect 4985 18921 4997 18955
rect 5031 18952 5043 18955
rect 5166 18952 5172 18964
rect 5031 18924 5172 18952
rect 5031 18921 5043 18924
rect 4985 18915 5043 18921
rect 4433 18751 4491 18757
rect 4433 18717 4445 18751
rect 4479 18748 4491 18751
rect 5000 18748 5028 18915
rect 5166 18912 5172 18924
rect 5224 18912 5230 18964
rect 12434 18912 12440 18964
rect 12492 18952 12498 18964
rect 13541 18955 13599 18961
rect 13541 18952 13553 18955
rect 12492 18924 13553 18952
rect 12492 18912 12498 18924
rect 13541 18921 13553 18924
rect 13587 18921 13599 18955
rect 13541 18915 13599 18921
rect 19426 18912 19432 18964
rect 19484 18952 19490 18964
rect 19521 18955 19579 18961
rect 19521 18952 19533 18955
rect 19484 18924 19533 18952
rect 19484 18912 19490 18924
rect 19521 18921 19533 18924
rect 19567 18921 19579 18955
rect 19521 18915 19579 18921
rect 4479 18720 5028 18748
rect 19613 18751 19671 18757
rect 4479 18717 4491 18720
rect 4433 18711 4491 18717
rect 19613 18717 19625 18751
rect 19659 18748 19671 18751
rect 19659 18720 20208 18748
rect 19659 18717 19671 18720
rect 19613 18711 19671 18717
rect 2774 18572 2780 18624
rect 2832 18612 2838 18624
rect 20180 18621 20208 18720
rect 4249 18615 4307 18621
rect 4249 18612 4261 18615
rect 2832 18584 4261 18612
rect 2832 18572 2838 18584
rect 4249 18581 4261 18584
rect 4295 18581 4307 18615
rect 4249 18575 4307 18581
rect 20165 18615 20223 18621
rect 20165 18581 20177 18615
rect 20211 18612 20223 18615
rect 22370 18612 22376 18624
rect 20211 18584 22376 18612
rect 20211 18581 20223 18584
rect 20165 18575 20223 18581
rect 22370 18572 22376 18584
rect 22428 18572 22434 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 1857 18275 1915 18281
rect 1857 18241 1869 18275
rect 1903 18272 1915 18275
rect 14274 18272 14280 18284
rect 1903 18244 14280 18272
rect 1903 18241 1915 18244
rect 1857 18235 1915 18241
rect 14274 18232 14280 18244
rect 14332 18232 14338 18284
rect 29457 18275 29515 18281
rect 29457 18241 29469 18275
rect 29503 18272 29515 18275
rect 38010 18272 38016 18284
rect 29503 18244 38016 18272
rect 29503 18241 29515 18244
rect 29457 18235 29515 18241
rect 38010 18232 38016 18244
rect 38068 18232 38074 18284
rect 1670 18068 1676 18080
rect 1631 18040 1676 18068
rect 1670 18028 1676 18040
rect 1728 18028 1734 18080
rect 17770 18028 17776 18080
rect 17828 18068 17834 18080
rect 29365 18071 29423 18077
rect 29365 18068 29377 18071
rect 17828 18040 29377 18068
rect 17828 18028 17834 18040
rect 29365 18037 29377 18040
rect 29411 18037 29423 18071
rect 29365 18031 29423 18037
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 17862 17280 17868 17332
rect 17920 17320 17926 17332
rect 19797 17323 19855 17329
rect 19797 17320 19809 17323
rect 17920 17292 19809 17320
rect 17920 17280 17926 17292
rect 19797 17289 19809 17292
rect 19843 17289 19855 17323
rect 19797 17283 19855 17289
rect 6825 17187 6883 17193
rect 6825 17153 6837 17187
rect 6871 17184 6883 17187
rect 7558 17184 7564 17196
rect 6871 17156 7564 17184
rect 6871 17153 6883 17156
rect 6825 17147 6883 17153
rect 7558 17144 7564 17156
rect 7616 17144 7622 17196
rect 19889 17187 19947 17193
rect 19889 17153 19901 17187
rect 19935 17184 19947 17187
rect 19935 17156 20484 17184
rect 19935 17153 19947 17156
rect 19889 17147 19947 17153
rect 6730 16980 6736 16992
rect 6691 16952 6736 16980
rect 6730 16940 6736 16952
rect 6788 16940 6794 16992
rect 20456 16989 20484 17156
rect 20441 16983 20499 16989
rect 20441 16949 20453 16983
rect 20487 16980 20499 16983
rect 24394 16980 24400 16992
rect 20487 16952 24400 16980
rect 20487 16949 20499 16952
rect 20441 16943 20499 16949
rect 24394 16940 24400 16952
rect 24452 16940 24458 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 1857 16099 1915 16105
rect 1857 16065 1869 16099
rect 1903 16096 1915 16099
rect 2774 16096 2780 16108
rect 1903 16068 2780 16096
rect 1903 16065 1915 16068
rect 1857 16059 1915 16065
rect 2774 16056 2780 16068
rect 2832 16056 2838 16108
rect 37642 16056 37648 16108
rect 37700 16096 37706 16108
rect 38013 16099 38071 16105
rect 38013 16096 38025 16099
rect 37700 16068 38025 16096
rect 37700 16056 37706 16068
rect 38013 16065 38025 16068
rect 38059 16065 38071 16099
rect 38013 16059 38071 16065
rect 38286 16028 38292 16040
rect 38247 16000 38292 16028
rect 38286 15988 38292 16000
rect 38344 15988 38350 16040
rect 1670 15892 1676 15904
rect 1631 15864 1676 15892
rect 1670 15852 1676 15864
rect 1728 15852 1734 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 38286 15688 38292 15700
rect 38247 15660 38292 15688
rect 38286 15648 38292 15660
rect 38344 15648 38350 15700
rect 7101 15487 7159 15493
rect 7101 15453 7113 15487
rect 7147 15484 7159 15487
rect 10042 15484 10048 15496
rect 7147 15456 10048 15484
rect 7147 15453 7159 15456
rect 7101 15447 7159 15453
rect 10042 15444 10048 15456
rect 10100 15444 10106 15496
rect 6822 15308 6828 15360
rect 6880 15348 6886 15360
rect 7009 15351 7067 15357
rect 7009 15348 7021 15351
rect 6880 15320 7021 15348
rect 6880 15308 6886 15320
rect 7009 15317 7021 15320
rect 7055 15317 7067 15351
rect 7009 15311 7067 15317
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 2501 14603 2559 14609
rect 2501 14569 2513 14603
rect 2547 14600 2559 14603
rect 4798 14600 4804 14612
rect 2547 14572 4804 14600
rect 2547 14569 2559 14572
rect 2501 14563 2559 14569
rect 1949 14399 2007 14405
rect 1949 14365 1961 14399
rect 1995 14396 2007 14399
rect 2516 14396 2544 14563
rect 4798 14560 4804 14572
rect 4856 14560 4862 14612
rect 38010 14464 38016 14476
rect 37971 14436 38016 14464
rect 38010 14424 38016 14436
rect 38068 14424 38074 14476
rect 38286 14396 38292 14408
rect 1995 14368 2544 14396
rect 38247 14368 38292 14396
rect 1995 14365 2007 14368
rect 1949 14359 2007 14365
rect 38286 14356 38292 14368
rect 38344 14356 38350 14408
rect 1765 14263 1823 14269
rect 1765 14229 1777 14263
rect 1811 14260 1823 14263
rect 1946 14260 1952 14272
rect 1811 14232 1952 14260
rect 1811 14229 1823 14232
rect 1765 14223 1823 14229
rect 1946 14220 1952 14232
rect 2004 14220 2010 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 38286 14056 38292 14068
rect 38247 14028 38292 14056
rect 38286 14016 38292 14028
rect 38344 14016 38350 14068
rect 1857 13991 1915 13997
rect 1857 13957 1869 13991
rect 1903 13988 1915 13991
rect 4706 13988 4712 14000
rect 1903 13960 4712 13988
rect 1903 13957 1915 13960
rect 1857 13951 1915 13957
rect 4706 13948 4712 13960
rect 4764 13948 4770 14000
rect 1578 13880 1584 13932
rect 1636 13920 1642 13932
rect 1673 13923 1731 13929
rect 1673 13920 1685 13923
rect 1636 13892 1685 13920
rect 1636 13880 1642 13892
rect 1673 13889 1685 13892
rect 1719 13889 1731 13923
rect 1673 13883 1731 13889
rect 2501 13923 2559 13929
rect 2501 13889 2513 13923
rect 2547 13920 2559 13923
rect 10318 13920 10324 13932
rect 2547 13892 10324 13920
rect 2547 13889 2559 13892
rect 2501 13883 2559 13889
rect 10318 13880 10324 13892
rect 10376 13880 10382 13932
rect 2406 13852 2412 13864
rect 2367 13824 2412 13852
rect 2406 13812 2412 13824
rect 2464 13812 2470 13864
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 1578 13512 1584 13524
rect 1539 13484 1584 13512
rect 1578 13472 1584 13484
rect 1636 13472 1642 13524
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 1857 12835 1915 12841
rect 1857 12801 1869 12835
rect 1903 12832 1915 12835
rect 6730 12832 6736 12844
rect 1903 12804 6736 12832
rect 1903 12801 1915 12804
rect 1857 12795 1915 12801
rect 6730 12792 6736 12804
rect 6788 12792 6794 12844
rect 37553 12835 37611 12841
rect 37553 12801 37565 12835
rect 37599 12832 37611 12835
rect 38194 12832 38200 12844
rect 37599 12804 38200 12832
rect 37599 12801 37611 12804
rect 37553 12795 37611 12801
rect 38194 12792 38200 12804
rect 38252 12792 38258 12844
rect 37274 12656 37280 12708
rect 37332 12696 37338 12708
rect 38013 12699 38071 12705
rect 38013 12696 38025 12699
rect 37332 12668 38025 12696
rect 37332 12656 37338 12668
rect 38013 12665 38025 12668
rect 38059 12665 38071 12699
rect 38013 12659 38071 12665
rect 1670 12628 1676 12640
rect 1631 12600 1676 12628
rect 1670 12588 1676 12600
rect 1728 12588 1734 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 15378 12384 15384 12436
rect 15436 12424 15442 12436
rect 15565 12427 15623 12433
rect 15565 12424 15577 12427
rect 15436 12396 15577 12424
rect 15436 12384 15442 12396
rect 15565 12393 15577 12396
rect 15611 12393 15623 12427
rect 15565 12387 15623 12393
rect 15657 12223 15715 12229
rect 15657 12189 15669 12223
rect 15703 12220 15715 12223
rect 37829 12223 37887 12229
rect 15703 12192 16160 12220
rect 15703 12189 15715 12192
rect 15657 12183 15715 12189
rect 16132 12096 16160 12192
rect 37829 12189 37841 12223
rect 37875 12220 37887 12223
rect 38010 12220 38016 12232
rect 37875 12192 38016 12220
rect 37875 12189 37887 12192
rect 37829 12183 37887 12189
rect 38010 12180 38016 12192
rect 38068 12180 38074 12232
rect 16114 12084 16120 12096
rect 16075 12056 16120 12084
rect 16114 12044 16120 12056
rect 16172 12044 16178 12096
rect 38010 12084 38016 12096
rect 37971 12056 38016 12084
rect 38010 12044 38016 12056
rect 38068 12044 38074 12096
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 8386 11092 8392 11144
rect 8444 11132 8450 11144
rect 10781 11135 10839 11141
rect 10781 11132 10793 11135
rect 8444 11104 10793 11132
rect 8444 11092 8450 11104
rect 10781 11101 10793 11104
rect 10827 11132 10839 11135
rect 11425 11135 11483 11141
rect 11425 11132 11437 11135
rect 10827 11104 11437 11132
rect 10827 11101 10839 11104
rect 10781 11095 10839 11101
rect 11425 11101 11437 11104
rect 11471 11101 11483 11135
rect 11425 11095 11483 11101
rect 37826 11092 37832 11144
rect 37884 11132 37890 11144
rect 38013 11135 38071 11141
rect 38013 11132 38025 11135
rect 37884 11104 38025 11132
rect 37884 11092 37890 11104
rect 38013 11101 38025 11104
rect 38059 11101 38071 11135
rect 38013 11095 38071 11101
rect 10870 11064 10876 11076
rect 10831 11036 10876 11064
rect 10870 11024 10876 11036
rect 10928 11024 10934 11076
rect 37553 11067 37611 11073
rect 37553 11033 37565 11067
rect 37599 11064 37611 11067
rect 38194 11064 38200 11076
rect 37599 11036 38200 11064
rect 37599 11033 37611 11036
rect 37553 11027 37611 11033
rect 38194 11024 38200 11036
rect 38252 11024 38258 11076
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 8938 10792 8944 10804
rect 8899 10764 8944 10792
rect 8938 10752 8944 10764
rect 8996 10752 9002 10804
rect 11793 10795 11851 10801
rect 11793 10761 11805 10795
rect 11839 10792 11851 10795
rect 12618 10792 12624 10804
rect 11839 10764 12624 10792
rect 11839 10761 11851 10764
rect 11793 10755 11851 10761
rect 12618 10752 12624 10764
rect 12676 10752 12682 10804
rect 19978 10752 19984 10804
rect 20036 10792 20042 10804
rect 25409 10795 25467 10801
rect 25409 10792 25421 10795
rect 20036 10764 25421 10792
rect 20036 10752 20042 10764
rect 25409 10761 25421 10764
rect 25455 10761 25467 10795
rect 25409 10755 25467 10761
rect 1857 10659 1915 10665
rect 1857 10625 1869 10659
rect 1903 10656 1915 10659
rect 2406 10656 2412 10668
rect 1903 10628 2412 10656
rect 1903 10625 1915 10628
rect 1857 10619 1915 10625
rect 2406 10616 2412 10628
rect 2464 10616 2470 10668
rect 8662 10616 8668 10668
rect 8720 10656 8726 10668
rect 8849 10659 8907 10665
rect 8849 10656 8861 10659
rect 8720 10628 8861 10656
rect 8720 10616 8726 10628
rect 8849 10625 8861 10628
rect 8895 10625 8907 10659
rect 8849 10619 8907 10625
rect 11885 10659 11943 10665
rect 11885 10625 11897 10659
rect 11931 10656 11943 10659
rect 11931 10628 12480 10656
rect 11931 10625 11943 10628
rect 11885 10619 11943 10625
rect 1670 10452 1676 10464
rect 1631 10424 1676 10452
rect 1670 10412 1676 10424
rect 1728 10412 1734 10464
rect 12452 10461 12480 10628
rect 14366 10616 14372 10668
rect 14424 10656 14430 10668
rect 18969 10659 19027 10665
rect 18969 10656 18981 10659
rect 14424 10628 18981 10656
rect 14424 10616 14430 10628
rect 18969 10625 18981 10628
rect 19015 10656 19027 10659
rect 19613 10659 19671 10665
rect 19613 10656 19625 10659
rect 19015 10628 19625 10656
rect 19015 10625 19027 10628
rect 18969 10619 19027 10625
rect 19613 10625 19625 10628
rect 19659 10625 19671 10659
rect 19613 10619 19671 10625
rect 25501 10659 25559 10665
rect 25501 10625 25513 10659
rect 25547 10656 25559 10659
rect 25961 10659 26019 10665
rect 25961 10656 25973 10659
rect 25547 10628 25973 10656
rect 25547 10625 25559 10628
rect 25501 10619 25559 10625
rect 25961 10625 25973 10628
rect 26007 10656 26019 10659
rect 28994 10656 29000 10668
rect 26007 10628 29000 10656
rect 26007 10625 26019 10628
rect 25961 10619 26019 10625
rect 28994 10616 29000 10628
rect 29052 10616 29058 10668
rect 19061 10523 19119 10529
rect 19061 10489 19073 10523
rect 19107 10520 19119 10523
rect 22002 10520 22008 10532
rect 19107 10492 22008 10520
rect 19107 10489 19119 10492
rect 19061 10483 19119 10489
rect 22002 10480 22008 10492
rect 22060 10480 22066 10532
rect 12437 10455 12495 10461
rect 12437 10421 12449 10455
rect 12483 10452 12495 10455
rect 12710 10452 12716 10464
rect 12483 10424 12716 10452
rect 12483 10421 12495 10424
rect 12437 10415 12495 10421
rect 12710 10412 12716 10424
rect 12768 10412 12774 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 16850 10248 16856 10260
rect 16811 10220 16856 10248
rect 16850 10208 16856 10220
rect 16908 10208 16914 10260
rect 16117 10047 16175 10053
rect 16117 10013 16129 10047
rect 16163 10044 16175 10047
rect 16850 10044 16856 10056
rect 16163 10016 16856 10044
rect 16163 10013 16175 10016
rect 16117 10007 16175 10013
rect 16850 10004 16856 10016
rect 16908 10004 16914 10056
rect 16209 9979 16267 9985
rect 16209 9945 16221 9979
rect 16255 9976 16267 9979
rect 18598 9976 18604 9988
rect 16255 9948 18604 9976
rect 16255 9945 16267 9948
rect 16209 9939 16267 9945
rect 18598 9936 18604 9948
rect 18656 9936 18662 9988
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 16301 9095 16359 9101
rect 16301 9061 16313 9095
rect 16347 9092 16359 9095
rect 18138 9092 18144 9104
rect 16347 9064 18144 9092
rect 16347 9061 16359 9064
rect 16301 9055 16359 9061
rect 18138 9052 18144 9064
rect 18196 9052 18202 9104
rect 13354 8916 13360 8968
rect 13412 8956 13418 8968
rect 14737 8959 14795 8965
rect 14737 8956 14749 8959
rect 13412 8928 14749 8956
rect 13412 8916 13418 8928
rect 14737 8925 14749 8928
rect 14783 8956 14795 8959
rect 15381 8959 15439 8965
rect 15381 8956 15393 8959
rect 14783 8928 15393 8956
rect 14783 8925 14795 8928
rect 14737 8919 14795 8925
rect 15381 8925 15393 8928
rect 15427 8925 15439 8959
rect 15381 8919 15439 8925
rect 16022 8916 16028 8968
rect 16080 8956 16086 8968
rect 16117 8959 16175 8965
rect 16117 8956 16129 8959
rect 16080 8928 16129 8956
rect 16080 8916 16086 8928
rect 16117 8925 16129 8928
rect 16163 8956 16175 8959
rect 16761 8959 16819 8965
rect 16761 8956 16773 8959
rect 16163 8928 16773 8956
rect 16163 8925 16175 8928
rect 16117 8919 16175 8925
rect 16761 8925 16773 8928
rect 16807 8925 16819 8959
rect 38010 8956 38016 8968
rect 37971 8928 38016 8956
rect 16761 8919 16819 8925
rect 38010 8916 38016 8928
rect 38068 8916 38074 8968
rect 1670 8888 1676 8900
rect 1631 8860 1676 8888
rect 1670 8848 1676 8860
rect 1728 8848 1734 8900
rect 16850 8888 16856 8900
rect 14936 8860 16856 8888
rect 1765 8823 1823 8829
rect 1765 8789 1777 8823
rect 1811 8820 1823 8823
rect 13630 8820 13636 8832
rect 1811 8792 13636 8820
rect 1811 8789 1823 8792
rect 1765 8783 1823 8789
rect 13630 8780 13636 8792
rect 13688 8780 13694 8832
rect 14936 8829 14964 8860
rect 16850 8848 16856 8860
rect 16908 8848 16914 8900
rect 14921 8823 14979 8829
rect 14921 8789 14933 8823
rect 14967 8789 14979 8823
rect 38194 8820 38200 8832
rect 38155 8792 38200 8820
rect 14921 8783 14979 8789
rect 38194 8780 38200 8792
rect 38252 8780 38258 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 1670 8616 1676 8628
rect 1631 8588 1676 8616
rect 1670 8576 1676 8588
rect 1728 8576 1734 8628
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 37274 7528 37280 7540
rect 26206 7500 37280 7528
rect 22370 7392 22376 7404
rect 22331 7364 22376 7392
rect 22370 7352 22376 7364
rect 22428 7392 22434 7404
rect 23017 7395 23075 7401
rect 23017 7392 23029 7395
rect 22428 7364 23029 7392
rect 22428 7352 22434 7364
rect 23017 7361 23029 7364
rect 23063 7392 23075 7395
rect 26206 7392 26234 7500
rect 37274 7488 37280 7500
rect 37332 7488 37338 7540
rect 37918 7420 37924 7472
rect 37976 7460 37982 7472
rect 38013 7463 38071 7469
rect 38013 7460 38025 7463
rect 37976 7432 38025 7460
rect 37976 7420 37982 7432
rect 38013 7429 38025 7432
rect 38059 7429 38071 7463
rect 38013 7423 38071 7429
rect 23063 7364 26234 7392
rect 37553 7395 37611 7401
rect 23063 7361 23075 7364
rect 23017 7355 23075 7361
rect 37553 7361 37565 7395
rect 37599 7392 37611 7395
rect 38194 7392 38200 7404
rect 37599 7364 38200 7392
rect 37599 7361 37611 7364
rect 37553 7355 37611 7361
rect 38194 7352 38200 7364
rect 38252 7352 38258 7404
rect 1578 7324 1584 7336
rect 1539 7296 1584 7324
rect 1578 7284 1584 7296
rect 1636 7284 1642 7336
rect 1857 7327 1915 7333
rect 1857 7293 1869 7327
rect 1903 7324 1915 7327
rect 10502 7324 10508 7336
rect 1903 7296 10508 7324
rect 1903 7293 1915 7296
rect 1857 7287 1915 7293
rect 10502 7284 10508 7296
rect 10560 7284 10566 7336
rect 22554 7188 22560 7200
rect 22515 7160 22560 7188
rect 22554 7148 22560 7160
rect 22612 7148 22618 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 1578 6984 1584 6996
rect 1539 6956 1584 6984
rect 1578 6944 1584 6956
rect 1636 6944 1642 6996
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 24394 6304 24400 6316
rect 24355 6276 24400 6304
rect 24394 6264 24400 6276
rect 24452 6304 24458 6316
rect 25041 6307 25099 6313
rect 25041 6304 25053 6307
rect 24452 6276 25053 6304
rect 24452 6264 24458 6276
rect 25041 6273 25053 6276
rect 25087 6304 25099 6307
rect 25087 6276 26234 6304
rect 25087 6273 25099 6276
rect 25041 6267 25099 6273
rect 24581 6103 24639 6109
rect 24581 6069 24593 6103
rect 24627 6100 24639 6103
rect 24946 6100 24952 6112
rect 24627 6072 24952 6100
rect 24627 6069 24639 6072
rect 24581 6063 24639 6069
rect 24946 6060 24952 6072
rect 25004 6060 25010 6112
rect 26206 6100 26234 6276
rect 37826 6100 37832 6112
rect 26206 6072 37832 6100
rect 37826 6060 37832 6072
rect 37884 6060 37890 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 38105 5899 38163 5905
rect 38105 5865 38117 5899
rect 38151 5896 38163 5899
rect 38378 5896 38384 5908
rect 38151 5868 38384 5896
rect 38151 5865 38163 5868
rect 38105 5859 38163 5865
rect 38378 5856 38384 5868
rect 38436 5856 38442 5908
rect 37553 5627 37611 5633
rect 37553 5593 37565 5627
rect 37599 5624 37611 5627
rect 38194 5624 38200 5636
rect 37599 5596 38200 5624
rect 37599 5593 37611 5596
rect 37553 5587 37611 5593
rect 38194 5584 38200 5596
rect 38252 5584 38258 5636
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 1762 5352 1768 5364
rect 1723 5324 1768 5352
rect 1762 5312 1768 5324
rect 1820 5312 1826 5364
rect 1578 5176 1584 5228
rect 1636 5216 1642 5228
rect 1673 5219 1731 5225
rect 1673 5216 1685 5219
rect 1636 5188 1685 5216
rect 1636 5176 1642 5188
rect 1673 5185 1685 5188
rect 1719 5185 1731 5219
rect 1673 5179 1731 5185
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 1578 4808 1584 4820
rect 1539 4780 1584 4808
rect 1578 4768 1584 4780
rect 1636 4768 1642 4820
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 1670 3924 1676 3936
rect 1631 3896 1676 3924
rect 1670 3884 1676 3896
rect 1728 3884 1734 3936
rect 38102 3884 38108 3936
rect 38160 3924 38166 3936
rect 38197 3927 38255 3933
rect 38197 3924 38209 3927
rect 38160 3896 38209 3924
rect 38160 3884 38166 3896
rect 38197 3893 38209 3896
rect 38243 3893 38255 3927
rect 38197 3887 38255 3893
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 1857 3655 1915 3661
rect 1857 3621 1869 3655
rect 1903 3652 1915 3655
rect 2866 3652 2872 3664
rect 1903 3624 2872 3652
rect 1903 3621 1915 3624
rect 1857 3615 1915 3621
rect 2866 3612 2872 3624
rect 2924 3612 2930 3664
rect 1670 3516 1676 3528
rect 1631 3488 1676 3516
rect 1670 3476 1676 3488
rect 1728 3476 1734 3528
rect 38013 3519 38071 3525
rect 38013 3516 38025 3519
rect 37476 3488 38025 3516
rect 37366 3340 37372 3392
rect 37424 3380 37430 3392
rect 37476 3389 37504 3488
rect 38013 3485 38025 3488
rect 38059 3485 38071 3519
rect 38013 3479 38071 3485
rect 37461 3383 37519 3389
rect 37461 3380 37473 3383
rect 37424 3352 37473 3380
rect 37424 3340 37430 3352
rect 37461 3349 37473 3352
rect 37507 3349 37519 3383
rect 38194 3380 38200 3392
rect 38155 3352 38200 3380
rect 37461 3343 37519 3349
rect 38194 3340 38200 3352
rect 38252 3340 38258 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 12710 3176 12716 3188
rect 12671 3148 12716 3176
rect 12710 3136 12716 3148
rect 12768 3136 12774 3188
rect 15930 3136 15936 3188
rect 15988 3176 15994 3188
rect 20717 3179 20775 3185
rect 20717 3176 20729 3179
rect 15988 3148 20729 3176
rect 15988 3136 15994 3148
rect 20717 3145 20729 3148
rect 20763 3145 20775 3179
rect 34698 3176 34704 3188
rect 20717 3139 20775 3145
rect 26206 3148 34704 3176
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3040 1915 3043
rect 1946 3040 1952 3052
rect 1903 3012 1952 3040
rect 1903 3009 1915 3012
rect 1857 3003 1915 3009
rect 1946 3000 1952 3012
rect 2004 3000 2010 3052
rect 8662 3040 8668 3052
rect 8623 3012 8668 3040
rect 8662 3000 8668 3012
rect 8720 3000 8726 3052
rect 12253 3043 12311 3049
rect 12253 3009 12265 3043
rect 12299 3040 12311 3043
rect 12728 3040 12756 3136
rect 14918 3068 14924 3120
rect 14976 3108 14982 3120
rect 20622 3108 20628 3120
rect 14976 3080 20628 3108
rect 14976 3068 14982 3080
rect 20622 3068 20628 3080
rect 20680 3068 20686 3120
rect 12299 3012 15700 3040
rect 12299 3009 12311 3012
rect 12253 3003 12311 3009
rect 2406 2972 2412 2984
rect 2319 2944 2412 2972
rect 2406 2932 2412 2944
rect 2464 2972 2470 2984
rect 15562 2972 15568 2984
rect 2464 2944 15568 2972
rect 2464 2932 2470 2944
rect 15562 2932 15568 2944
rect 15620 2932 15626 2984
rect 15672 2972 15700 3012
rect 15746 3000 15752 3052
rect 15804 3040 15810 3052
rect 16114 3040 16120 3052
rect 15804 3012 16120 3040
rect 15804 3000 15810 3012
rect 16114 3000 16120 3012
rect 16172 3040 16178 3052
rect 18693 3043 18751 3049
rect 18693 3040 18705 3043
rect 16172 3012 18705 3040
rect 16172 3000 16178 3012
rect 18693 3009 18705 3012
rect 18739 3040 18751 3043
rect 19337 3043 19395 3049
rect 19337 3040 19349 3043
rect 18739 3012 19349 3040
rect 18739 3009 18751 3012
rect 18693 3003 18751 3009
rect 19337 3009 19349 3012
rect 19383 3009 19395 3043
rect 20732 3040 20760 3139
rect 20806 3068 20812 3120
rect 20864 3108 20870 3120
rect 26206 3108 26234 3148
rect 34698 3136 34704 3148
rect 34756 3136 34762 3188
rect 20864 3080 26234 3108
rect 29733 3111 29791 3117
rect 20864 3068 20870 3080
rect 29733 3077 29745 3111
rect 29779 3108 29791 3111
rect 37274 3108 37280 3120
rect 29779 3080 37280 3108
rect 29779 3077 29791 3080
rect 29733 3071 29791 3077
rect 21269 3043 21327 3049
rect 21269 3040 21281 3043
rect 20732 3012 21281 3040
rect 19337 3003 19395 3009
rect 21269 3009 21281 3012
rect 21315 3009 21327 3043
rect 28994 3040 29000 3052
rect 28907 3012 29000 3040
rect 21269 3003 21327 3009
rect 28994 3000 29000 3012
rect 29052 3040 29058 3052
rect 29748 3040 29776 3071
rect 37274 3068 37280 3080
rect 37332 3068 37338 3120
rect 37734 3068 37740 3120
rect 37792 3108 37798 3120
rect 38013 3111 38071 3117
rect 38013 3108 38025 3111
rect 37792 3080 38025 3108
rect 37792 3068 37798 3080
rect 38013 3077 38025 3080
rect 38059 3077 38071 3111
rect 38013 3071 38071 3077
rect 29052 3012 29776 3040
rect 36909 3043 36967 3049
rect 29052 3000 29058 3012
rect 36909 3009 36921 3043
rect 36955 3040 36967 3043
rect 38194 3040 38200 3052
rect 36955 3012 38200 3040
rect 36955 3009 36967 3012
rect 36909 3003 36967 3009
rect 38194 3000 38200 3012
rect 38252 3000 38258 3052
rect 30282 2972 30288 2984
rect 15672 2944 30288 2972
rect 30282 2932 30288 2944
rect 30340 2932 30346 2984
rect 36722 2932 36728 2984
rect 36780 2972 36786 2984
rect 37461 2975 37519 2981
rect 37461 2972 37473 2975
rect 36780 2944 37473 2972
rect 36780 2932 36786 2944
rect 37461 2941 37473 2944
rect 37507 2941 37519 2975
rect 37461 2935 37519 2941
rect 4706 2864 4712 2916
rect 4764 2904 4770 2916
rect 12069 2907 12127 2913
rect 12069 2904 12081 2907
rect 4764 2876 12081 2904
rect 4764 2864 4770 2876
rect 12069 2873 12081 2876
rect 12115 2873 12127 2907
rect 12069 2867 12127 2873
rect 18877 2907 18935 2913
rect 18877 2873 18889 2907
rect 18923 2904 18935 2907
rect 37366 2904 37372 2916
rect 18923 2876 37372 2904
rect 18923 2873 18935 2876
rect 18877 2867 18935 2873
rect 37366 2864 37372 2876
rect 37424 2864 37430 2916
rect 1670 2836 1676 2848
rect 1631 2808 1676 2836
rect 1670 2796 1676 2808
rect 1728 2796 1734 2848
rect 4525 2839 4583 2845
rect 4525 2805 4537 2839
rect 4571 2836 4583 2839
rect 4614 2836 4620 2848
rect 4571 2808 4620 2836
rect 4571 2805 4583 2808
rect 4525 2799 4583 2805
rect 4614 2796 4620 2808
rect 4672 2796 4678 2848
rect 8481 2839 8539 2845
rect 8481 2805 8493 2839
rect 8527 2836 8539 2839
rect 8570 2836 8576 2848
rect 8527 2808 8576 2836
rect 8527 2805 8539 2808
rect 8481 2799 8539 2805
rect 8570 2796 8576 2808
rect 8628 2796 8634 2848
rect 21361 2839 21419 2845
rect 21361 2805 21373 2839
rect 21407 2836 21419 2839
rect 23382 2836 23388 2848
rect 21407 2808 23388 2836
rect 21407 2805 21419 2808
rect 21361 2799 21419 2805
rect 23382 2796 23388 2808
rect 23440 2796 23446 2848
rect 29178 2836 29184 2848
rect 29139 2808 29184 2836
rect 29178 2796 29184 2808
rect 29236 2796 29242 2848
rect 36354 2836 36360 2848
rect 36315 2808 36360 2836
rect 36354 2796 36360 2808
rect 36412 2796 36418 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 4157 2635 4215 2641
rect 4157 2601 4169 2635
rect 4203 2632 4215 2635
rect 8662 2632 8668 2644
rect 4203 2604 8668 2632
rect 4203 2601 4215 2604
rect 4157 2595 4215 2601
rect 8662 2592 8668 2604
rect 8720 2592 8726 2644
rect 15746 2632 15752 2644
rect 10060 2604 15752 2632
rect 14 2524 20 2576
rect 72 2564 78 2576
rect 2409 2567 2467 2573
rect 2409 2564 2421 2567
rect 72 2536 2421 2564
rect 72 2524 78 2536
rect 2409 2533 2421 2536
rect 2455 2533 2467 2567
rect 2409 2527 2467 2533
rect 2958 2524 2964 2576
rect 3016 2564 3022 2576
rect 4617 2567 4675 2573
rect 4617 2564 4629 2567
rect 3016 2536 4629 2564
rect 3016 2524 3022 2536
rect 4617 2533 4629 2536
rect 4663 2533 4675 2567
rect 4617 2527 4675 2533
rect 4706 2496 4712 2508
rect 2608 2468 4712 2496
rect 1857 2431 1915 2437
rect 1857 2397 1869 2431
rect 1903 2428 1915 2431
rect 2406 2428 2412 2440
rect 1903 2400 2412 2428
rect 1903 2397 1915 2400
rect 1857 2391 1915 2397
rect 2406 2388 2412 2400
rect 2464 2388 2470 2440
rect 2608 2437 2636 2468
rect 4706 2456 4712 2468
rect 4764 2456 4770 2508
rect 10060 2505 10088 2604
rect 15746 2592 15752 2604
rect 15804 2592 15810 2644
rect 28534 2632 28540 2644
rect 28495 2604 28540 2632
rect 28534 2592 28540 2604
rect 28592 2592 28598 2644
rect 33686 2632 33692 2644
rect 33647 2604 33692 2632
rect 33686 2592 33692 2604
rect 33744 2592 33750 2644
rect 35989 2635 36047 2641
rect 35989 2632 36001 2635
rect 33796 2604 36001 2632
rect 11974 2564 11980 2576
rect 11935 2536 11980 2564
rect 11974 2524 11980 2536
rect 12032 2524 12038 2576
rect 15197 2567 15255 2573
rect 15197 2533 15209 2567
rect 15243 2564 15255 2567
rect 15654 2564 15660 2576
rect 15243 2536 15660 2564
rect 15243 2533 15255 2536
rect 15197 2527 15255 2533
rect 15654 2524 15660 2536
rect 15712 2524 15718 2576
rect 30282 2524 30288 2576
rect 30340 2564 30346 2576
rect 32309 2567 32367 2573
rect 32309 2564 32321 2567
rect 30340 2536 32321 2564
rect 30340 2524 30346 2536
rect 32309 2533 32321 2536
rect 32355 2533 32367 2567
rect 32309 2527 32367 2533
rect 10045 2499 10103 2505
rect 10045 2465 10057 2499
rect 10091 2465 10103 2499
rect 10045 2459 10103 2465
rect 15378 2456 15384 2508
rect 15436 2496 15442 2508
rect 33796 2496 33824 2604
rect 35989 2601 36001 2604
rect 36035 2601 36047 2635
rect 35989 2595 36047 2601
rect 34790 2524 34796 2576
rect 34848 2564 34854 2576
rect 36633 2567 36691 2573
rect 36633 2564 36645 2567
rect 34848 2536 36645 2564
rect 34848 2524 34854 2536
rect 36633 2533 36645 2536
rect 36679 2533 36691 2567
rect 36633 2527 36691 2533
rect 15436 2468 33824 2496
rect 15436 2456 15442 2468
rect 37274 2456 37280 2508
rect 37332 2496 37338 2508
rect 38013 2499 38071 2505
rect 38013 2496 38025 2499
rect 37332 2468 38025 2496
rect 37332 2456 37338 2468
rect 38013 2465 38025 2468
rect 38059 2465 38071 2499
rect 38013 2459 38071 2465
rect 2593 2431 2651 2437
rect 2593 2397 2605 2431
rect 2639 2397 2651 2431
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 2593 2391 2651 2397
rect 3344 2400 3985 2428
rect 1302 2252 1308 2304
rect 1360 2292 1366 2304
rect 1673 2295 1731 2301
rect 1673 2292 1685 2295
rect 1360 2264 1685 2292
rect 1360 2252 1366 2264
rect 1673 2261 1685 2264
rect 1719 2261 1731 2295
rect 1673 2255 1731 2261
rect 3234 2252 3240 2304
rect 3292 2292 3298 2304
rect 3344 2301 3372 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 6822 2428 6828 2440
rect 6783 2400 6828 2428
rect 3973 2391 4031 2397
rect 6822 2388 6828 2400
rect 6880 2388 6886 2440
rect 8570 2428 8576 2440
rect 8531 2400 8576 2428
rect 8570 2388 8576 2400
rect 8628 2388 8634 2440
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2428 9367 2431
rect 9674 2428 9680 2440
rect 9355 2400 9680 2428
rect 9355 2397 9367 2400
rect 9309 2391 9367 2397
rect 9674 2388 9680 2400
rect 9732 2428 9738 2440
rect 9769 2431 9827 2437
rect 9769 2428 9781 2431
rect 9732 2400 9781 2428
rect 9732 2388 9738 2400
rect 9769 2397 9781 2400
rect 9815 2397 9827 2431
rect 9769 2391 9827 2397
rect 10870 2388 10876 2440
rect 10928 2428 10934 2440
rect 12989 2431 13047 2437
rect 12989 2428 13001 2431
rect 10928 2400 13001 2428
rect 10928 2388 10934 2400
rect 12989 2397 13001 2400
rect 13035 2397 13047 2431
rect 16850 2428 16856 2440
rect 16811 2400 16856 2428
rect 12989 2391 13047 2397
rect 16850 2388 16856 2400
rect 16908 2388 16914 2440
rect 18138 2428 18144 2440
rect 18099 2400 18144 2428
rect 18138 2388 18144 2400
rect 18196 2388 18202 2440
rect 18598 2388 18604 2440
rect 18656 2428 18662 2440
rect 20073 2431 20131 2437
rect 20073 2428 20085 2431
rect 18656 2400 20085 2428
rect 18656 2388 18662 2400
rect 20073 2397 20085 2400
rect 20119 2397 20131 2431
rect 22002 2428 22008 2440
rect 21963 2400 22008 2428
rect 20073 2391 20131 2397
rect 22002 2388 22008 2400
rect 22060 2388 22066 2440
rect 22554 2388 22560 2440
rect 22612 2428 22618 2440
rect 23293 2431 23351 2437
rect 23293 2428 23305 2431
rect 22612 2400 23305 2428
rect 22612 2388 22618 2400
rect 23293 2397 23305 2400
rect 23339 2397 23351 2431
rect 23293 2391 23351 2397
rect 24946 2388 24952 2440
rect 25004 2428 25010 2440
rect 25225 2431 25283 2437
rect 25225 2428 25237 2431
rect 25004 2400 25237 2428
rect 25004 2388 25010 2400
rect 25225 2397 25237 2400
rect 25271 2397 25283 2431
rect 27157 2431 27215 2437
rect 27157 2428 27169 2431
rect 25225 2391 25283 2397
rect 26206 2400 27169 2428
rect 4522 2320 4528 2372
rect 4580 2360 4586 2372
rect 4801 2363 4859 2369
rect 4801 2360 4813 2363
rect 4580 2332 4813 2360
rect 4580 2320 4586 2332
rect 4801 2329 4813 2332
rect 4847 2329 4859 2363
rect 4801 2323 4859 2329
rect 11149 2363 11207 2369
rect 11149 2329 11161 2363
rect 11195 2360 11207 2363
rect 11606 2360 11612 2372
rect 11195 2332 11612 2360
rect 11195 2329 11207 2332
rect 11149 2323 11207 2329
rect 11606 2320 11612 2332
rect 11664 2360 11670 2372
rect 11793 2363 11851 2369
rect 11793 2360 11805 2363
rect 11664 2332 11805 2360
rect 11664 2320 11670 2332
rect 11793 2329 11805 2332
rect 11839 2329 11851 2363
rect 11793 2323 11851 2329
rect 14461 2363 14519 2369
rect 14461 2329 14473 2363
rect 14507 2360 14519 2363
rect 14826 2360 14832 2372
rect 14507 2332 14832 2360
rect 14507 2329 14519 2332
rect 14461 2323 14519 2329
rect 14826 2320 14832 2332
rect 14884 2360 14890 2372
rect 15013 2363 15071 2369
rect 15013 2360 15025 2363
rect 14884 2332 15025 2360
rect 14884 2320 14890 2332
rect 15013 2329 15025 2332
rect 15059 2329 15071 2363
rect 15013 2323 15071 2329
rect 23382 2320 23388 2372
rect 23440 2360 23446 2372
rect 26206 2360 26234 2400
rect 27157 2397 27169 2400
rect 27203 2397 27215 2431
rect 27157 2391 27215 2397
rect 29178 2388 29184 2440
rect 29236 2428 29242 2440
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29236 2400 29745 2428
rect 29236 2388 29242 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 34698 2388 34704 2440
rect 34756 2428 34762 2440
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 34756 2400 34897 2428
rect 34756 2388 34762 2400
rect 34885 2397 34897 2400
rect 34931 2397 34943 2431
rect 34885 2391 34943 2397
rect 36173 2431 36231 2437
rect 36173 2397 36185 2431
rect 36219 2428 36231 2431
rect 36354 2428 36360 2440
rect 36219 2400 36360 2428
rect 36219 2397 36231 2400
rect 36173 2391 36231 2397
rect 36354 2388 36360 2400
rect 36412 2428 36418 2440
rect 37182 2428 37188 2440
rect 36412 2400 37188 2428
rect 36412 2388 36418 2400
rect 37182 2388 37188 2400
rect 37240 2388 37246 2440
rect 38102 2388 38108 2440
rect 38160 2428 38166 2440
rect 38289 2431 38347 2437
rect 38289 2428 38301 2431
rect 38160 2400 38301 2428
rect 38160 2388 38166 2400
rect 38289 2397 38301 2400
rect 38335 2397 38347 2431
rect 38289 2391 38347 2397
rect 23440 2332 26234 2360
rect 27985 2363 28043 2369
rect 23440 2320 23446 2332
rect 27985 2329 27997 2363
rect 28031 2360 28043 2363
rect 28350 2360 28356 2372
rect 28031 2332 28356 2360
rect 28031 2329 28043 2332
rect 27985 2323 28043 2329
rect 28350 2320 28356 2332
rect 28408 2360 28414 2372
rect 28629 2363 28687 2369
rect 28629 2360 28641 2363
rect 28408 2332 28641 2360
rect 28408 2320 28414 2332
rect 28629 2329 28641 2332
rect 28675 2329 28687 2363
rect 32493 2363 32551 2369
rect 32493 2360 32505 2363
rect 28629 2323 28687 2329
rect 31772 2332 32505 2360
rect 31772 2304 31800 2332
rect 32493 2329 32505 2332
rect 32539 2329 32551 2363
rect 32493 2323 32551 2329
rect 33137 2363 33195 2369
rect 33137 2329 33149 2363
rect 33183 2360 33195 2363
rect 33502 2360 33508 2372
rect 33183 2332 33508 2360
rect 33183 2329 33195 2332
rect 33137 2323 33195 2329
rect 33502 2320 33508 2332
rect 33560 2360 33566 2372
rect 33781 2363 33839 2369
rect 33781 2360 33793 2363
rect 33560 2332 33793 2360
rect 33560 2320 33566 2332
rect 33781 2329 33793 2332
rect 33827 2329 33839 2363
rect 33781 2323 33839 2329
rect 36722 2320 36728 2372
rect 36780 2360 36786 2372
rect 36817 2363 36875 2369
rect 36817 2360 36829 2363
rect 36780 2332 36829 2360
rect 36780 2320 36786 2332
rect 36817 2329 36829 2332
rect 36863 2329 36875 2363
rect 36817 2323 36875 2329
rect 3329 2295 3387 2301
rect 3329 2292 3341 2295
rect 3292 2264 3341 2292
rect 3292 2252 3298 2264
rect 3329 2261 3341 2264
rect 3375 2261 3387 2295
rect 3329 2255 3387 2261
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 6641 2295 6699 2301
rect 6641 2292 6653 2295
rect 6512 2264 6653 2292
rect 6512 2252 6518 2264
rect 6641 2261 6653 2264
rect 6687 2261 6699 2295
rect 8386 2292 8392 2304
rect 8347 2264 8392 2292
rect 6641 2255 6699 2261
rect 8386 2252 8392 2264
rect 8444 2252 8450 2304
rect 12894 2252 12900 2304
rect 12952 2292 12958 2304
rect 13173 2295 13231 2301
rect 13173 2292 13185 2295
rect 12952 2264 13185 2292
rect 12952 2252 12958 2264
rect 13173 2261 13185 2264
rect 13219 2261 13231 2295
rect 13173 2255 13231 2261
rect 16758 2252 16764 2304
rect 16816 2292 16822 2304
rect 17037 2295 17095 2301
rect 17037 2292 17049 2295
rect 16816 2264 17049 2292
rect 16816 2252 16822 2264
rect 17037 2261 17049 2264
rect 17083 2261 17095 2295
rect 17037 2255 17095 2261
rect 18046 2252 18052 2304
rect 18104 2292 18110 2304
rect 18325 2295 18383 2301
rect 18325 2292 18337 2295
rect 18104 2264 18337 2292
rect 18104 2252 18110 2264
rect 18325 2261 18337 2264
rect 18371 2261 18383 2295
rect 18325 2255 18383 2261
rect 19978 2252 19984 2304
rect 20036 2292 20042 2304
rect 20257 2295 20315 2301
rect 20257 2292 20269 2295
rect 20036 2264 20269 2292
rect 20036 2252 20042 2264
rect 20257 2261 20269 2264
rect 20303 2261 20315 2295
rect 20257 2255 20315 2261
rect 21266 2252 21272 2304
rect 21324 2292 21330 2304
rect 22189 2295 22247 2301
rect 22189 2292 22201 2295
rect 21324 2264 22201 2292
rect 21324 2252 21330 2264
rect 22189 2261 22201 2264
rect 22235 2261 22247 2295
rect 22189 2255 22247 2261
rect 23198 2252 23204 2304
rect 23256 2292 23262 2304
rect 23477 2295 23535 2301
rect 23477 2292 23489 2295
rect 23256 2264 23489 2292
rect 23256 2252 23262 2264
rect 23477 2261 23489 2264
rect 23523 2261 23535 2295
rect 23477 2255 23535 2261
rect 25130 2252 25136 2304
rect 25188 2292 25194 2304
rect 25409 2295 25467 2301
rect 25409 2292 25421 2295
rect 25188 2264 25421 2292
rect 25188 2252 25194 2264
rect 25409 2261 25421 2264
rect 25455 2261 25467 2295
rect 25409 2255 25467 2261
rect 26418 2252 26424 2304
rect 26476 2292 26482 2304
rect 27341 2295 27399 2301
rect 27341 2292 27353 2295
rect 26476 2264 27353 2292
rect 26476 2252 26482 2264
rect 27341 2261 27353 2264
rect 27387 2261 27399 2295
rect 27341 2255 27399 2261
rect 29638 2252 29644 2304
rect 29696 2292 29702 2304
rect 29917 2295 29975 2301
rect 29917 2292 29929 2295
rect 29696 2264 29929 2292
rect 29696 2252 29702 2264
rect 29917 2261 29929 2264
rect 29963 2261 29975 2295
rect 31754 2292 31760 2304
rect 31715 2264 31760 2292
rect 29917 2255 29975 2261
rect 31754 2252 31760 2264
rect 31812 2252 31818 2304
rect 34790 2252 34796 2304
rect 34848 2292 34854 2304
rect 35069 2295 35127 2301
rect 35069 2292 35081 2295
rect 34848 2264 35081 2292
rect 34848 2252 34854 2264
rect 35069 2261 35081 2264
rect 35115 2261 35127 2295
rect 35069 2255 35127 2261
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 14280 37680 14332 37732
rect 21548 37680 21600 37732
rect 13176 37612 13228 37664
rect 16120 37612 16172 37664
rect 16488 37612 16540 37664
rect 18880 37612 18932 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 8208 37408 8260 37460
rect 22836 37408 22888 37460
rect 38200 37408 38252 37460
rect 38660 37408 38712 37460
rect 16028 37383 16080 37392
rect 20 37272 72 37324
rect 2320 37272 2372 37324
rect 6552 37272 6604 37324
rect 16028 37349 16037 37383
rect 16037 37349 16071 37383
rect 16071 37349 16080 37383
rect 16028 37340 16080 37349
rect 16396 37340 16448 37392
rect 1676 37247 1728 37256
rect 1676 37213 1685 37247
rect 1685 37213 1719 37247
rect 1719 37213 1728 37247
rect 1676 37204 1728 37213
rect 4620 37204 4672 37256
rect 1860 37136 1912 37188
rect 2688 37136 2740 37188
rect 3884 37136 3936 37188
rect 8208 37204 8260 37256
rect 3332 37068 3384 37120
rect 4252 37111 4304 37120
rect 4252 37077 4261 37111
rect 4261 37077 4295 37111
rect 4295 37077 4304 37111
rect 4252 37068 4304 37077
rect 11244 37272 11296 37324
rect 13176 37315 13228 37324
rect 13176 37281 13185 37315
rect 13185 37281 13219 37315
rect 13219 37281 13228 37315
rect 13176 37272 13228 37281
rect 14556 37272 14608 37324
rect 9128 37204 9180 37256
rect 14004 37204 14056 37256
rect 16488 37204 16540 37256
rect 16672 37272 16724 37324
rect 21548 37340 21600 37392
rect 16856 37204 16908 37256
rect 17132 37247 17184 37256
rect 17132 37213 17141 37247
rect 17141 37213 17175 37247
rect 17175 37213 17184 37247
rect 17132 37204 17184 37213
rect 19248 37272 19300 37324
rect 23940 37315 23992 37324
rect 9588 37136 9640 37188
rect 10692 37136 10744 37188
rect 12716 37136 12768 37188
rect 12900 37136 12952 37188
rect 14188 37136 14240 37188
rect 14648 37136 14700 37188
rect 19432 37247 19484 37256
rect 19432 37213 19441 37247
rect 19441 37213 19475 37247
rect 19475 37213 19484 37247
rect 19432 37204 19484 37213
rect 19984 37204 20036 37256
rect 20720 37204 20772 37256
rect 23940 37281 23949 37315
rect 23949 37281 23983 37315
rect 23983 37281 23992 37315
rect 23940 37272 23992 37281
rect 22744 37247 22796 37256
rect 22744 37213 22753 37247
rect 22753 37213 22787 37247
rect 22787 37213 22796 37247
rect 22744 37204 22796 37213
rect 6000 37068 6052 37120
rect 10968 37068 11020 37120
rect 11152 37111 11204 37120
rect 11152 37077 11161 37111
rect 11161 37077 11195 37111
rect 11195 37077 11204 37111
rect 11152 37068 11204 37077
rect 11704 37111 11756 37120
rect 11704 37077 11713 37111
rect 11713 37077 11747 37111
rect 11747 37077 11756 37111
rect 11704 37068 11756 37077
rect 12532 37068 12584 37120
rect 16028 37068 16080 37120
rect 16580 37068 16632 37120
rect 16764 37068 16816 37120
rect 17684 37111 17736 37120
rect 17684 37077 17693 37111
rect 17693 37077 17727 37111
rect 17727 37077 17736 37111
rect 17684 37068 17736 37077
rect 18696 37068 18748 37120
rect 20444 37136 20496 37188
rect 29184 37272 29236 37324
rect 35440 37272 35492 37324
rect 25320 37247 25372 37256
rect 21916 37068 21968 37120
rect 22652 37068 22704 37120
rect 22928 37068 22980 37120
rect 25320 37213 25329 37247
rect 25329 37213 25363 37247
rect 25363 37213 25372 37247
rect 25320 37204 25372 37213
rect 26516 37204 26568 37256
rect 29736 37247 29788 37256
rect 29736 37213 29745 37247
rect 29745 37213 29779 37247
rect 29779 37213 29788 37247
rect 29736 37204 29788 37213
rect 30380 37204 30432 37256
rect 32312 37247 32364 37256
rect 32312 37213 32321 37247
rect 32321 37213 32355 37247
rect 32355 37213 32364 37247
rect 32312 37204 32364 37213
rect 33968 37204 34020 37256
rect 24768 37111 24820 37120
rect 24768 37077 24777 37111
rect 24777 37077 24811 37111
rect 24811 37077 24820 37111
rect 24768 37068 24820 37077
rect 25136 37068 25188 37120
rect 26516 37111 26568 37120
rect 26516 37077 26525 37111
rect 26525 37077 26559 37111
rect 26559 37077 26568 37111
rect 26516 37068 26568 37077
rect 27068 37068 27120 37120
rect 28448 37111 28500 37120
rect 28448 37077 28457 37111
rect 28457 37077 28491 37111
rect 28491 37077 28500 37111
rect 28448 37068 28500 37077
rect 29000 37068 29052 37120
rect 30564 37136 30616 37188
rect 32220 37068 32272 37120
rect 33508 37068 33560 37120
rect 36820 37111 36872 37120
rect 36820 37077 36829 37111
rect 36829 37077 36863 37111
rect 36863 37077 36872 37111
rect 36820 37068 36872 37077
rect 37372 37068 37424 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 1676 36864 1728 36916
rect 3884 36864 3936 36916
rect 940 36796 992 36848
rect 5908 36864 5960 36916
rect 11888 36864 11940 36916
rect 6276 36796 6328 36848
rect 9680 36796 9732 36848
rect 10968 36796 11020 36848
rect 11152 36796 11204 36848
rect 14556 36864 14608 36916
rect 15752 36864 15804 36916
rect 17224 36864 17276 36916
rect 22744 36864 22796 36916
rect 23848 36864 23900 36916
rect 24768 36864 24820 36916
rect 29736 36864 29788 36916
rect 3884 36728 3936 36780
rect 4068 36660 4120 36712
rect 6368 36660 6420 36712
rect 6828 36703 6880 36712
rect 6828 36669 6837 36703
rect 6837 36669 6871 36703
rect 6871 36669 6880 36703
rect 6828 36660 6880 36669
rect 7196 36660 7248 36712
rect 8116 36660 8168 36712
rect 9036 36660 9088 36712
rect 9128 36660 9180 36712
rect 11612 36728 11664 36780
rect 17040 36728 17092 36780
rect 17500 36728 17552 36780
rect 17868 36728 17920 36780
rect 18972 36728 19024 36780
rect 20444 36771 20496 36780
rect 20444 36737 20453 36771
rect 20453 36737 20487 36771
rect 20487 36737 20496 36771
rect 20444 36728 20496 36737
rect 20720 36796 20772 36848
rect 22560 36796 22612 36848
rect 11060 36660 11112 36712
rect 14004 36703 14056 36712
rect 14004 36669 14013 36703
rect 14013 36669 14047 36703
rect 14047 36669 14056 36703
rect 14004 36660 14056 36669
rect 4252 36524 4304 36576
rect 4988 36524 5040 36576
rect 6276 36524 6328 36576
rect 11612 36592 11664 36644
rect 13084 36592 13136 36644
rect 17224 36660 17276 36712
rect 20168 36703 20220 36712
rect 20168 36669 20177 36703
rect 20177 36669 20211 36703
rect 20211 36669 20220 36703
rect 20168 36660 20220 36669
rect 20628 36660 20680 36712
rect 23020 36728 23072 36780
rect 27068 36796 27120 36848
rect 36820 36796 36872 36848
rect 38200 36839 38252 36848
rect 38200 36805 38209 36839
rect 38209 36805 38243 36839
rect 38243 36805 38252 36839
rect 38200 36796 38252 36805
rect 32312 36728 32364 36780
rect 22744 36660 22796 36712
rect 24032 36703 24084 36712
rect 24032 36669 24041 36703
rect 24041 36669 24075 36703
rect 24075 36669 24084 36703
rect 24032 36660 24084 36669
rect 25688 36660 25740 36712
rect 25780 36660 25832 36712
rect 29644 36703 29696 36712
rect 29644 36669 29653 36703
rect 29653 36669 29687 36703
rect 29687 36669 29696 36703
rect 29644 36660 29696 36669
rect 27068 36592 27120 36644
rect 38016 36635 38068 36644
rect 38016 36601 38025 36635
rect 38025 36601 38059 36635
rect 38059 36601 38068 36635
rect 38016 36592 38068 36601
rect 11796 36524 11848 36576
rect 12992 36524 13044 36576
rect 14280 36567 14332 36576
rect 14280 36533 14310 36567
rect 14310 36533 14332 36567
rect 14280 36524 14332 36533
rect 16120 36524 16172 36576
rect 16304 36567 16356 36576
rect 16304 36533 16313 36567
rect 16313 36533 16347 36567
rect 16347 36533 16356 36567
rect 16304 36524 16356 36533
rect 16672 36524 16724 36576
rect 18604 36567 18656 36576
rect 18604 36533 18613 36567
rect 18613 36533 18647 36567
rect 18647 36533 18656 36567
rect 18604 36524 18656 36533
rect 19156 36524 19208 36576
rect 22560 36524 22612 36576
rect 22836 36524 22888 36576
rect 24676 36567 24728 36576
rect 24676 36533 24685 36567
rect 24685 36533 24719 36567
rect 24719 36533 24728 36567
rect 24676 36524 24728 36533
rect 28448 36524 28500 36576
rect 37464 36524 37516 36576
rect 37924 36524 37976 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 4620 36320 4672 36372
rect 7196 36320 7248 36372
rect 3700 36184 3752 36236
rect 3884 36184 3936 36236
rect 6828 36227 6880 36236
rect 6828 36193 6837 36227
rect 6837 36193 6871 36227
rect 6871 36193 6880 36227
rect 6828 36184 6880 36193
rect 7748 36184 7800 36236
rect 1676 36159 1728 36168
rect 1676 36125 1685 36159
rect 1685 36125 1719 36159
rect 1719 36125 1728 36159
rect 1676 36116 1728 36125
rect 3976 36159 4028 36168
rect 3976 36125 3985 36159
rect 3985 36125 4019 36159
rect 4019 36125 4028 36159
rect 3976 36116 4028 36125
rect 8208 36116 8260 36168
rect 2964 36048 3016 36100
rect 4988 36048 5040 36100
rect 4068 35980 4120 36032
rect 6920 35980 6972 36032
rect 7196 36048 7248 36100
rect 10968 36184 11020 36236
rect 11612 36320 11664 36372
rect 13728 36320 13780 36372
rect 12716 36252 12768 36304
rect 11612 36227 11664 36236
rect 11612 36193 11621 36227
rect 11621 36193 11655 36227
rect 11655 36193 11664 36227
rect 11612 36184 11664 36193
rect 12624 36184 12676 36236
rect 13084 36227 13136 36236
rect 13084 36193 13093 36227
rect 13093 36193 13127 36227
rect 13127 36193 13136 36227
rect 13084 36184 13136 36193
rect 14280 36184 14332 36236
rect 19432 36320 19484 36372
rect 17040 36252 17092 36304
rect 19064 36184 19116 36236
rect 20720 36252 20772 36304
rect 23020 36320 23072 36372
rect 23848 36363 23900 36372
rect 23848 36329 23857 36363
rect 23857 36329 23891 36363
rect 23891 36329 23900 36363
rect 23848 36320 23900 36329
rect 37188 36320 37240 36372
rect 38292 36320 38344 36372
rect 21640 36252 21692 36304
rect 8576 36116 8628 36168
rect 9128 36159 9180 36168
rect 9128 36125 9137 36159
rect 9137 36125 9171 36159
rect 9171 36125 9180 36159
rect 9128 36116 9180 36125
rect 11060 36116 11112 36168
rect 9496 36048 9548 36100
rect 11888 36048 11940 36100
rect 13452 36048 13504 36100
rect 10692 35980 10744 36032
rect 10876 36023 10928 36032
rect 10876 35989 10885 36023
rect 10885 35989 10919 36023
rect 10919 35989 10928 36023
rect 10876 35980 10928 35989
rect 10968 35980 11020 36032
rect 13176 35980 13228 36032
rect 13268 35980 13320 36032
rect 13912 35980 13964 36032
rect 16764 36116 16816 36168
rect 17224 36159 17276 36168
rect 17224 36125 17233 36159
rect 17233 36125 17267 36159
rect 17267 36125 17276 36159
rect 17224 36116 17276 36125
rect 17868 36159 17920 36168
rect 17868 36125 17877 36159
rect 17877 36125 17911 36159
rect 17911 36125 17920 36159
rect 17868 36116 17920 36125
rect 18972 36116 19024 36168
rect 15108 36048 15160 36100
rect 15752 36091 15804 36100
rect 15752 36057 15761 36091
rect 15761 36057 15795 36091
rect 15795 36057 15804 36091
rect 15752 36048 15804 36057
rect 18788 36048 18840 36100
rect 22744 36227 22796 36236
rect 22744 36193 22753 36227
rect 22753 36193 22787 36227
rect 22787 36193 22796 36227
rect 22744 36184 22796 36193
rect 20444 36116 20496 36168
rect 20628 36116 20680 36168
rect 37832 36116 37884 36168
rect 37924 36116 37976 36168
rect 20720 36048 20772 36100
rect 22652 36091 22704 36100
rect 16580 35980 16632 36032
rect 17408 35980 17460 36032
rect 17960 36023 18012 36032
rect 17960 35989 17969 36023
rect 17969 35989 18003 36023
rect 18003 35989 18012 36023
rect 17960 35980 18012 35989
rect 18052 35980 18104 36032
rect 22652 36057 22661 36091
rect 22661 36057 22695 36091
rect 22695 36057 22704 36091
rect 22652 36048 22704 36057
rect 24676 36023 24728 36032
rect 24676 35989 24685 36023
rect 24685 35989 24719 36023
rect 24719 35989 24728 36023
rect 24676 35980 24728 35989
rect 27344 36023 27396 36032
rect 27344 35989 27353 36023
rect 27353 35989 27387 36023
rect 27387 35989 27396 36023
rect 27344 35980 27396 35989
rect 27896 36023 27948 36032
rect 27896 35989 27905 36023
rect 27905 35989 27939 36023
rect 27939 35989 27948 36023
rect 27896 35980 27948 35989
rect 28448 36023 28500 36032
rect 28448 35989 28457 36023
rect 28457 35989 28491 36023
rect 28491 35989 28500 36023
rect 28448 35980 28500 35989
rect 29000 36023 29052 36032
rect 29000 35989 29009 36023
rect 29009 35989 29043 36023
rect 29043 35989 29052 36023
rect 29000 35980 29052 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 3884 35776 3936 35828
rect 1308 35708 1360 35760
rect 5264 35708 5316 35760
rect 5724 35751 5776 35760
rect 5724 35717 5733 35751
rect 5733 35717 5767 35751
rect 5767 35717 5776 35751
rect 5724 35708 5776 35717
rect 1676 35640 1728 35692
rect 8392 35776 8444 35828
rect 9128 35776 9180 35828
rect 9220 35776 9272 35828
rect 9772 35776 9824 35828
rect 10324 35776 10376 35828
rect 11612 35776 11664 35828
rect 8852 35708 8904 35760
rect 7104 35683 7156 35692
rect 7104 35649 7113 35683
rect 7113 35649 7147 35683
rect 7147 35649 7156 35683
rect 7104 35640 7156 35649
rect 10876 35708 10928 35760
rect 14924 35708 14976 35760
rect 15108 35708 15160 35760
rect 15476 35708 15528 35760
rect 10784 35640 10836 35692
rect 14096 35640 14148 35692
rect 16396 35640 16448 35692
rect 16672 35640 16724 35692
rect 16948 35640 17000 35692
rect 19984 35776 20036 35828
rect 19432 35708 19484 35760
rect 19800 35708 19852 35760
rect 20076 35708 20128 35760
rect 27160 35751 27212 35760
rect 2412 35572 2464 35624
rect 4988 35572 5040 35624
rect 4712 35504 4764 35556
rect 9220 35572 9272 35624
rect 8300 35504 8352 35556
rect 11060 35572 11112 35624
rect 12624 35572 12676 35624
rect 13820 35572 13872 35624
rect 13084 35504 13136 35556
rect 14372 35504 14424 35556
rect 3700 35436 3752 35488
rect 6460 35436 6512 35488
rect 7196 35436 7248 35488
rect 10600 35436 10652 35488
rect 13636 35436 13688 35488
rect 14280 35436 14332 35488
rect 16580 35572 16632 35624
rect 19984 35640 20036 35692
rect 20168 35640 20220 35692
rect 20812 35640 20864 35692
rect 27160 35717 27169 35751
rect 27169 35717 27203 35751
rect 27203 35717 27212 35751
rect 27160 35708 27212 35717
rect 22744 35640 22796 35692
rect 22836 35640 22888 35692
rect 30564 35640 30616 35692
rect 18880 35572 18932 35624
rect 23204 35615 23256 35624
rect 23204 35581 23213 35615
rect 23213 35581 23247 35615
rect 23247 35581 23256 35615
rect 23204 35572 23256 35581
rect 16764 35504 16816 35556
rect 22376 35504 22428 35556
rect 17040 35436 17092 35488
rect 18236 35436 18288 35488
rect 20260 35479 20312 35488
rect 20260 35445 20269 35479
rect 20269 35445 20303 35479
rect 20303 35445 20312 35479
rect 20260 35436 20312 35445
rect 22100 35479 22152 35488
rect 22100 35445 22109 35479
rect 22109 35445 22143 35479
rect 22143 35445 22152 35479
rect 22744 35479 22796 35488
rect 22100 35436 22152 35445
rect 22744 35445 22753 35479
rect 22753 35445 22787 35479
rect 22787 35445 22796 35479
rect 22744 35436 22796 35445
rect 23756 35479 23808 35488
rect 23756 35445 23765 35479
rect 23765 35445 23799 35479
rect 23799 35445 23808 35479
rect 23756 35436 23808 35445
rect 24032 35436 24084 35488
rect 24676 35436 24728 35488
rect 26240 35436 26292 35488
rect 28448 35504 28500 35556
rect 27988 35436 28040 35488
rect 38200 35479 38252 35488
rect 38200 35445 38209 35479
rect 38209 35445 38243 35479
rect 38243 35445 38252 35479
rect 38200 35436 38252 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 3976 35232 4028 35284
rect 3792 35164 3844 35216
rect 7196 35232 7248 35284
rect 7656 35232 7708 35284
rect 7840 35232 7892 35284
rect 13084 35232 13136 35284
rect 14188 35232 14240 35284
rect 19800 35232 19852 35284
rect 3424 35139 3476 35148
rect 3424 35105 3433 35139
rect 3433 35105 3467 35139
rect 3467 35105 3476 35139
rect 3424 35096 3476 35105
rect 3884 35096 3936 35148
rect 9404 35164 9456 35216
rect 14372 35164 14424 35216
rect 19064 35164 19116 35216
rect 25688 35275 25740 35284
rect 25688 35241 25697 35275
rect 25697 35241 25731 35275
rect 25731 35241 25740 35275
rect 25688 35232 25740 35241
rect 26240 35275 26292 35284
rect 26240 35241 26249 35275
rect 26249 35241 26283 35275
rect 26283 35241 26292 35275
rect 26240 35232 26292 35241
rect 21364 35164 21416 35216
rect 22836 35164 22888 35216
rect 11060 35096 11112 35148
rect 2044 35028 2096 35080
rect 3700 35028 3752 35080
rect 3976 35071 4028 35080
rect 3976 35037 3985 35071
rect 3985 35037 4019 35071
rect 4019 35037 4028 35071
rect 3976 35028 4028 35037
rect 8576 35071 8628 35080
rect 8576 35037 8585 35071
rect 8585 35037 8619 35071
rect 8619 35037 8628 35071
rect 9128 35071 9180 35080
rect 8576 35028 8628 35037
rect 9128 35037 9137 35071
rect 9137 35037 9171 35071
rect 9171 35037 9180 35071
rect 9128 35028 9180 35037
rect 15660 35096 15712 35148
rect 13268 35071 13320 35080
rect 5172 34960 5224 35012
rect 2412 34892 2464 34944
rect 3976 34892 4028 34944
rect 5632 34892 5684 34944
rect 6552 34892 6604 34944
rect 7840 34960 7892 35012
rect 8208 34892 8260 34944
rect 8668 34960 8720 35012
rect 13268 35037 13277 35071
rect 13277 35037 13311 35071
rect 13311 35037 13320 35071
rect 13268 35028 13320 35037
rect 13820 35028 13872 35080
rect 15016 35071 15068 35080
rect 15016 35037 15025 35071
rect 15025 35037 15059 35071
rect 15059 35037 15068 35071
rect 15016 35028 15068 35037
rect 15384 35028 15436 35080
rect 9496 34960 9548 35012
rect 12256 34960 12308 35012
rect 8484 34892 8536 34944
rect 8760 34892 8812 34944
rect 12348 34892 12400 34944
rect 12532 34892 12584 34944
rect 13728 34960 13780 35012
rect 19432 35096 19484 35148
rect 20076 35139 20128 35148
rect 20076 35105 20085 35139
rect 20085 35105 20119 35139
rect 20119 35105 20128 35139
rect 20076 35096 20128 35105
rect 25780 35164 25832 35216
rect 25136 35139 25188 35148
rect 16396 35028 16448 35080
rect 16856 35028 16908 35080
rect 17316 35071 17368 35080
rect 17316 35037 17325 35071
rect 17325 35037 17359 35071
rect 17359 35037 17368 35071
rect 17316 35028 17368 35037
rect 15844 34960 15896 35012
rect 16488 34960 16540 35012
rect 18696 35028 18748 35080
rect 18052 34960 18104 35012
rect 19064 34960 19116 35012
rect 19984 34960 20036 35012
rect 21088 35028 21140 35080
rect 25136 35105 25145 35139
rect 25145 35105 25179 35139
rect 25179 35105 25188 35139
rect 25136 35096 25188 35105
rect 20996 34960 21048 35012
rect 23204 34960 23256 35012
rect 14280 34935 14332 34944
rect 14280 34901 14289 34935
rect 14289 34901 14323 34935
rect 14323 34901 14332 34935
rect 14280 34892 14332 34901
rect 15016 34892 15068 34944
rect 16028 34892 16080 34944
rect 16396 34892 16448 34944
rect 22376 34935 22428 34944
rect 22376 34901 22385 34935
rect 22385 34901 22419 34935
rect 22419 34901 22428 34935
rect 22376 34892 22428 34901
rect 24032 34935 24084 34944
rect 24032 34901 24041 34935
rect 24041 34901 24075 34935
rect 24075 34901 24084 34935
rect 24032 34892 24084 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 3792 34688 3844 34740
rect 3884 34688 3936 34740
rect 3148 34620 3200 34672
rect 3700 34620 3752 34672
rect 4620 34620 4672 34672
rect 5540 34595 5592 34604
rect 5540 34561 5549 34595
rect 5549 34561 5583 34595
rect 5583 34561 5592 34595
rect 5540 34552 5592 34561
rect 1952 34484 2004 34536
rect 3700 34484 3752 34536
rect 7196 34620 7248 34672
rect 5816 34552 5868 34604
rect 8208 34688 8260 34740
rect 8852 34688 8904 34740
rect 10692 34688 10744 34740
rect 12164 34688 12216 34740
rect 6920 34484 6972 34536
rect 7288 34484 7340 34536
rect 8208 34484 8260 34536
rect 8944 34527 8996 34536
rect 8944 34493 8953 34527
rect 8953 34493 8987 34527
rect 8987 34493 8996 34527
rect 8944 34484 8996 34493
rect 7932 34416 7984 34468
rect 5264 34391 5316 34400
rect 5264 34357 5285 34391
rect 5285 34357 5316 34391
rect 5264 34348 5316 34357
rect 5448 34348 5500 34400
rect 7012 34348 7064 34400
rect 7564 34348 7616 34400
rect 7840 34348 7892 34400
rect 8576 34348 8628 34400
rect 9680 34620 9732 34672
rect 13268 34620 13320 34672
rect 9864 34595 9916 34604
rect 9864 34561 9873 34595
rect 9873 34561 9907 34595
rect 9907 34561 9916 34595
rect 10508 34595 10560 34604
rect 9864 34552 9916 34561
rect 10508 34561 10517 34595
rect 10517 34561 10551 34595
rect 10551 34561 10560 34595
rect 11152 34595 11204 34604
rect 10508 34552 10560 34561
rect 11152 34561 11161 34595
rect 11161 34561 11195 34595
rect 11195 34561 11204 34595
rect 11152 34552 11204 34561
rect 14280 34688 14332 34740
rect 14372 34688 14424 34740
rect 15108 34688 15160 34740
rect 15660 34688 15712 34740
rect 19248 34688 19300 34740
rect 21364 34731 21416 34740
rect 21364 34697 21373 34731
rect 21373 34697 21407 34731
rect 21407 34697 21416 34731
rect 21364 34688 21416 34697
rect 22744 34688 22796 34740
rect 14096 34620 14148 34672
rect 17408 34663 17460 34672
rect 13544 34552 13596 34604
rect 14648 34552 14700 34604
rect 14832 34595 14884 34604
rect 14832 34561 14841 34595
rect 14841 34561 14875 34595
rect 14875 34561 14884 34595
rect 14832 34552 14884 34561
rect 15292 34552 15344 34604
rect 9404 34484 9456 34536
rect 13084 34484 13136 34536
rect 13636 34484 13688 34536
rect 14556 34484 14608 34536
rect 15660 34484 15712 34536
rect 15752 34484 15804 34536
rect 17408 34629 17417 34663
rect 17417 34629 17451 34663
rect 17451 34629 17460 34663
rect 17408 34620 17460 34629
rect 17684 34620 17736 34672
rect 17868 34620 17920 34672
rect 16856 34595 16908 34604
rect 16856 34561 16865 34595
rect 16865 34561 16899 34595
rect 16899 34561 16908 34595
rect 16856 34552 16908 34561
rect 18972 34595 19024 34604
rect 18972 34561 18981 34595
rect 18981 34561 19015 34595
rect 19015 34561 19024 34595
rect 18972 34552 19024 34561
rect 19984 34552 20036 34604
rect 21824 34620 21876 34672
rect 23204 34663 23256 34672
rect 23204 34629 23213 34663
rect 23213 34629 23247 34663
rect 23247 34629 23256 34663
rect 29000 34688 29052 34740
rect 23204 34620 23256 34629
rect 24308 34527 24360 34536
rect 9312 34348 9364 34400
rect 9680 34348 9732 34400
rect 11612 34348 11664 34400
rect 11980 34348 12032 34400
rect 19432 34416 19484 34468
rect 24308 34493 24317 34527
rect 24317 34493 24351 34527
rect 24351 34493 24360 34527
rect 37740 34620 37792 34672
rect 24308 34484 24360 34493
rect 24032 34416 24084 34468
rect 25688 34416 25740 34468
rect 15200 34348 15252 34400
rect 15384 34348 15436 34400
rect 20720 34348 20772 34400
rect 20812 34391 20864 34400
rect 20812 34357 20821 34391
rect 20821 34357 20855 34391
rect 20855 34357 20864 34391
rect 23664 34391 23716 34400
rect 20812 34348 20864 34357
rect 23664 34357 23673 34391
rect 23673 34357 23707 34391
rect 23707 34357 23716 34391
rect 23664 34348 23716 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 2504 34144 2556 34196
rect 2964 34008 3016 34060
rect 3424 34008 3476 34060
rect 1124 33804 1176 33856
rect 3424 33847 3476 33856
rect 3424 33813 3433 33847
rect 3433 33813 3467 33847
rect 3467 33813 3476 33847
rect 3424 33804 3476 33813
rect 5080 34144 5132 34196
rect 5264 34144 5316 34196
rect 7656 34144 7708 34196
rect 7840 34144 7892 34196
rect 8300 34144 8352 34196
rect 9772 34187 9824 34196
rect 9772 34153 9781 34187
rect 9781 34153 9815 34187
rect 9815 34153 9824 34187
rect 9772 34144 9824 34153
rect 4804 33940 4856 33992
rect 5540 34008 5592 34060
rect 9588 34076 9640 34128
rect 10784 34076 10836 34128
rect 12348 34144 12400 34196
rect 14280 34144 14332 34196
rect 14372 34144 14424 34196
rect 21732 34144 21784 34196
rect 4988 33940 5040 33992
rect 5448 33940 5500 33992
rect 5632 33940 5684 33992
rect 7472 33940 7524 33992
rect 7748 33940 7800 33992
rect 7932 33940 7984 33992
rect 11152 34008 11204 34060
rect 12164 34051 12216 34060
rect 12164 34017 12173 34051
rect 12173 34017 12207 34051
rect 12207 34017 12216 34051
rect 12164 34008 12216 34017
rect 12440 34076 12492 34128
rect 8300 33940 8352 33992
rect 9956 33940 10008 33992
rect 10600 33940 10652 33992
rect 5632 33804 5684 33856
rect 7012 33872 7064 33924
rect 8760 33872 8812 33924
rect 11428 33872 11480 33924
rect 11796 33872 11848 33924
rect 7932 33847 7984 33856
rect 7932 33813 7941 33847
rect 7941 33813 7975 33847
rect 7975 33813 7984 33847
rect 7932 33804 7984 33813
rect 11520 33804 11572 33856
rect 11612 33804 11664 33856
rect 13268 33940 13320 33992
rect 13544 33940 13596 33992
rect 12440 33872 12492 33924
rect 15200 33940 15252 33992
rect 16488 34008 16540 34060
rect 19524 34051 19576 34060
rect 17224 33940 17276 33992
rect 17868 33940 17920 33992
rect 14924 33872 14976 33924
rect 15016 33872 15068 33924
rect 15844 33872 15896 33924
rect 16120 33872 16172 33924
rect 16488 33915 16540 33924
rect 16488 33881 16497 33915
rect 16497 33881 16531 33915
rect 16531 33881 16540 33915
rect 16488 33872 16540 33881
rect 13728 33804 13780 33856
rect 14280 33804 14332 33856
rect 17224 33804 17276 33856
rect 17500 33872 17552 33924
rect 17960 33872 18012 33924
rect 18144 33915 18196 33924
rect 18144 33881 18153 33915
rect 18153 33881 18187 33915
rect 18187 33881 18196 33915
rect 18144 33872 18196 33881
rect 18236 33915 18288 33924
rect 18236 33881 18245 33915
rect 18245 33881 18279 33915
rect 18279 33881 18288 33915
rect 18788 33915 18840 33924
rect 18236 33872 18288 33881
rect 18788 33881 18797 33915
rect 18797 33881 18831 33915
rect 18831 33881 18840 33915
rect 18788 33872 18840 33881
rect 17684 33804 17736 33856
rect 19524 34017 19533 34051
rect 19533 34017 19567 34051
rect 19567 34017 19576 34051
rect 19524 34008 19576 34017
rect 20536 34076 20588 34128
rect 20720 34076 20772 34128
rect 22836 34144 22888 34196
rect 23204 34187 23256 34196
rect 23204 34153 23213 34187
rect 23213 34153 23247 34187
rect 23247 34153 23256 34187
rect 23204 34144 23256 34153
rect 25688 34187 25740 34196
rect 25688 34153 25697 34187
rect 25697 34153 25731 34187
rect 25731 34153 25740 34187
rect 25688 34144 25740 34153
rect 26332 34144 26384 34196
rect 37464 34144 37516 34196
rect 25412 34076 25464 34128
rect 19984 33983 20036 33992
rect 19984 33949 19993 33983
rect 19993 33949 20027 33983
rect 20027 33949 20036 33983
rect 19984 33940 20036 33949
rect 20812 33940 20864 33992
rect 25228 33940 25280 33992
rect 25412 33940 25464 33992
rect 38016 34076 38068 34128
rect 20536 33872 20588 33924
rect 20904 33847 20956 33856
rect 20904 33813 20913 33847
rect 20913 33813 20947 33847
rect 20947 33813 20956 33847
rect 20904 33804 20956 33813
rect 22100 33847 22152 33856
rect 22100 33813 22109 33847
rect 22109 33813 22143 33847
rect 22143 33813 22152 33847
rect 22100 33804 22152 33813
rect 22744 33872 22796 33924
rect 23664 33847 23716 33856
rect 23664 33813 23673 33847
rect 23673 33813 23707 33847
rect 23707 33813 23716 33847
rect 23664 33804 23716 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 1032 33464 1084 33516
rect 2780 33532 2832 33584
rect 4620 33532 4672 33584
rect 5908 33532 5960 33584
rect 7288 33575 7340 33584
rect 7288 33541 7297 33575
rect 7297 33541 7331 33575
rect 7331 33541 7340 33575
rect 7288 33532 7340 33541
rect 7932 33532 7984 33584
rect 11428 33600 11480 33652
rect 14372 33600 14424 33652
rect 14464 33600 14516 33652
rect 19248 33600 19300 33652
rect 19432 33600 19484 33652
rect 23204 33600 23256 33652
rect 25228 33600 25280 33652
rect 12256 33532 12308 33584
rect 13452 33532 13504 33584
rect 13544 33532 13596 33584
rect 15844 33532 15896 33584
rect 16028 33575 16080 33584
rect 16028 33541 16037 33575
rect 16037 33541 16071 33575
rect 16071 33541 16080 33575
rect 16028 33532 16080 33541
rect 17500 33532 17552 33584
rect 17868 33532 17920 33584
rect 2872 33464 2924 33516
rect 3424 33464 3476 33516
rect 5540 33507 5592 33516
rect 5540 33473 5549 33507
rect 5549 33473 5583 33507
rect 5583 33473 5592 33507
rect 5540 33464 5592 33473
rect 9312 33507 9364 33516
rect 9312 33473 9321 33507
rect 9321 33473 9355 33507
rect 9355 33473 9364 33507
rect 9312 33464 9364 33473
rect 9680 33396 9732 33448
rect 9956 33396 10008 33448
rect 11060 33464 11112 33516
rect 14372 33464 14424 33516
rect 11980 33439 12032 33448
rect 11980 33405 11989 33439
rect 11989 33405 12023 33439
rect 12023 33405 12032 33439
rect 11980 33396 12032 33405
rect 13176 33396 13228 33448
rect 16672 33464 16724 33516
rect 17960 33507 18012 33516
rect 17960 33473 17969 33507
rect 17969 33473 18003 33507
rect 18003 33473 18012 33507
rect 17960 33464 18012 33473
rect 18972 33507 19024 33516
rect 18972 33473 18981 33507
rect 18981 33473 19015 33507
rect 19015 33473 19024 33507
rect 18972 33464 19024 33473
rect 19340 33464 19392 33516
rect 20812 33532 20864 33584
rect 20628 33507 20680 33516
rect 20628 33473 20637 33507
rect 20637 33473 20671 33507
rect 20671 33473 20680 33507
rect 20628 33464 20680 33473
rect 22836 33464 22888 33516
rect 26424 33507 26476 33516
rect 26424 33473 26433 33507
rect 26433 33473 26467 33507
rect 26467 33473 26476 33507
rect 26424 33464 26476 33473
rect 38200 33507 38252 33516
rect 38200 33473 38209 33507
rect 38209 33473 38243 33507
rect 38243 33473 38252 33507
rect 38200 33464 38252 33473
rect 15844 33439 15896 33448
rect 15844 33405 15853 33439
rect 15853 33405 15887 33439
rect 15887 33405 15896 33439
rect 15844 33396 15896 33405
rect 15936 33396 15988 33448
rect 20720 33396 20772 33448
rect 3792 33303 3844 33312
rect 3792 33269 3801 33303
rect 3801 33269 3835 33303
rect 3835 33269 3844 33303
rect 3792 33260 3844 33269
rect 7840 33260 7892 33312
rect 7932 33260 7984 33312
rect 9312 33260 9364 33312
rect 11336 33260 11388 33312
rect 14464 33260 14516 33312
rect 14740 33260 14792 33312
rect 15568 33328 15620 33380
rect 25872 33371 25924 33380
rect 25872 33337 25881 33371
rect 25881 33337 25915 33371
rect 25915 33337 25924 33371
rect 25872 33328 25924 33337
rect 37372 33328 37424 33380
rect 16488 33260 16540 33312
rect 17868 33260 17920 33312
rect 18604 33260 18656 33312
rect 22100 33303 22152 33312
rect 22100 33269 22109 33303
rect 22109 33269 22143 33303
rect 22143 33269 22152 33303
rect 22100 33260 22152 33269
rect 24032 33260 24084 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 3332 33056 3384 33108
rect 7012 33056 7064 33108
rect 7288 33056 7340 33108
rect 11152 33056 11204 33108
rect 5540 32988 5592 33040
rect 7104 32988 7156 33040
rect 16396 33056 16448 33108
rect 16580 33056 16632 33108
rect 17408 33056 17460 33108
rect 19248 33056 19300 33108
rect 20904 33056 20956 33108
rect 21732 33099 21784 33108
rect 21732 33065 21741 33099
rect 21741 33065 21775 33099
rect 21775 33065 21784 33099
rect 21732 33056 21784 33065
rect 23204 33056 23256 33108
rect 23664 33056 23716 33108
rect 25228 33099 25280 33108
rect 25228 33065 25237 33099
rect 25237 33065 25271 33099
rect 25271 33065 25280 33099
rect 25228 33056 25280 33065
rect 12624 32988 12676 33040
rect 22192 32988 22244 33040
rect 2964 32920 3016 32972
rect 5448 32920 5500 32972
rect 7288 32920 7340 32972
rect 4988 32852 5040 32904
rect 7472 32852 7524 32904
rect 8300 32852 8352 32904
rect 8852 32852 8904 32904
rect 9312 32852 9364 32904
rect 11060 32920 11112 32972
rect 11520 32963 11572 32972
rect 11520 32929 11529 32963
rect 11529 32929 11563 32963
rect 11563 32929 11572 32963
rect 11520 32920 11572 32929
rect 12164 32920 12216 32972
rect 13452 32920 13504 32972
rect 14280 32920 14332 32972
rect 16120 32920 16172 32972
rect 16580 32963 16632 32972
rect 16580 32929 16589 32963
rect 16589 32929 16623 32963
rect 16623 32929 16632 32963
rect 16580 32920 16632 32929
rect 16948 32963 17000 32972
rect 16948 32929 16957 32963
rect 16957 32929 16991 32963
rect 16991 32929 17000 32963
rect 16948 32920 17000 32929
rect 17224 32920 17276 32972
rect 20720 32920 20772 32972
rect 12624 32852 12676 32904
rect 13360 32852 13412 32904
rect 14648 32852 14700 32904
rect 18328 32895 18380 32904
rect 18328 32861 18337 32895
rect 18337 32861 18371 32895
rect 18371 32861 18380 32895
rect 18328 32852 18380 32861
rect 19340 32852 19392 32904
rect 20628 32852 20680 32904
rect 22284 32852 22336 32904
rect 25688 32895 25740 32904
rect 25688 32861 25697 32895
rect 25697 32861 25731 32895
rect 25731 32861 25740 32895
rect 25688 32852 25740 32861
rect 1216 32716 1268 32768
rect 5632 32784 5684 32836
rect 6644 32827 6696 32836
rect 6644 32793 6653 32827
rect 6653 32793 6687 32827
rect 6687 32793 6696 32827
rect 6644 32784 6696 32793
rect 11428 32784 11480 32836
rect 13268 32827 13320 32836
rect 13268 32793 13277 32827
rect 13277 32793 13311 32827
rect 13311 32793 13320 32827
rect 13268 32784 13320 32793
rect 6000 32716 6052 32768
rect 7748 32716 7800 32768
rect 8484 32759 8536 32768
rect 8484 32725 8493 32759
rect 8493 32725 8527 32759
rect 8527 32725 8536 32759
rect 8484 32716 8536 32725
rect 9220 32759 9272 32768
rect 9220 32725 9229 32759
rect 9229 32725 9263 32759
rect 9263 32725 9272 32759
rect 9220 32716 9272 32725
rect 9496 32716 9548 32768
rect 10508 32716 10560 32768
rect 10692 32759 10744 32768
rect 10692 32725 10701 32759
rect 10701 32725 10735 32759
rect 10735 32725 10744 32759
rect 10692 32716 10744 32725
rect 12256 32716 12308 32768
rect 14740 32784 14792 32836
rect 16396 32784 16448 32836
rect 16580 32716 16632 32768
rect 16764 32784 16816 32836
rect 20076 32784 20128 32836
rect 17040 32716 17092 32768
rect 18512 32716 18564 32768
rect 20352 32716 20404 32768
rect 22100 32716 22152 32768
rect 24032 32759 24084 32768
rect 24032 32725 24041 32759
rect 24041 32725 24075 32759
rect 24075 32725 24084 32759
rect 24032 32716 24084 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 1676 32419 1728 32428
rect 1676 32385 1685 32419
rect 1685 32385 1719 32419
rect 1719 32385 1728 32419
rect 1676 32376 1728 32385
rect 2596 32419 2648 32428
rect 2596 32385 2605 32419
rect 2605 32385 2639 32419
rect 2639 32385 2648 32419
rect 2596 32376 2648 32385
rect 2964 32512 3016 32564
rect 2872 32444 2924 32496
rect 5080 32512 5132 32564
rect 5540 32512 5592 32564
rect 7012 32512 7064 32564
rect 3516 32444 3568 32496
rect 7748 32444 7800 32496
rect 9036 32444 9088 32496
rect 11612 32444 11664 32496
rect 11152 32376 11204 32428
rect 12900 32512 12952 32564
rect 15384 32512 15436 32564
rect 16856 32512 16908 32564
rect 12992 32444 13044 32496
rect 2320 32240 2372 32292
rect 3700 32283 3752 32292
rect 3700 32249 3709 32283
rect 3709 32249 3743 32283
rect 3743 32249 3752 32283
rect 3700 32240 3752 32249
rect 3884 32308 3936 32360
rect 8392 32308 8444 32360
rect 8760 32351 8812 32360
rect 8760 32317 8769 32351
rect 8769 32317 8803 32351
rect 8803 32317 8812 32351
rect 9404 32351 9456 32360
rect 8760 32308 8812 32317
rect 9404 32317 9413 32351
rect 9413 32317 9447 32351
rect 9447 32317 9456 32351
rect 9404 32308 9456 32317
rect 5448 32240 5500 32292
rect 7104 32240 7156 32292
rect 12072 32308 12124 32360
rect 11520 32240 11572 32292
rect 12808 32308 12860 32360
rect 15108 32444 15160 32496
rect 22192 32512 22244 32564
rect 18328 32487 18380 32496
rect 18328 32453 18337 32487
rect 18337 32453 18371 32487
rect 18371 32453 18380 32487
rect 18328 32444 18380 32453
rect 18696 32444 18748 32496
rect 18788 32444 18840 32496
rect 19432 32376 19484 32428
rect 19984 32376 20036 32428
rect 20260 32419 20312 32428
rect 20260 32385 20269 32419
rect 20269 32385 20303 32419
rect 20303 32385 20312 32419
rect 20260 32376 20312 32385
rect 20904 32376 20956 32428
rect 22192 32419 22244 32428
rect 22192 32385 22201 32419
rect 22201 32385 22235 32419
rect 22235 32385 22244 32419
rect 22192 32376 22244 32385
rect 38016 32419 38068 32428
rect 38016 32385 38025 32419
rect 38025 32385 38059 32419
rect 38059 32385 38068 32419
rect 38016 32376 38068 32385
rect 10968 32172 11020 32224
rect 12072 32172 12124 32224
rect 15200 32308 15252 32360
rect 17500 32351 17552 32360
rect 17500 32317 17509 32351
rect 17509 32317 17543 32351
rect 17543 32317 17552 32351
rect 17500 32308 17552 32317
rect 17960 32308 18012 32360
rect 20720 32351 20772 32360
rect 20720 32317 20729 32351
rect 20729 32317 20763 32351
rect 20763 32317 20772 32351
rect 20720 32308 20772 32317
rect 22100 32308 22152 32360
rect 24032 32308 24084 32360
rect 18420 32240 18472 32292
rect 22284 32172 22336 32224
rect 38200 32215 38252 32224
rect 38200 32181 38209 32215
rect 38209 32181 38243 32215
rect 38243 32181 38252 32215
rect 38200 32172 38252 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 2780 31968 2832 32020
rect 2964 31968 3016 32020
rect 3424 31968 3476 32020
rect 7104 31968 7156 32020
rect 7288 31968 7340 32020
rect 9312 31968 9364 32020
rect 7564 31900 7616 31952
rect 10232 31968 10284 32020
rect 3608 31832 3660 31884
rect 5540 31832 5592 31884
rect 8760 31832 8812 31884
rect 3424 31807 3476 31816
rect 3424 31773 3433 31807
rect 3433 31773 3467 31807
rect 3467 31773 3476 31807
rect 3424 31764 3476 31773
rect 5448 31764 5500 31816
rect 6000 31764 6052 31816
rect 2136 31696 2188 31748
rect 5632 31696 5684 31748
rect 7196 31696 7248 31748
rect 9312 31764 9364 31816
rect 12072 31968 12124 32020
rect 12440 31968 12492 32020
rect 13452 31968 13504 32020
rect 13544 31968 13596 32020
rect 15384 31968 15436 32020
rect 15568 31968 15620 32020
rect 20812 31968 20864 32020
rect 21824 31968 21876 32020
rect 22100 31968 22152 32020
rect 13636 31900 13688 31952
rect 9588 31764 9640 31816
rect 10600 31832 10652 31884
rect 11060 31832 11112 31884
rect 12992 31832 13044 31884
rect 13360 31832 13412 31884
rect 10140 31807 10192 31816
rect 10140 31773 10149 31807
rect 10149 31773 10183 31807
rect 10183 31773 10192 31807
rect 13636 31807 13688 31816
rect 10140 31764 10192 31773
rect 13636 31773 13645 31807
rect 13645 31773 13679 31807
rect 13679 31773 13688 31807
rect 13636 31764 13688 31773
rect 14004 31832 14056 31884
rect 14648 31832 14700 31884
rect 16028 31900 16080 31952
rect 16396 31943 16448 31952
rect 16396 31909 16405 31943
rect 16405 31909 16439 31943
rect 16439 31909 16448 31943
rect 16396 31900 16448 31909
rect 16948 31900 17000 31952
rect 20168 31900 20220 31952
rect 22836 31943 22888 31952
rect 22836 31909 22845 31943
rect 22845 31909 22879 31943
rect 22879 31909 22888 31943
rect 22836 31900 22888 31909
rect 15384 31875 15436 31884
rect 15384 31841 15393 31875
rect 15393 31841 15427 31875
rect 15427 31841 15436 31875
rect 15752 31875 15804 31884
rect 15384 31832 15436 31841
rect 15752 31841 15761 31875
rect 15761 31841 15795 31875
rect 15795 31841 15804 31875
rect 15752 31832 15804 31841
rect 16580 31832 16632 31884
rect 17592 31832 17644 31884
rect 17960 31832 18012 31884
rect 18788 31807 18840 31816
rect 18788 31773 18797 31807
rect 18797 31773 18831 31807
rect 18831 31773 18840 31807
rect 18788 31764 18840 31773
rect 19432 31764 19484 31816
rect 4252 31628 4304 31680
rect 6092 31628 6144 31680
rect 9496 31696 9548 31748
rect 8576 31628 8628 31680
rect 11336 31628 11388 31680
rect 12256 31739 12308 31748
rect 12256 31705 12265 31739
rect 12265 31705 12299 31739
rect 12299 31705 12308 31739
rect 12256 31696 12308 31705
rect 13912 31696 13964 31748
rect 15660 31739 15712 31748
rect 15660 31705 15669 31739
rect 15669 31705 15703 31739
rect 15703 31705 15712 31739
rect 15660 31696 15712 31705
rect 16764 31696 16816 31748
rect 17592 31739 17644 31748
rect 12532 31628 12584 31680
rect 14188 31628 14240 31680
rect 16580 31628 16632 31680
rect 17592 31705 17601 31739
rect 17601 31705 17635 31739
rect 17635 31705 17644 31739
rect 17592 31696 17644 31705
rect 17684 31739 17736 31748
rect 17684 31705 17693 31739
rect 17693 31705 17727 31739
rect 17727 31705 17736 31739
rect 18236 31739 18288 31748
rect 17684 31696 17736 31705
rect 18236 31705 18245 31739
rect 18245 31705 18279 31739
rect 18279 31705 18288 31739
rect 18236 31696 18288 31705
rect 19340 31696 19392 31748
rect 20076 31764 20128 31816
rect 19984 31696 20036 31748
rect 20720 31764 20772 31816
rect 22192 31832 22244 31884
rect 17500 31628 17552 31680
rect 20904 31628 20956 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 8300 31424 8352 31476
rect 10692 31424 10744 31476
rect 3148 31356 3200 31408
rect 4252 31356 4304 31408
rect 8484 31356 8536 31408
rect 8852 31356 8904 31408
rect 1676 31331 1728 31340
rect 1676 31297 1685 31331
rect 1685 31297 1719 31331
rect 1719 31297 1728 31331
rect 1676 31288 1728 31297
rect 2228 31288 2280 31340
rect 2596 31288 2648 31340
rect 5448 31288 5500 31340
rect 7472 31288 7524 31340
rect 9404 31331 9456 31340
rect 9404 31297 9413 31331
rect 9413 31297 9447 31331
rect 9447 31297 9456 31331
rect 11704 31356 11756 31408
rect 12716 31356 12768 31408
rect 13176 31356 13228 31408
rect 9404 31288 9456 31297
rect 10876 31288 10928 31340
rect 17316 31399 17368 31408
rect 17316 31365 17325 31399
rect 17325 31365 17359 31399
rect 17359 31365 17368 31399
rect 17316 31356 17368 31365
rect 18236 31356 18288 31408
rect 18512 31399 18564 31408
rect 18512 31365 18521 31399
rect 18521 31365 18555 31399
rect 18555 31365 18564 31399
rect 18512 31356 18564 31365
rect 19156 31424 19208 31476
rect 19248 31424 19300 31476
rect 20352 31424 20404 31476
rect 20904 31467 20956 31476
rect 20904 31433 20913 31467
rect 20913 31433 20947 31467
rect 20947 31433 20956 31467
rect 20904 31424 20956 31433
rect 22100 31467 22152 31476
rect 22100 31433 22109 31467
rect 22109 31433 22143 31467
rect 22143 31433 22152 31467
rect 22560 31467 22612 31476
rect 22100 31424 22152 31433
rect 22560 31433 22569 31467
rect 22569 31433 22603 31467
rect 22603 31433 22612 31467
rect 22560 31424 22612 31433
rect 23664 31424 23716 31476
rect 19340 31356 19392 31408
rect 20260 31356 20312 31408
rect 14280 31288 14332 31340
rect 16028 31331 16080 31340
rect 16028 31297 16037 31331
rect 16037 31297 16071 31331
rect 16071 31297 16080 31331
rect 16028 31288 16080 31297
rect 19432 31288 19484 31340
rect 19984 31288 20036 31340
rect 3976 31220 4028 31272
rect 1860 31195 1912 31204
rect 1860 31161 1869 31195
rect 1869 31161 1903 31195
rect 1903 31161 1912 31195
rect 1860 31152 1912 31161
rect 6000 31220 6052 31272
rect 9128 31263 9180 31272
rect 9128 31229 9137 31263
rect 9137 31229 9171 31263
rect 9171 31229 9180 31263
rect 9128 31220 9180 31229
rect 11336 31220 11388 31272
rect 11704 31220 11756 31272
rect 13176 31220 13228 31272
rect 13268 31263 13320 31272
rect 13268 31229 13277 31263
rect 13277 31229 13311 31263
rect 13311 31229 13320 31263
rect 13268 31220 13320 31229
rect 7748 31152 7800 31204
rect 2320 31127 2372 31136
rect 2320 31093 2329 31127
rect 2329 31093 2363 31127
rect 2363 31093 2372 31127
rect 2320 31084 2372 31093
rect 5172 31084 5224 31136
rect 5448 31084 5500 31136
rect 10968 31152 11020 31204
rect 10416 31127 10468 31136
rect 10416 31093 10425 31127
rect 10425 31093 10459 31127
rect 10459 31093 10468 31127
rect 10416 31084 10468 31093
rect 11612 31084 11664 31136
rect 12808 31084 12860 31136
rect 13084 31084 13136 31136
rect 15016 31220 15068 31272
rect 15200 31263 15252 31272
rect 15200 31229 15209 31263
rect 15209 31229 15243 31263
rect 15243 31229 15252 31263
rect 15200 31220 15252 31229
rect 15844 31220 15896 31272
rect 17224 31263 17276 31272
rect 17224 31229 17233 31263
rect 17233 31229 17267 31263
rect 17267 31229 17276 31263
rect 17224 31220 17276 31229
rect 20444 31220 20496 31272
rect 13912 31152 13964 31204
rect 15292 31084 15344 31136
rect 15384 31084 15436 31136
rect 16212 31084 16264 31136
rect 18144 31084 18196 31136
rect 19432 31084 19484 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 4804 30880 4856 30932
rect 5264 30880 5316 30932
rect 7656 30880 7708 30932
rect 4712 30744 4764 30796
rect 4896 30744 4948 30796
rect 5632 30744 5684 30796
rect 8760 30812 8812 30864
rect 9404 30880 9456 30932
rect 11060 30880 11112 30932
rect 11244 30880 11296 30932
rect 12348 30880 12400 30932
rect 12716 30880 12768 30932
rect 20168 30923 20220 30932
rect 9404 30744 9456 30796
rect 9864 30812 9916 30864
rect 10508 30812 10560 30864
rect 10876 30812 10928 30864
rect 16212 30855 16264 30864
rect 16212 30821 16221 30855
rect 16221 30821 16255 30855
rect 16255 30821 16264 30855
rect 16212 30812 16264 30821
rect 17960 30812 18012 30864
rect 20168 30889 20177 30923
rect 20177 30889 20211 30923
rect 20211 30889 20220 30923
rect 20168 30880 20220 30889
rect 20720 30923 20772 30932
rect 20720 30889 20729 30923
rect 20729 30889 20763 30923
rect 20763 30889 20772 30923
rect 20720 30880 20772 30889
rect 37280 30812 37332 30864
rect 3424 30719 3476 30728
rect 3424 30685 3433 30719
rect 3433 30685 3467 30719
rect 3467 30685 3476 30719
rect 3976 30719 4028 30728
rect 3424 30676 3476 30685
rect 3976 30685 3985 30719
rect 3985 30685 4019 30719
rect 4019 30685 4028 30719
rect 3976 30676 4028 30685
rect 5908 30676 5960 30728
rect 6184 30676 6236 30728
rect 9956 30676 10008 30728
rect 10416 30744 10468 30796
rect 15016 30787 15068 30796
rect 11244 30676 11296 30728
rect 12992 30719 13044 30728
rect 12992 30685 13001 30719
rect 13001 30685 13035 30719
rect 13035 30685 13044 30719
rect 12992 30676 13044 30685
rect 13176 30676 13228 30728
rect 2504 30608 2556 30660
rect 1768 30540 1820 30592
rect 3240 30540 3292 30592
rect 5264 30608 5316 30660
rect 5632 30540 5684 30592
rect 6920 30608 6972 30660
rect 8576 30608 8628 30660
rect 9588 30608 9640 30660
rect 8852 30540 8904 30592
rect 12256 30608 12308 30660
rect 12808 30608 12860 30660
rect 13268 30608 13320 30660
rect 15016 30753 15025 30787
rect 15025 30753 15059 30787
rect 15059 30753 15068 30787
rect 15016 30744 15068 30753
rect 16304 30744 16356 30796
rect 14280 30719 14332 30728
rect 14280 30685 14289 30719
rect 14289 30685 14323 30719
rect 14323 30685 14332 30719
rect 14280 30676 14332 30685
rect 18420 30676 18472 30728
rect 20352 30744 20404 30796
rect 20260 30719 20312 30728
rect 20260 30685 20269 30719
rect 20269 30685 20303 30719
rect 20303 30685 20312 30719
rect 20260 30676 20312 30685
rect 22192 30676 22244 30728
rect 15844 30608 15896 30660
rect 13084 30540 13136 30592
rect 14188 30540 14240 30592
rect 14280 30540 14332 30592
rect 15016 30540 15068 30592
rect 16120 30540 16172 30592
rect 16764 30651 16816 30660
rect 16764 30617 16773 30651
rect 16773 30617 16807 30651
rect 16807 30617 16816 30651
rect 16764 30608 16816 30617
rect 17592 30608 17644 30660
rect 17868 30651 17920 30660
rect 17868 30617 17877 30651
rect 17877 30617 17911 30651
rect 17911 30617 17920 30651
rect 17868 30608 17920 30617
rect 20812 30608 20864 30660
rect 21824 30540 21876 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 7288 30336 7340 30388
rect 7656 30336 7708 30388
rect 9128 30336 9180 30388
rect 3700 30268 3752 30320
rect 5264 30268 5316 30320
rect 6000 30268 6052 30320
rect 8300 30268 8352 30320
rect 9220 30268 9272 30320
rect 12256 30336 12308 30388
rect 21824 30336 21876 30388
rect 11336 30268 11388 30320
rect 12716 30268 12768 30320
rect 14924 30311 14976 30320
rect 14924 30277 14933 30311
rect 14933 30277 14967 30311
rect 14967 30277 14976 30311
rect 14924 30268 14976 30277
rect 15292 30268 15344 30320
rect 17040 30311 17092 30320
rect 17040 30277 17049 30311
rect 17049 30277 17083 30311
rect 17083 30277 17092 30311
rect 17040 30268 17092 30277
rect 2044 30200 2096 30252
rect 3792 30200 3844 30252
rect 4068 30200 4120 30252
rect 20352 30268 20404 30320
rect 3424 30175 3476 30184
rect 3424 30141 3433 30175
rect 3433 30141 3467 30175
rect 3467 30141 3476 30175
rect 3424 30132 3476 30141
rect 3976 30132 4028 30184
rect 5908 30132 5960 30184
rect 7748 30132 7800 30184
rect 8024 30132 8076 30184
rect 10784 30132 10836 30184
rect 10876 30175 10928 30184
rect 10876 30141 10885 30175
rect 10885 30141 10919 30175
rect 10919 30141 10928 30175
rect 10876 30132 10928 30141
rect 11704 30175 11756 30184
rect 1676 30107 1728 30116
rect 1676 30073 1685 30107
rect 1685 30073 1719 30107
rect 1719 30073 1728 30107
rect 1676 30064 1728 30073
rect 3608 29996 3660 30048
rect 3792 29996 3844 30048
rect 7472 29996 7524 30048
rect 7932 29996 7984 30048
rect 10692 29996 10744 30048
rect 10876 29996 10928 30048
rect 11704 30141 11713 30175
rect 11713 30141 11747 30175
rect 11747 30141 11756 30175
rect 11704 30132 11756 30141
rect 11520 30064 11572 30116
rect 12532 30132 12584 30184
rect 13176 30175 13228 30184
rect 13176 30141 13185 30175
rect 13185 30141 13219 30175
rect 13219 30141 13228 30175
rect 13176 30132 13228 30141
rect 12992 29996 13044 30048
rect 14096 30132 14148 30184
rect 14832 30064 14884 30116
rect 16120 30132 16172 30184
rect 16580 30132 16632 30184
rect 16948 30175 17000 30184
rect 16948 30141 16957 30175
rect 16957 30141 16991 30175
rect 16991 30141 17000 30175
rect 16948 30132 17000 30141
rect 17408 30175 17460 30184
rect 17408 30141 17417 30175
rect 17417 30141 17451 30175
rect 17451 30141 17460 30175
rect 17408 30132 17460 30141
rect 16488 30064 16540 30116
rect 18880 30200 18932 30252
rect 19616 30243 19668 30252
rect 19616 30209 19625 30243
rect 19625 30209 19659 30243
rect 19659 30209 19668 30243
rect 19616 30200 19668 30209
rect 20720 30200 20772 30252
rect 17868 30132 17920 30184
rect 19432 30132 19484 30184
rect 29184 30132 29236 30184
rect 37280 30200 37332 30252
rect 37648 30132 37700 30184
rect 14740 29996 14792 30048
rect 20352 30064 20404 30116
rect 18236 29996 18288 30048
rect 18696 29996 18748 30048
rect 18972 29996 19024 30048
rect 20260 29996 20312 30048
rect 29460 30039 29512 30048
rect 29460 30005 29469 30039
rect 29469 30005 29503 30039
rect 29503 30005 29512 30039
rect 29460 29996 29512 30005
rect 38200 30039 38252 30048
rect 38200 30005 38209 30039
rect 38209 30005 38243 30039
rect 38243 30005 38252 30039
rect 38200 29996 38252 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 3884 29792 3936 29844
rect 4804 29792 4856 29844
rect 7748 29792 7800 29844
rect 8024 29792 8076 29844
rect 8392 29792 8444 29844
rect 9588 29792 9640 29844
rect 3424 29656 3476 29708
rect 3884 29656 3936 29708
rect 3608 29588 3660 29640
rect 5816 29656 5868 29708
rect 9680 29724 9732 29776
rect 9956 29792 10008 29844
rect 10416 29724 10468 29776
rect 5908 29588 5960 29640
rect 3976 29520 4028 29572
rect 4712 29520 4764 29572
rect 6368 29520 6420 29572
rect 7104 29588 7156 29640
rect 5540 29452 5592 29504
rect 8116 29520 8168 29572
rect 6920 29452 6972 29504
rect 9404 29520 9456 29572
rect 11520 29656 11572 29708
rect 12532 29792 12584 29844
rect 16488 29792 16540 29844
rect 16580 29792 16632 29844
rect 12900 29724 12952 29776
rect 14464 29724 14516 29776
rect 15936 29724 15988 29776
rect 19432 29724 19484 29776
rect 19616 29792 19668 29844
rect 20812 29835 20864 29844
rect 20812 29801 20821 29835
rect 20821 29801 20855 29835
rect 20855 29801 20864 29835
rect 20812 29792 20864 29801
rect 21548 29792 21600 29844
rect 22560 29835 22612 29844
rect 22560 29801 22569 29835
rect 22569 29801 22603 29835
rect 22603 29801 22612 29835
rect 22560 29792 22612 29801
rect 38016 29835 38068 29844
rect 38016 29801 38025 29835
rect 38025 29801 38059 29835
rect 38059 29801 38068 29835
rect 38016 29792 38068 29801
rect 29460 29724 29512 29776
rect 15568 29699 15620 29708
rect 15568 29665 15577 29699
rect 15577 29665 15611 29699
rect 15611 29665 15620 29699
rect 15568 29656 15620 29665
rect 17316 29588 17368 29640
rect 10876 29520 10928 29572
rect 11520 29520 11572 29572
rect 12256 29452 12308 29504
rect 12440 29452 12492 29504
rect 12808 29452 12860 29504
rect 13084 29563 13136 29572
rect 13084 29529 13093 29563
rect 13093 29529 13127 29563
rect 13127 29529 13136 29563
rect 13084 29520 13136 29529
rect 13360 29520 13412 29572
rect 14556 29520 14608 29572
rect 14740 29520 14792 29572
rect 14924 29520 14976 29572
rect 19340 29588 19392 29640
rect 19432 29631 19484 29640
rect 19432 29597 19441 29631
rect 19441 29597 19475 29631
rect 19475 29597 19484 29631
rect 21548 29656 21600 29708
rect 19432 29588 19484 29597
rect 20720 29631 20772 29640
rect 20720 29597 20729 29631
rect 20729 29597 20763 29631
rect 20763 29597 20772 29631
rect 20720 29588 20772 29597
rect 18144 29563 18196 29572
rect 18144 29529 18153 29563
rect 18153 29529 18187 29563
rect 18187 29529 18196 29563
rect 18144 29520 18196 29529
rect 18236 29563 18288 29572
rect 18236 29529 18245 29563
rect 18245 29529 18279 29563
rect 18279 29529 18288 29563
rect 18236 29520 18288 29529
rect 18420 29520 18472 29572
rect 18788 29563 18840 29572
rect 18788 29529 18797 29563
rect 18797 29529 18831 29563
rect 18831 29529 18840 29563
rect 18788 29520 18840 29529
rect 18880 29520 18932 29572
rect 27344 29656 27396 29708
rect 15476 29452 15528 29504
rect 17500 29452 17552 29504
rect 37648 29452 37700 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 1676 29223 1728 29232
rect 1676 29189 1685 29223
rect 1685 29189 1719 29223
rect 1719 29189 1728 29223
rect 1676 29180 1728 29189
rect 3056 29180 3108 29232
rect 9496 29248 9548 29300
rect 7932 29180 7984 29232
rect 8208 29223 8260 29232
rect 8208 29189 8217 29223
rect 8217 29189 8251 29223
rect 8251 29189 8260 29223
rect 8208 29180 8260 29189
rect 8392 29180 8444 29232
rect 9312 29180 9364 29232
rect 1768 29112 1820 29164
rect 5540 29112 5592 29164
rect 3148 29044 3200 29096
rect 848 28976 900 29028
rect 5908 29044 5960 29096
rect 6092 29112 6144 29164
rect 6276 29044 6328 29096
rect 6920 29087 6972 29096
rect 6920 29053 6929 29087
rect 6929 29053 6963 29087
rect 6963 29053 6972 29087
rect 6920 29044 6972 29053
rect 9404 29044 9456 29096
rect 13360 29248 13412 29300
rect 10140 29180 10192 29232
rect 10876 29180 10928 29232
rect 11980 29223 12032 29232
rect 11152 29155 11204 29164
rect 11152 29121 11161 29155
rect 11161 29121 11195 29155
rect 11195 29121 11204 29155
rect 11980 29189 11989 29223
rect 11989 29189 12023 29223
rect 12023 29189 12032 29223
rect 11980 29180 12032 29189
rect 13820 29180 13872 29232
rect 11152 29112 11204 29121
rect 10324 29044 10376 29096
rect 16948 29248 17000 29300
rect 14188 29223 14240 29232
rect 14188 29189 14197 29223
rect 14197 29189 14231 29223
rect 14231 29189 14240 29223
rect 14188 29180 14240 29189
rect 15384 29223 15436 29232
rect 15384 29189 15393 29223
rect 15393 29189 15427 29223
rect 15427 29189 15436 29223
rect 15384 29180 15436 29189
rect 16120 29180 16172 29232
rect 16212 29180 16264 29232
rect 18880 29248 18932 29300
rect 22928 29248 22980 29300
rect 17500 29223 17552 29232
rect 17500 29189 17509 29223
rect 17509 29189 17543 29223
rect 17543 29189 17552 29223
rect 17500 29180 17552 29189
rect 17592 29223 17644 29232
rect 17592 29189 17601 29223
rect 17601 29189 17635 29223
rect 17635 29189 17644 29223
rect 17592 29180 17644 29189
rect 18972 29180 19024 29232
rect 19432 29155 19484 29164
rect 19432 29121 19441 29155
rect 19441 29121 19475 29155
rect 19475 29121 19484 29155
rect 19432 29112 19484 29121
rect 20260 29155 20312 29164
rect 20260 29121 20269 29155
rect 20269 29121 20303 29155
rect 20303 29121 20312 29155
rect 20260 29112 20312 29121
rect 14096 29087 14148 29096
rect 14096 29053 14106 29087
rect 14106 29053 14140 29087
rect 14140 29053 14148 29087
rect 14096 29044 14148 29053
rect 15292 29087 15344 29096
rect 3424 28908 3476 28960
rect 4068 28908 4120 28960
rect 5080 28908 5132 28960
rect 5632 28908 5684 28960
rect 8208 28976 8260 29028
rect 8668 28976 8720 29028
rect 10232 28976 10284 29028
rect 11244 28976 11296 29028
rect 13176 28976 13228 29028
rect 5816 28908 5868 28960
rect 6276 28908 6328 28960
rect 7656 28908 7708 28960
rect 7748 28908 7800 28960
rect 10140 28908 10192 28960
rect 11980 28908 12032 28960
rect 13360 28908 13412 28960
rect 14648 29019 14700 29028
rect 14648 28985 14657 29019
rect 14657 28985 14691 29019
rect 14691 28985 14700 29019
rect 14648 28976 14700 28985
rect 15292 29053 15301 29087
rect 15301 29053 15335 29087
rect 15335 29053 15344 29087
rect 15292 29044 15344 29053
rect 17316 29087 17368 29096
rect 17316 29053 17325 29087
rect 17325 29053 17359 29087
rect 17359 29053 17368 29087
rect 17316 29044 17368 29053
rect 17868 29044 17920 29096
rect 18236 29087 18288 29096
rect 18236 29053 18245 29087
rect 18245 29053 18279 29087
rect 18279 29053 18288 29087
rect 18236 29044 18288 29053
rect 18512 29087 18564 29096
rect 18512 29053 18521 29087
rect 18521 29053 18555 29087
rect 18555 29053 18564 29087
rect 18512 29044 18564 29053
rect 20720 29044 20772 29096
rect 20904 29155 20956 29164
rect 20904 29121 20913 29155
rect 20913 29121 20947 29155
rect 20947 29121 20956 29155
rect 37372 29180 37424 29232
rect 20904 29112 20956 29121
rect 34520 29112 34572 29164
rect 18972 28976 19024 29028
rect 38200 29019 38252 29028
rect 38200 28985 38209 29019
rect 38209 28985 38243 29019
rect 38243 28985 38252 29019
rect 38200 28976 38252 28985
rect 16212 28908 16264 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 6920 28704 6972 28756
rect 7564 28704 7616 28756
rect 11888 28704 11940 28756
rect 13360 28704 13412 28756
rect 16028 28704 16080 28756
rect 9864 28636 9916 28688
rect 10968 28636 11020 28688
rect 11704 28636 11756 28688
rect 11980 28636 12032 28688
rect 13544 28636 13596 28688
rect 2596 28543 2648 28552
rect 1860 28432 1912 28484
rect 2596 28509 2605 28543
rect 2605 28509 2639 28543
rect 2639 28509 2648 28543
rect 2596 28500 2648 28509
rect 3424 28543 3476 28552
rect 3424 28509 3433 28543
rect 3433 28509 3467 28543
rect 3467 28509 3476 28543
rect 3424 28500 3476 28509
rect 2872 28432 2924 28484
rect 4160 28568 4212 28620
rect 6184 28568 6236 28620
rect 7748 28568 7800 28620
rect 7564 28500 7616 28552
rect 10140 28568 10192 28620
rect 11244 28568 11296 28620
rect 10600 28500 10652 28552
rect 12624 28568 12676 28620
rect 15568 28636 15620 28688
rect 15936 28636 15988 28688
rect 14832 28568 14884 28620
rect 16120 28568 16172 28620
rect 16856 28704 16908 28756
rect 17040 28704 17092 28756
rect 17316 28704 17368 28756
rect 22836 28704 22888 28756
rect 33968 28747 34020 28756
rect 33968 28713 33977 28747
rect 33977 28713 34011 28747
rect 34011 28713 34020 28747
rect 33968 28704 34020 28713
rect 16672 28636 16724 28688
rect 34520 28636 34572 28688
rect 16948 28611 17000 28620
rect 16948 28577 16957 28611
rect 16957 28577 16991 28611
rect 16991 28577 17000 28611
rect 16948 28568 17000 28577
rect 18972 28568 19024 28620
rect 19156 28500 19208 28552
rect 30748 28543 30800 28552
rect 30748 28509 30757 28543
rect 30757 28509 30791 28543
rect 30791 28509 30800 28543
rect 30748 28500 30800 28509
rect 34152 28543 34204 28552
rect 34152 28509 34161 28543
rect 34161 28509 34195 28543
rect 34195 28509 34204 28543
rect 34152 28500 34204 28509
rect 4068 28475 4120 28484
rect 4068 28441 4077 28475
rect 4077 28441 4111 28475
rect 4111 28441 4120 28475
rect 4068 28432 4120 28441
rect 5080 28432 5132 28484
rect 4620 28364 4672 28416
rect 6644 28432 6696 28484
rect 5724 28364 5776 28416
rect 6276 28364 6328 28416
rect 7748 28364 7800 28416
rect 7932 28432 7984 28484
rect 8392 28432 8444 28484
rect 9404 28475 9456 28484
rect 9404 28441 9413 28475
rect 9413 28441 9447 28475
rect 9447 28441 9456 28475
rect 9404 28432 9456 28441
rect 9496 28475 9548 28484
rect 9496 28441 9505 28475
rect 9505 28441 9539 28475
rect 9539 28441 9548 28475
rect 11428 28475 11480 28484
rect 9496 28432 9548 28441
rect 11428 28441 11437 28475
rect 11437 28441 11471 28475
rect 11471 28441 11480 28475
rect 11428 28432 11480 28441
rect 11520 28475 11572 28484
rect 11520 28441 11529 28475
rect 11529 28441 11563 28475
rect 11563 28441 11572 28475
rect 11520 28432 11572 28441
rect 11704 28432 11756 28484
rect 12624 28475 12676 28484
rect 12624 28441 12633 28475
rect 12633 28441 12667 28475
rect 12667 28441 12676 28475
rect 12624 28432 12676 28441
rect 13636 28432 13688 28484
rect 16212 28475 16264 28484
rect 10324 28364 10376 28416
rect 11060 28364 11112 28416
rect 16212 28441 16221 28475
rect 16221 28441 16255 28475
rect 16255 28441 16264 28475
rect 16212 28432 16264 28441
rect 16396 28364 16448 28416
rect 18512 28432 18564 28484
rect 18696 28475 18748 28484
rect 18696 28441 18705 28475
rect 18705 28441 18739 28475
rect 18739 28441 18748 28475
rect 18696 28432 18748 28441
rect 19248 28432 19300 28484
rect 18236 28364 18288 28416
rect 18420 28364 18472 28416
rect 19984 28364 20036 28416
rect 20076 28407 20128 28416
rect 20076 28373 20085 28407
rect 20085 28373 20119 28407
rect 20119 28373 20128 28407
rect 20076 28364 20128 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 4068 28160 4120 28212
rect 4988 28092 5040 28144
rect 5540 28092 5592 28144
rect 9588 28160 9640 28212
rect 11980 28160 12032 28212
rect 16396 28160 16448 28212
rect 18144 28160 18196 28212
rect 9680 28092 9732 28144
rect 10692 28092 10744 28144
rect 2320 28024 2372 28076
rect 3332 28067 3384 28076
rect 3332 28033 3341 28067
rect 3341 28033 3375 28067
rect 3375 28033 3384 28067
rect 3332 28024 3384 28033
rect 4068 28024 4120 28076
rect 4528 28067 4580 28076
rect 4528 28033 4537 28067
rect 4537 28033 4571 28067
rect 4571 28033 4580 28067
rect 4528 28024 4580 28033
rect 5448 28024 5500 28076
rect 3148 27956 3200 28008
rect 5724 27956 5776 28008
rect 6644 28024 6696 28076
rect 6920 28067 6972 28076
rect 6920 28033 6929 28067
rect 6929 28033 6963 28067
rect 6963 28033 6972 28067
rect 6920 28024 6972 28033
rect 7472 28024 7524 28076
rect 9956 28067 10008 28076
rect 9956 28033 9965 28067
rect 9965 28033 9999 28067
rect 9999 28033 10008 28067
rect 12256 28067 12308 28076
rect 9956 28024 10008 28033
rect 12256 28033 12265 28067
rect 12265 28033 12299 28067
rect 12299 28033 12308 28067
rect 12256 28024 12308 28033
rect 6184 27956 6236 28008
rect 7656 27999 7708 28008
rect 7656 27965 7665 27999
rect 7665 27965 7699 27999
rect 7699 27965 7708 27999
rect 7656 27956 7708 27965
rect 8392 27956 8444 28008
rect 9036 27956 9088 28008
rect 10324 27956 10376 28008
rect 12900 27956 12952 28008
rect 1676 27931 1728 27940
rect 1676 27897 1685 27931
rect 1685 27897 1719 27931
rect 1719 27897 1728 27931
rect 1676 27888 1728 27897
rect 7564 27888 7616 27940
rect 5908 27820 5960 27872
rect 6552 27820 6604 27872
rect 10784 27888 10836 27940
rect 11060 27931 11112 27940
rect 11060 27897 11069 27931
rect 11069 27897 11103 27931
rect 11103 27897 11112 27931
rect 13636 28092 13688 28144
rect 14280 28135 14332 28144
rect 14280 28101 14289 28135
rect 14289 28101 14323 28135
rect 14323 28101 14332 28135
rect 14280 28092 14332 28101
rect 14464 28092 14516 28144
rect 16028 28024 16080 28076
rect 16580 28092 16632 28144
rect 16488 28024 16540 28076
rect 23572 28160 23624 28212
rect 18604 28092 18656 28144
rect 22652 28092 22704 28144
rect 19984 28067 20036 28076
rect 19984 28033 19993 28067
rect 19993 28033 20027 28067
rect 20027 28033 20036 28067
rect 19984 28024 20036 28033
rect 14648 27999 14700 28008
rect 14648 27965 14657 27999
rect 14657 27965 14691 27999
rect 14691 27965 14700 27999
rect 14648 27956 14700 27965
rect 15016 27956 15068 28008
rect 16948 27999 17000 28008
rect 11060 27888 11112 27897
rect 15568 27888 15620 27940
rect 14372 27820 14424 27872
rect 15200 27820 15252 27872
rect 16948 27965 16957 27999
rect 16957 27965 16991 27999
rect 16991 27965 17000 27999
rect 16948 27956 17000 27965
rect 16856 27888 16908 27940
rect 18696 27956 18748 28008
rect 18880 27999 18932 28008
rect 18880 27965 18889 27999
rect 18889 27965 18923 27999
rect 18923 27965 18932 27999
rect 18880 27956 18932 27965
rect 19340 27956 19392 28008
rect 18512 27888 18564 27940
rect 26240 27888 26292 27940
rect 19156 27820 19208 27872
rect 19248 27820 19300 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 2872 27616 2924 27668
rect 8116 27616 8168 27668
rect 10692 27616 10744 27668
rect 11520 27616 11572 27668
rect 16856 27616 16908 27668
rect 18880 27659 18932 27668
rect 18880 27625 18889 27659
rect 18889 27625 18923 27659
rect 18923 27625 18932 27659
rect 18880 27616 18932 27625
rect 22652 27616 22704 27668
rect 22836 27659 22888 27668
rect 22836 27625 22845 27659
rect 22845 27625 22879 27659
rect 22879 27625 22888 27659
rect 22836 27616 22888 27625
rect 2044 27548 2096 27600
rect 4620 27548 4672 27600
rect 2872 27480 2924 27532
rect 10324 27548 10376 27600
rect 14648 27591 14700 27600
rect 14648 27557 14657 27591
rect 14657 27557 14691 27591
rect 14691 27557 14700 27591
rect 14648 27548 14700 27557
rect 3700 27412 3752 27464
rect 5540 27412 5592 27464
rect 6460 27455 6512 27464
rect 3608 27276 3660 27328
rect 3884 27276 3936 27328
rect 6092 27344 6144 27396
rect 6460 27421 6469 27455
rect 6469 27421 6503 27455
rect 6503 27421 6512 27455
rect 6460 27412 6512 27421
rect 7104 27455 7156 27464
rect 7104 27421 7113 27455
rect 7113 27421 7147 27455
rect 7147 27421 7156 27455
rect 7104 27412 7156 27421
rect 7380 27412 7432 27464
rect 8760 27412 8812 27464
rect 9036 27412 9088 27464
rect 9312 27455 9364 27464
rect 9312 27421 9321 27455
rect 9321 27421 9355 27455
rect 9355 27421 9364 27455
rect 9312 27412 9364 27421
rect 9404 27412 9456 27464
rect 6920 27344 6972 27396
rect 4896 27276 4948 27328
rect 6460 27276 6512 27328
rect 7564 27276 7616 27328
rect 8300 27276 8352 27328
rect 9680 27276 9732 27328
rect 9772 27319 9824 27328
rect 9772 27285 9781 27319
rect 9781 27285 9815 27319
rect 9815 27285 9824 27319
rect 10140 27344 10192 27396
rect 11244 27387 11296 27396
rect 11244 27353 11253 27387
rect 11253 27353 11287 27387
rect 11287 27353 11296 27387
rect 12440 27480 12492 27532
rect 12900 27480 12952 27532
rect 15844 27523 15896 27532
rect 15844 27489 15853 27523
rect 15853 27489 15887 27523
rect 15887 27489 15896 27523
rect 15844 27480 15896 27489
rect 16488 27480 16540 27532
rect 14556 27412 14608 27464
rect 20076 27480 20128 27532
rect 20444 27523 20496 27532
rect 20444 27489 20453 27523
rect 20453 27489 20487 27523
rect 20487 27489 20496 27523
rect 20444 27480 20496 27489
rect 18236 27455 18288 27464
rect 11244 27344 11296 27353
rect 13084 27387 13136 27396
rect 13084 27353 13093 27387
rect 13093 27353 13127 27387
rect 13127 27353 13136 27387
rect 15108 27387 15160 27396
rect 13084 27344 13136 27353
rect 9772 27276 9824 27285
rect 11888 27276 11940 27328
rect 12992 27276 13044 27328
rect 15108 27353 15117 27387
rect 15117 27353 15151 27387
rect 15151 27353 15160 27387
rect 15108 27344 15160 27353
rect 16672 27344 16724 27396
rect 16856 27387 16908 27396
rect 16856 27353 16865 27387
rect 16865 27353 16899 27387
rect 16899 27353 16908 27387
rect 16856 27344 16908 27353
rect 18236 27421 18245 27455
rect 18245 27421 18279 27455
rect 18279 27421 18288 27455
rect 18236 27412 18288 27421
rect 17684 27344 17736 27396
rect 20352 27344 20404 27396
rect 16948 27276 17000 27328
rect 21180 27319 21232 27328
rect 21180 27285 21189 27319
rect 21189 27285 21223 27319
rect 21223 27285 21232 27319
rect 21180 27276 21232 27285
rect 34152 27344 34204 27396
rect 34796 27344 34848 27396
rect 37924 27276 37976 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 2504 27072 2556 27124
rect 3056 27115 3108 27124
rect 3056 27081 3065 27115
rect 3065 27081 3099 27115
rect 3099 27081 3108 27115
rect 3056 27072 3108 27081
rect 3884 27072 3936 27124
rect 4896 27004 4948 27056
rect 1768 26936 1820 26988
rect 2504 26979 2556 26988
rect 2504 26945 2513 26979
rect 2513 26945 2547 26979
rect 2547 26945 2556 26979
rect 2504 26936 2556 26945
rect 2964 26979 3016 26988
rect 2320 26868 2372 26920
rect 2964 26945 2973 26979
rect 2973 26945 3007 26979
rect 3007 26945 3016 26979
rect 2964 26936 3016 26945
rect 3240 26936 3292 26988
rect 5080 26936 5132 26988
rect 5448 27072 5500 27124
rect 5824 26985 5876 26994
rect 5824 26951 5833 26985
rect 5833 26951 5867 26985
rect 5867 26951 5876 26985
rect 6184 27072 6236 27124
rect 8208 27072 8260 27124
rect 9312 27072 9364 27124
rect 11060 27072 11112 27124
rect 11244 27072 11296 27124
rect 16120 27072 16172 27124
rect 16580 27072 16632 27124
rect 18236 27072 18288 27124
rect 20352 27115 20404 27124
rect 7840 27004 7892 27056
rect 9128 27004 9180 27056
rect 9220 27047 9272 27056
rect 9220 27013 9229 27047
rect 9229 27013 9263 27047
rect 9263 27013 9272 27047
rect 9220 27004 9272 27013
rect 5824 26942 5876 26951
rect 7380 26936 7432 26988
rect 8024 26868 8076 26920
rect 9128 26911 9180 26920
rect 9128 26877 9137 26911
rect 9137 26877 9171 26911
rect 9171 26877 9180 26911
rect 9128 26868 9180 26877
rect 9036 26800 9088 26852
rect 9680 26843 9732 26852
rect 9680 26809 9689 26843
rect 9689 26809 9723 26843
rect 9723 26809 9732 26843
rect 9680 26800 9732 26809
rect 1676 26775 1728 26784
rect 1676 26741 1685 26775
rect 1685 26741 1719 26775
rect 1719 26741 1728 26775
rect 1676 26732 1728 26741
rect 3056 26732 3108 26784
rect 4896 26732 4948 26784
rect 6184 26732 6236 26784
rect 10600 27004 10652 27056
rect 10968 27047 11020 27056
rect 10968 27013 10977 27047
rect 10977 27013 11011 27047
rect 11011 27013 11020 27047
rect 10968 27004 11020 27013
rect 11888 27047 11940 27056
rect 11888 27013 11897 27047
rect 11897 27013 11931 27047
rect 11931 27013 11940 27047
rect 11888 27004 11940 27013
rect 13084 27004 13136 27056
rect 14372 27047 14424 27056
rect 14372 27013 14381 27047
rect 14381 27013 14415 27047
rect 14415 27013 14424 27047
rect 14372 27004 14424 27013
rect 14924 27047 14976 27056
rect 14924 27013 14933 27047
rect 14933 27013 14967 27047
rect 14967 27013 14976 27047
rect 14924 27004 14976 27013
rect 15108 27004 15160 27056
rect 17960 27004 18012 27056
rect 19340 27004 19392 27056
rect 19524 27004 19576 27056
rect 20352 27081 20361 27115
rect 20361 27081 20395 27115
rect 20395 27081 20404 27115
rect 20352 27072 20404 27081
rect 13452 26936 13504 26988
rect 16120 26979 16172 26988
rect 10324 26911 10376 26920
rect 10324 26877 10333 26911
rect 10333 26877 10367 26911
rect 10367 26877 10376 26911
rect 10324 26868 10376 26877
rect 9864 26800 9916 26852
rect 12256 26868 12308 26920
rect 14096 26868 14148 26920
rect 16120 26945 16129 26979
rect 16129 26945 16163 26979
rect 16163 26945 16172 26979
rect 16120 26936 16172 26945
rect 17684 26936 17736 26988
rect 18604 26936 18656 26988
rect 17224 26868 17276 26920
rect 17868 26800 17920 26852
rect 19340 26868 19392 26920
rect 21180 27004 21232 27056
rect 20720 26936 20772 26988
rect 21640 26936 21692 26988
rect 18604 26800 18656 26852
rect 22652 27072 22704 27124
rect 25320 27072 25372 27124
rect 22284 27004 22336 27056
rect 37740 27004 37792 27056
rect 23572 26979 23624 26988
rect 23572 26945 23581 26979
rect 23581 26945 23615 26979
rect 23615 26945 23624 26979
rect 23572 26936 23624 26945
rect 38200 26979 38252 26988
rect 38200 26945 38209 26979
rect 38209 26945 38243 26979
rect 38243 26945 38252 26979
rect 38200 26936 38252 26945
rect 38292 26800 38344 26852
rect 10324 26732 10376 26784
rect 12808 26732 12860 26784
rect 13636 26775 13688 26784
rect 13636 26741 13645 26775
rect 13645 26741 13679 26775
rect 13679 26741 13688 26775
rect 13636 26732 13688 26741
rect 15384 26732 15436 26784
rect 16120 26732 16172 26784
rect 22284 26732 22336 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 2136 26528 2188 26580
rect 2412 26528 2464 26580
rect 1308 26460 1360 26512
rect 848 26392 900 26444
rect 3056 26392 3108 26444
rect 3148 26392 3200 26444
rect 3884 26392 3936 26444
rect 2320 26324 2372 26376
rect 1952 26256 2004 26308
rect 2136 26256 2188 26308
rect 2412 26188 2464 26240
rect 2780 26324 2832 26376
rect 3608 26324 3660 26376
rect 4528 26324 4580 26376
rect 5080 26528 5132 26580
rect 7012 26528 7064 26580
rect 7380 26528 7432 26580
rect 7564 26528 7616 26580
rect 7656 26528 7708 26580
rect 9772 26528 9824 26580
rect 10048 26528 10100 26580
rect 11888 26528 11940 26580
rect 12440 26528 12492 26580
rect 13728 26528 13780 26580
rect 15108 26571 15160 26580
rect 15108 26537 15117 26571
rect 15117 26537 15151 26571
rect 15151 26537 15160 26571
rect 15108 26528 15160 26537
rect 17132 26571 17184 26580
rect 17132 26537 17141 26571
rect 17141 26537 17175 26571
rect 17175 26537 17184 26571
rect 17132 26528 17184 26537
rect 17224 26528 17276 26580
rect 18696 26528 18748 26580
rect 18880 26571 18932 26580
rect 18880 26537 18889 26571
rect 18889 26537 18923 26571
rect 18923 26537 18932 26571
rect 18880 26528 18932 26537
rect 19616 26528 19668 26580
rect 20536 26528 20588 26580
rect 20720 26528 20772 26580
rect 4896 26324 4948 26376
rect 5632 26324 5684 26376
rect 6644 26367 6696 26376
rect 6644 26333 6653 26367
rect 6653 26333 6687 26367
rect 6687 26333 6696 26367
rect 6644 26324 6696 26333
rect 4804 26256 4856 26308
rect 3148 26188 3200 26240
rect 5080 26188 5132 26240
rect 6460 26256 6512 26308
rect 7012 26324 7064 26376
rect 7288 26324 7340 26376
rect 9036 26392 9088 26444
rect 9404 26324 9456 26376
rect 9956 26367 10008 26376
rect 9956 26333 9965 26367
rect 9965 26333 9999 26367
rect 9999 26333 10008 26367
rect 9956 26324 10008 26333
rect 10324 26392 10376 26444
rect 10784 26435 10836 26444
rect 10784 26401 10793 26435
rect 10793 26401 10827 26435
rect 10827 26401 10836 26435
rect 10784 26392 10836 26401
rect 13084 26460 13136 26512
rect 11520 26324 11572 26376
rect 11888 26367 11940 26376
rect 11888 26333 11897 26367
rect 11897 26333 11931 26367
rect 11931 26333 11940 26367
rect 11888 26324 11940 26333
rect 7656 26256 7708 26308
rect 7932 26299 7984 26308
rect 7932 26265 7941 26299
rect 7941 26265 7975 26299
rect 7975 26265 7984 26299
rect 7932 26256 7984 26265
rect 8024 26299 8076 26308
rect 8024 26265 8033 26299
rect 8033 26265 8067 26299
rect 8067 26265 8076 26299
rect 8024 26256 8076 26265
rect 8300 26256 8352 26308
rect 8760 26256 8812 26308
rect 9312 26256 9364 26308
rect 9680 26256 9732 26308
rect 9220 26188 9272 26240
rect 9496 26188 9548 26240
rect 12716 26188 12768 26240
rect 14924 26392 14976 26444
rect 15384 26392 15436 26444
rect 16396 26460 16448 26512
rect 12900 26324 12952 26376
rect 18144 26392 18196 26444
rect 18328 26392 18380 26444
rect 16948 26367 17000 26376
rect 14556 26256 14608 26308
rect 13912 26188 13964 26240
rect 14648 26188 14700 26240
rect 15476 26188 15528 26240
rect 16948 26333 16957 26367
rect 16957 26333 16991 26367
rect 16991 26333 17000 26367
rect 16948 26324 17000 26333
rect 17500 26324 17552 26376
rect 18420 26367 18472 26376
rect 18420 26333 18429 26367
rect 18429 26333 18463 26367
rect 18463 26333 18472 26367
rect 18420 26324 18472 26333
rect 17960 26256 18012 26308
rect 16304 26188 16356 26240
rect 20628 26324 20680 26376
rect 18696 26256 18748 26308
rect 37740 26256 37792 26308
rect 18604 26188 18656 26240
rect 38384 26188 38436 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 2044 25984 2096 26036
rect 4068 26027 4120 26036
rect 4068 25993 4077 26027
rect 4077 25993 4111 26027
rect 4111 25993 4120 26027
rect 4068 25984 4120 25993
rect 4988 25984 5040 26036
rect 13728 26027 13780 26036
rect 4712 25916 4764 25968
rect 6184 25916 6236 25968
rect 9036 25959 9088 25968
rect 9036 25925 9045 25959
rect 9045 25925 9079 25959
rect 9079 25925 9088 25959
rect 9036 25916 9088 25925
rect 9312 25916 9364 25968
rect 9772 25916 9824 25968
rect 13728 25993 13737 26027
rect 13737 25993 13771 26027
rect 13771 25993 13780 26027
rect 13728 25984 13780 25993
rect 13912 25984 13964 26036
rect 13084 25959 13136 25968
rect 13084 25925 13093 25959
rect 13093 25925 13127 25959
rect 13127 25925 13136 25959
rect 13084 25916 13136 25925
rect 14096 25916 14148 25968
rect 18328 25984 18380 26036
rect 18420 25984 18472 26036
rect 20536 25984 20588 26036
rect 37832 26027 37884 26036
rect 37832 25993 37841 26027
rect 37841 25993 37875 26027
rect 37875 25993 37884 26027
rect 37832 25984 37884 25993
rect 19432 25916 19484 25968
rect 20720 25916 20772 25968
rect 2780 25848 2832 25900
rect 3148 25891 3200 25900
rect 3148 25857 3157 25891
rect 3157 25857 3191 25891
rect 3191 25857 3200 25891
rect 3148 25848 3200 25857
rect 2964 25780 3016 25832
rect 4068 25848 4120 25900
rect 4620 25848 4672 25900
rect 5080 25848 5132 25900
rect 3792 25780 3844 25832
rect 5724 25848 5776 25900
rect 6736 25848 6788 25900
rect 10968 25891 11020 25900
rect 10968 25857 10977 25891
rect 10977 25857 11011 25891
rect 11011 25857 11020 25891
rect 10968 25848 11020 25857
rect 11796 25848 11848 25900
rect 13636 25848 13688 25900
rect 14832 25848 14884 25900
rect 15660 25891 15712 25900
rect 15660 25857 15669 25891
rect 15669 25857 15703 25891
rect 15703 25857 15712 25891
rect 15660 25848 15712 25857
rect 16304 25891 16356 25900
rect 16304 25857 16313 25891
rect 16313 25857 16347 25891
rect 16347 25857 16356 25891
rect 16304 25848 16356 25857
rect 17500 25848 17552 25900
rect 17960 25891 18012 25900
rect 17960 25857 17969 25891
rect 17969 25857 18003 25891
rect 18003 25857 18012 25891
rect 17960 25848 18012 25857
rect 5632 25780 5684 25832
rect 7564 25780 7616 25832
rect 8300 25780 8352 25832
rect 9772 25823 9824 25832
rect 5172 25712 5224 25764
rect 2412 25644 2464 25696
rect 3148 25644 3200 25696
rect 6276 25644 6328 25696
rect 8668 25712 8720 25764
rect 8208 25644 8260 25696
rect 9772 25789 9781 25823
rect 9781 25789 9815 25823
rect 9815 25789 9824 25823
rect 9772 25780 9824 25789
rect 9220 25712 9272 25764
rect 10600 25712 10652 25764
rect 12440 25712 12492 25764
rect 12900 25712 12952 25764
rect 13544 25780 13596 25832
rect 13912 25780 13964 25832
rect 14188 25823 14240 25832
rect 14188 25789 14197 25823
rect 14197 25789 14231 25823
rect 14231 25789 14240 25823
rect 14188 25780 14240 25789
rect 18236 25780 18288 25832
rect 14464 25712 14516 25764
rect 17040 25712 17092 25764
rect 20996 25848 21048 25900
rect 19892 25823 19944 25832
rect 19892 25789 19901 25823
rect 19901 25789 19935 25823
rect 19935 25789 19944 25823
rect 19892 25780 19944 25789
rect 21088 25780 21140 25832
rect 19248 25712 19300 25764
rect 38384 25848 38436 25900
rect 11888 25644 11940 25696
rect 12532 25644 12584 25696
rect 13176 25644 13228 25696
rect 13728 25644 13780 25696
rect 13820 25644 13872 25696
rect 15568 25687 15620 25696
rect 15568 25653 15577 25687
rect 15577 25653 15611 25687
rect 15611 25653 15620 25687
rect 15568 25644 15620 25653
rect 15660 25644 15712 25696
rect 20996 25644 21048 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 1216 25440 1268 25492
rect 3516 25440 3568 25492
rect 3976 25440 4028 25492
rect 5264 25440 5316 25492
rect 6184 25483 6236 25492
rect 6184 25449 6193 25483
rect 6193 25449 6227 25483
rect 6227 25449 6236 25483
rect 6184 25440 6236 25449
rect 7932 25483 7984 25492
rect 7932 25449 7941 25483
rect 7941 25449 7975 25483
rect 7975 25449 7984 25483
rect 7932 25440 7984 25449
rect 8024 25440 8076 25492
rect 9036 25372 9088 25424
rect 9312 25372 9364 25424
rect 11704 25372 11756 25424
rect 12624 25440 12676 25492
rect 13544 25372 13596 25424
rect 13636 25372 13688 25424
rect 14924 25415 14976 25424
rect 2964 25304 3016 25356
rect 3700 25304 3752 25356
rect 5632 25347 5684 25356
rect 2504 25279 2556 25288
rect 2504 25245 2513 25279
rect 2513 25245 2547 25279
rect 2547 25245 2556 25279
rect 2504 25236 2556 25245
rect 2780 25236 2832 25288
rect 4160 25279 4212 25288
rect 4160 25245 4169 25279
rect 4169 25245 4203 25279
rect 4203 25245 4212 25279
rect 4804 25279 4856 25288
rect 4160 25236 4212 25245
rect 4804 25245 4813 25279
rect 4813 25245 4847 25279
rect 4847 25245 4856 25279
rect 4804 25236 4856 25245
rect 5632 25313 5641 25347
rect 5641 25313 5675 25347
rect 5675 25313 5684 25347
rect 5632 25304 5684 25313
rect 6000 25304 6052 25356
rect 9496 25304 9548 25356
rect 9864 25304 9916 25356
rect 11428 25304 11480 25356
rect 12440 25347 12492 25356
rect 12440 25313 12449 25347
rect 12449 25313 12483 25347
rect 12483 25313 12492 25347
rect 12440 25304 12492 25313
rect 13084 25304 13136 25356
rect 13820 25304 13872 25356
rect 14924 25381 14933 25415
rect 14933 25381 14967 25415
rect 14967 25381 14976 25415
rect 14924 25372 14976 25381
rect 4988 25168 5040 25220
rect 5172 25168 5224 25220
rect 6368 25168 6420 25220
rect 5632 25100 5684 25152
rect 7288 25236 7340 25288
rect 9128 25168 9180 25220
rect 9772 25211 9824 25220
rect 9772 25177 9781 25211
rect 9781 25177 9815 25211
rect 9815 25177 9824 25211
rect 13636 25236 13688 25288
rect 9772 25168 9824 25177
rect 8024 25100 8076 25152
rect 8300 25100 8352 25152
rect 8484 25100 8536 25152
rect 8576 25100 8628 25152
rect 11704 25168 11756 25220
rect 10232 25100 10284 25152
rect 11428 25100 11480 25152
rect 14372 25168 14424 25220
rect 14464 25211 14516 25220
rect 14464 25177 14473 25211
rect 14473 25177 14507 25211
rect 14507 25177 14516 25211
rect 17776 25440 17828 25492
rect 21088 25483 21140 25492
rect 21088 25449 21097 25483
rect 21097 25449 21131 25483
rect 21131 25449 21140 25483
rect 21088 25440 21140 25449
rect 20444 25415 20496 25424
rect 20444 25381 20453 25415
rect 20453 25381 20487 25415
rect 20487 25381 20496 25415
rect 20444 25372 20496 25381
rect 17500 25304 17552 25356
rect 18236 25347 18288 25356
rect 18236 25313 18245 25347
rect 18245 25313 18279 25347
rect 18279 25313 18288 25347
rect 18236 25304 18288 25313
rect 26240 25304 26292 25356
rect 16396 25279 16448 25288
rect 16396 25245 16405 25279
rect 16405 25245 16439 25279
rect 16439 25245 16448 25279
rect 16396 25236 16448 25245
rect 17040 25279 17092 25288
rect 17040 25245 17049 25279
rect 17049 25245 17083 25279
rect 17083 25245 17092 25279
rect 17040 25236 17092 25245
rect 17684 25279 17736 25288
rect 17684 25245 17693 25279
rect 17693 25245 17727 25279
rect 17727 25245 17736 25279
rect 17684 25236 17736 25245
rect 20996 25236 21048 25288
rect 14464 25168 14516 25177
rect 18328 25211 18380 25220
rect 18328 25177 18337 25211
rect 18337 25177 18371 25211
rect 18371 25177 18380 25211
rect 18328 25168 18380 25177
rect 19432 25168 19484 25220
rect 19892 25211 19944 25220
rect 19892 25177 19901 25211
rect 19901 25177 19935 25211
rect 19935 25177 19944 25211
rect 19892 25168 19944 25177
rect 19984 25211 20036 25220
rect 19984 25177 19993 25211
rect 19993 25177 20027 25211
rect 20027 25177 20036 25211
rect 19984 25168 20036 25177
rect 13820 25100 13872 25152
rect 15844 25100 15896 25152
rect 17868 25100 17920 25152
rect 37740 25236 37792 25288
rect 38108 25236 38160 25288
rect 37280 25168 37332 25220
rect 36820 25100 36872 25152
rect 38016 25143 38068 25152
rect 38016 25109 38025 25143
rect 38025 25109 38059 25143
rect 38059 25109 38068 25143
rect 38016 25100 38068 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 14188 24896 14240 24948
rect 14832 24896 14884 24948
rect 20076 24896 20128 24948
rect 1124 24624 1176 24676
rect 2780 24760 2832 24812
rect 3700 24803 3752 24812
rect 3700 24769 3709 24803
rect 3709 24769 3743 24803
rect 3743 24769 3752 24803
rect 3700 24760 3752 24769
rect 8024 24828 8076 24880
rect 9496 24828 9548 24880
rect 10600 24871 10652 24880
rect 3976 24760 4028 24812
rect 4712 24760 4764 24812
rect 5632 24760 5684 24812
rect 4620 24692 4672 24744
rect 6000 24760 6052 24812
rect 8300 24760 8352 24812
rect 8484 24803 8536 24812
rect 8484 24769 8493 24803
rect 8493 24769 8527 24803
rect 8527 24769 8536 24803
rect 8484 24760 8536 24769
rect 8852 24760 8904 24812
rect 10600 24837 10609 24871
rect 10609 24837 10643 24871
rect 10643 24837 10652 24871
rect 10600 24828 10652 24837
rect 11888 24828 11940 24880
rect 12716 24828 12768 24880
rect 7012 24692 7064 24744
rect 9128 24735 9180 24744
rect 9128 24701 9137 24735
rect 9137 24701 9171 24735
rect 9171 24701 9180 24735
rect 9128 24692 9180 24701
rect 9220 24692 9272 24744
rect 12900 24803 12952 24812
rect 12900 24769 12909 24803
rect 12909 24769 12943 24803
rect 12943 24769 12952 24803
rect 15476 24828 15528 24880
rect 15844 24828 15896 24880
rect 12900 24760 12952 24769
rect 14556 24803 14608 24812
rect 14556 24769 14565 24803
rect 14565 24769 14599 24803
rect 14599 24769 14608 24803
rect 14556 24760 14608 24769
rect 14740 24803 14792 24812
rect 14740 24769 14749 24803
rect 14749 24769 14783 24803
rect 14783 24769 14792 24803
rect 14740 24760 14792 24769
rect 11520 24692 11572 24744
rect 13084 24692 13136 24744
rect 13268 24692 13320 24744
rect 15660 24735 15712 24744
rect 1676 24599 1728 24608
rect 1676 24565 1685 24599
rect 1685 24565 1719 24599
rect 1719 24565 1728 24599
rect 1676 24556 1728 24565
rect 2504 24556 2556 24608
rect 4160 24556 4212 24608
rect 5356 24599 5408 24608
rect 5356 24565 5365 24599
rect 5365 24565 5399 24599
rect 5399 24565 5408 24599
rect 5356 24556 5408 24565
rect 9680 24556 9732 24608
rect 9956 24624 10008 24676
rect 12992 24624 13044 24676
rect 13176 24624 13228 24676
rect 14372 24667 14424 24676
rect 11428 24556 11480 24608
rect 13360 24556 13412 24608
rect 13544 24599 13596 24608
rect 13544 24565 13553 24599
rect 13553 24565 13587 24599
rect 13587 24565 13596 24599
rect 13544 24556 13596 24565
rect 13728 24556 13780 24608
rect 14004 24556 14056 24608
rect 14372 24633 14381 24667
rect 14381 24633 14415 24667
rect 14415 24633 14424 24667
rect 14372 24624 14424 24633
rect 15108 24624 15160 24676
rect 15660 24701 15669 24735
rect 15669 24701 15703 24735
rect 15703 24701 15712 24735
rect 15660 24692 15712 24701
rect 16856 24735 16908 24744
rect 16856 24701 16865 24735
rect 16865 24701 16899 24735
rect 16899 24701 16908 24735
rect 16856 24692 16908 24701
rect 17408 24760 17460 24812
rect 38016 24803 38068 24812
rect 17868 24692 17920 24744
rect 38016 24769 38025 24803
rect 38025 24769 38059 24803
rect 38059 24769 38068 24803
rect 38016 24760 38068 24769
rect 19892 24735 19944 24744
rect 19892 24701 19901 24735
rect 19901 24701 19935 24735
rect 19935 24701 19944 24735
rect 19892 24692 19944 24701
rect 20628 24692 20680 24744
rect 18512 24624 18564 24676
rect 18696 24624 18748 24676
rect 19340 24667 19392 24676
rect 19340 24633 19349 24667
rect 19349 24633 19383 24667
rect 19383 24633 19392 24667
rect 19340 24624 19392 24633
rect 17684 24556 17736 24608
rect 18144 24556 18196 24608
rect 38200 24599 38252 24608
rect 38200 24565 38209 24599
rect 38209 24565 38243 24599
rect 38243 24565 38252 24599
rect 38200 24556 38252 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 1952 24395 2004 24404
rect 1952 24361 1961 24395
rect 1961 24361 1995 24395
rect 1995 24361 2004 24395
rect 1952 24352 2004 24361
rect 2688 24352 2740 24404
rect 3976 24395 4028 24404
rect 3976 24361 3985 24395
rect 3985 24361 4019 24395
rect 4019 24361 4028 24395
rect 3976 24352 4028 24361
rect 5816 24352 5868 24404
rect 8576 24352 8628 24404
rect 8668 24352 8720 24404
rect 9680 24352 9732 24404
rect 13820 24352 13872 24404
rect 14004 24352 14056 24404
rect 17040 24352 17092 24404
rect 17500 24395 17552 24404
rect 17500 24361 17509 24395
rect 17509 24361 17543 24395
rect 17543 24361 17552 24395
rect 17500 24352 17552 24361
rect 18052 24395 18104 24404
rect 18052 24361 18061 24395
rect 18061 24361 18095 24395
rect 18095 24361 18104 24395
rect 18052 24352 18104 24361
rect 18328 24352 18380 24404
rect 19984 24352 20036 24404
rect 20076 24352 20128 24404
rect 1768 24284 1820 24336
rect 8484 24284 8536 24336
rect 2504 24191 2556 24200
rect 2504 24157 2513 24191
rect 2513 24157 2547 24191
rect 2547 24157 2556 24191
rect 8300 24216 8352 24268
rect 2504 24148 2556 24157
rect 7748 24191 7800 24200
rect 2780 24080 2832 24132
rect 7748 24157 7757 24191
rect 7757 24157 7791 24191
rect 7791 24157 7800 24191
rect 7748 24148 7800 24157
rect 7840 24148 7892 24200
rect 9312 24216 9364 24268
rect 13176 24284 13228 24336
rect 9680 24259 9732 24268
rect 9680 24225 9689 24259
rect 9689 24225 9723 24259
rect 9723 24225 9732 24259
rect 9680 24216 9732 24225
rect 12532 24216 12584 24268
rect 10692 24191 10744 24200
rect 10692 24157 10701 24191
rect 10701 24157 10735 24191
rect 10735 24157 10744 24191
rect 10692 24148 10744 24157
rect 10876 24191 10928 24200
rect 10876 24157 10885 24191
rect 10885 24157 10919 24191
rect 10919 24157 10928 24191
rect 10876 24148 10928 24157
rect 12256 24191 12308 24200
rect 12256 24157 12265 24191
rect 12265 24157 12299 24191
rect 12299 24157 12308 24191
rect 15568 24284 15620 24336
rect 13360 24216 13412 24268
rect 15660 24259 15712 24268
rect 12256 24148 12308 24157
rect 13636 24148 13688 24200
rect 8576 24080 8628 24132
rect 8944 24080 8996 24132
rect 4804 24055 4856 24064
rect 4804 24021 4813 24055
rect 4813 24021 4847 24055
rect 4847 24021 4856 24055
rect 4804 24012 4856 24021
rect 7196 24055 7248 24064
rect 7196 24021 7205 24055
rect 7205 24021 7239 24055
rect 7239 24021 7248 24055
rect 7196 24012 7248 24021
rect 8300 24012 8352 24064
rect 8760 24012 8812 24064
rect 9312 24123 9364 24132
rect 9312 24089 9321 24123
rect 9321 24089 9355 24123
rect 9355 24089 9364 24123
rect 15660 24225 15669 24259
rect 15669 24225 15703 24259
rect 15703 24225 15712 24259
rect 15660 24216 15712 24225
rect 16764 24216 16816 24268
rect 14648 24148 14700 24200
rect 20720 24284 20772 24336
rect 17868 24216 17920 24268
rect 9312 24080 9364 24089
rect 14924 24080 14976 24132
rect 9588 24012 9640 24064
rect 11704 24012 11756 24064
rect 14740 24012 14792 24064
rect 15752 24123 15804 24132
rect 15752 24089 15761 24123
rect 15761 24089 15795 24123
rect 15795 24089 15804 24123
rect 15752 24080 15804 24089
rect 18052 24148 18104 24200
rect 18328 24080 18380 24132
rect 16580 24012 16632 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 940 23808 992 23860
rect 2780 23808 2832 23860
rect 4068 23808 4120 23860
rect 4988 23808 5040 23860
rect 5264 23808 5316 23860
rect 11704 23851 11756 23860
rect 2136 23740 2188 23792
rect 7196 23740 7248 23792
rect 2504 23672 2556 23724
rect 7104 23715 7156 23724
rect 7104 23681 7113 23715
rect 7113 23681 7147 23715
rect 7147 23681 7156 23715
rect 7104 23672 7156 23681
rect 7748 23715 7800 23724
rect 7748 23681 7757 23715
rect 7757 23681 7791 23715
rect 7791 23681 7800 23715
rect 7748 23672 7800 23681
rect 9496 23740 9548 23792
rect 11704 23817 11713 23851
rect 11713 23817 11747 23851
rect 11747 23817 11756 23851
rect 11704 23808 11756 23817
rect 13360 23808 13412 23860
rect 15568 23808 15620 23860
rect 15752 23808 15804 23860
rect 17040 23808 17092 23860
rect 18328 23808 18380 23860
rect 11244 23740 11296 23792
rect 11612 23740 11664 23792
rect 13544 23740 13596 23792
rect 18144 23783 18196 23792
rect 18144 23749 18153 23783
rect 18153 23749 18187 23783
rect 18187 23749 18196 23783
rect 18144 23740 18196 23749
rect 18696 23783 18748 23792
rect 18696 23749 18705 23783
rect 18705 23749 18739 23783
rect 18739 23749 18748 23783
rect 18696 23740 18748 23749
rect 7840 23604 7892 23656
rect 4620 23536 4672 23588
rect 7196 23579 7248 23588
rect 7196 23545 7205 23579
rect 7205 23545 7239 23579
rect 7239 23545 7248 23579
rect 7196 23536 7248 23545
rect 2688 23468 2740 23520
rect 8852 23604 8904 23656
rect 9036 23647 9088 23656
rect 9036 23613 9045 23647
rect 9045 23613 9079 23647
rect 9079 23613 9088 23647
rect 9036 23604 9088 23613
rect 12256 23672 12308 23724
rect 14004 23672 14056 23724
rect 17040 23715 17092 23724
rect 17040 23681 17049 23715
rect 17049 23681 17083 23715
rect 17083 23681 17092 23715
rect 17040 23672 17092 23681
rect 10048 23604 10100 23656
rect 10324 23536 10376 23588
rect 11060 23604 11112 23656
rect 13820 23604 13872 23656
rect 14372 23536 14424 23588
rect 8576 23468 8628 23520
rect 13360 23468 13412 23520
rect 13636 23468 13688 23520
rect 15200 23579 15252 23588
rect 15200 23545 15209 23579
rect 15209 23545 15243 23579
rect 15243 23545 15252 23579
rect 16856 23604 16908 23656
rect 17776 23604 17828 23656
rect 15200 23536 15252 23545
rect 15384 23468 15436 23520
rect 27252 23808 27304 23860
rect 37280 23672 37332 23724
rect 17592 23468 17644 23520
rect 38200 23511 38252 23520
rect 38200 23477 38209 23511
rect 38209 23477 38243 23511
rect 38243 23477 38252 23511
rect 38200 23468 38252 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 2780 23264 2832 23316
rect 4620 23307 4672 23316
rect 4620 23273 4629 23307
rect 4629 23273 4663 23307
rect 4663 23273 4672 23307
rect 4620 23264 4672 23273
rect 5540 23264 5592 23316
rect 5724 23307 5776 23316
rect 5724 23273 5733 23307
rect 5733 23273 5767 23307
rect 5767 23273 5776 23307
rect 5724 23264 5776 23273
rect 6828 23264 6880 23316
rect 11060 23264 11112 23316
rect 11704 23264 11756 23316
rect 17684 23264 17736 23316
rect 27252 23307 27304 23316
rect 10692 23196 10744 23248
rect 14372 23239 14424 23248
rect 14372 23205 14381 23239
rect 14381 23205 14415 23239
rect 14415 23205 14424 23239
rect 14372 23196 14424 23205
rect 18604 23196 18656 23248
rect 9036 23128 9088 23180
rect 1768 23060 1820 23112
rect 10508 23128 10560 23180
rect 10784 23171 10836 23180
rect 10784 23137 10793 23171
rect 10793 23137 10827 23171
rect 10827 23137 10836 23171
rect 10784 23128 10836 23137
rect 11796 23128 11848 23180
rect 10968 23060 11020 23112
rect 12532 23103 12584 23112
rect 12532 23069 12541 23103
rect 12541 23069 12575 23103
rect 12575 23069 12584 23103
rect 12532 23060 12584 23069
rect 16764 23128 16816 23180
rect 27252 23273 27261 23307
rect 27261 23273 27295 23307
rect 27295 23273 27304 23307
rect 27252 23264 27304 23273
rect 27988 23307 28040 23316
rect 27988 23273 27997 23307
rect 27997 23273 28031 23307
rect 28031 23273 28040 23307
rect 27988 23264 28040 23273
rect 33692 23128 33744 23180
rect 10324 23035 10376 23044
rect 10324 23001 10333 23035
rect 10333 23001 10367 23035
rect 10367 23001 10376 23035
rect 10324 22992 10376 23001
rect 10416 23035 10468 23044
rect 10416 23001 10425 23035
rect 10425 23001 10459 23035
rect 10459 23001 10468 23035
rect 10416 22992 10468 23001
rect 11152 22992 11204 23044
rect 12348 22992 12400 23044
rect 14004 23060 14056 23112
rect 17868 23060 17920 23112
rect 27252 23060 27304 23112
rect 14096 22992 14148 23044
rect 15568 22992 15620 23044
rect 16028 23035 16080 23044
rect 16028 23001 16037 23035
rect 16037 23001 16071 23035
rect 16071 23001 16080 23035
rect 16028 22992 16080 23001
rect 16488 22992 16540 23044
rect 1860 22924 1912 22976
rect 11520 22967 11572 22976
rect 11520 22933 11529 22967
rect 11529 22933 11563 22967
rect 11563 22933 11572 22967
rect 11520 22924 11572 22933
rect 13360 22967 13412 22976
rect 13360 22933 13369 22967
rect 13369 22933 13403 22967
rect 13403 22933 13412 22967
rect 13360 22924 13412 22933
rect 17132 22924 17184 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 3148 22720 3200 22772
rect 3516 22720 3568 22772
rect 3884 22720 3936 22772
rect 5172 22720 5224 22772
rect 5448 22720 5500 22772
rect 5540 22720 5592 22772
rect 7748 22720 7800 22772
rect 10416 22720 10468 22772
rect 11520 22720 11572 22772
rect 5264 22652 5316 22704
rect 9312 22652 9364 22704
rect 10600 22652 10652 22704
rect 1860 22627 1912 22636
rect 1860 22593 1869 22627
rect 1869 22593 1903 22627
rect 1903 22593 1912 22627
rect 1860 22584 1912 22593
rect 3424 22584 3476 22636
rect 9588 22627 9640 22636
rect 9588 22593 9597 22627
rect 9597 22593 9631 22627
rect 9631 22593 9640 22627
rect 9588 22584 9640 22593
rect 10232 22627 10284 22636
rect 10232 22593 10241 22627
rect 10241 22593 10275 22627
rect 10275 22593 10284 22627
rect 10232 22584 10284 22593
rect 10508 22584 10560 22636
rect 6000 22559 6052 22568
rect 6000 22525 6009 22559
rect 6009 22525 6043 22559
rect 6043 22525 6052 22559
rect 6000 22516 6052 22525
rect 6552 22516 6604 22568
rect 1676 22491 1728 22500
rect 1676 22457 1685 22491
rect 1685 22457 1719 22491
rect 1719 22457 1728 22491
rect 1676 22448 1728 22457
rect 7932 22448 7984 22500
rect 17132 22695 17184 22704
rect 17132 22661 17141 22695
rect 17141 22661 17175 22695
rect 17175 22661 17184 22695
rect 17132 22652 17184 22661
rect 11244 22584 11296 22636
rect 12624 22584 12676 22636
rect 14740 22584 14792 22636
rect 15384 22627 15436 22636
rect 15384 22593 15393 22627
rect 15393 22593 15427 22627
rect 15427 22593 15436 22627
rect 15384 22584 15436 22593
rect 18328 22627 18380 22636
rect 18328 22593 18337 22627
rect 18337 22593 18371 22627
rect 18371 22593 18380 22627
rect 18328 22584 18380 22593
rect 2780 22380 2832 22432
rect 2964 22380 3016 22432
rect 13544 22516 13596 22568
rect 14096 22559 14148 22568
rect 14096 22525 14105 22559
rect 14105 22525 14139 22559
rect 14139 22525 14148 22559
rect 14096 22516 14148 22525
rect 17132 22516 17184 22568
rect 14372 22448 14424 22500
rect 15200 22448 15252 22500
rect 15568 22491 15620 22500
rect 15568 22457 15577 22491
rect 15577 22457 15611 22491
rect 15611 22457 15620 22491
rect 15568 22448 15620 22457
rect 16764 22448 16816 22500
rect 17868 22516 17920 22568
rect 19340 22559 19392 22568
rect 19340 22525 19349 22559
rect 19349 22525 19383 22559
rect 19383 22525 19392 22559
rect 19340 22516 19392 22525
rect 10968 22423 11020 22432
rect 10968 22389 10977 22423
rect 10977 22389 11011 22423
rect 11011 22389 11020 22423
rect 10968 22380 11020 22389
rect 12164 22423 12216 22432
rect 12164 22389 12173 22423
rect 12173 22389 12207 22423
rect 12207 22389 12216 22423
rect 12164 22380 12216 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 5264 22176 5316 22228
rect 6000 22219 6052 22228
rect 6000 22185 6009 22219
rect 6009 22185 6043 22219
rect 6043 22185 6052 22219
rect 6000 22176 6052 22185
rect 8852 22176 8904 22228
rect 9588 22176 9640 22228
rect 2780 22040 2832 22092
rect 4068 22040 4120 22092
rect 5080 22040 5132 22092
rect 7380 22040 7432 22092
rect 8208 22040 8260 22092
rect 10416 22083 10468 22092
rect 10416 22049 10425 22083
rect 10425 22049 10459 22083
rect 10459 22049 10468 22083
rect 10416 22040 10468 22049
rect 3516 21972 3568 22024
rect 4896 21972 4948 22024
rect 10600 21947 10652 21956
rect 10600 21913 10609 21947
rect 10609 21913 10643 21947
rect 10643 21913 10652 21947
rect 10600 21904 10652 21913
rect 10692 21947 10744 21956
rect 10692 21913 10701 21947
rect 10701 21913 10735 21947
rect 10735 21913 10744 21947
rect 10692 21904 10744 21913
rect 2964 21836 3016 21888
rect 10508 21836 10560 21888
rect 12348 22108 12400 22160
rect 11704 22040 11756 22092
rect 13360 22040 13412 22092
rect 13820 22040 13872 22092
rect 12624 22015 12676 22024
rect 12624 21981 12633 22015
rect 12633 21981 12667 22015
rect 12667 21981 12676 22015
rect 12624 21972 12676 21981
rect 15292 21972 15344 22024
rect 12072 21904 12124 21956
rect 13544 21836 13596 21888
rect 15660 21836 15712 21888
rect 17132 21836 17184 21888
rect 17776 21879 17828 21888
rect 17776 21845 17785 21879
rect 17785 21845 17819 21879
rect 17819 21845 17828 21879
rect 17776 21836 17828 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 2780 21632 2832 21684
rect 2872 21632 2924 21684
rect 4988 21675 5040 21684
rect 4988 21641 4997 21675
rect 4997 21641 5031 21675
rect 5031 21641 5040 21675
rect 4988 21632 5040 21641
rect 6184 21632 6236 21684
rect 6552 21675 6604 21684
rect 6552 21641 6561 21675
rect 6561 21641 6595 21675
rect 6595 21641 6604 21675
rect 6552 21632 6604 21641
rect 12164 21675 12216 21684
rect 12164 21641 12173 21675
rect 12173 21641 12207 21675
rect 12207 21641 12216 21675
rect 12164 21632 12216 21641
rect 6460 21564 6512 21616
rect 10600 21564 10652 21616
rect 10692 21564 10744 21616
rect 13912 21564 13964 21616
rect 14096 21607 14148 21616
rect 14096 21573 14105 21607
rect 14105 21573 14139 21607
rect 14139 21573 14148 21607
rect 14096 21564 14148 21573
rect 1584 21496 1636 21548
rect 5724 21496 5776 21548
rect 10508 21539 10560 21548
rect 10508 21505 10517 21539
rect 10517 21505 10551 21539
rect 10551 21505 10560 21539
rect 10508 21496 10560 21505
rect 10232 21428 10284 21480
rect 13268 21496 13320 21548
rect 15292 21496 15344 21548
rect 15660 21539 15712 21548
rect 15660 21505 15669 21539
rect 15669 21505 15703 21539
rect 15703 21505 15712 21539
rect 15660 21496 15712 21505
rect 36820 21496 36872 21548
rect 11060 21428 11112 21480
rect 11612 21428 11664 21480
rect 12808 21471 12860 21480
rect 12808 21437 12817 21471
rect 12817 21437 12851 21471
rect 12851 21437 12860 21471
rect 12808 21428 12860 21437
rect 15384 21428 15436 21480
rect 16028 21428 16080 21480
rect 16672 21428 16724 21480
rect 17868 21428 17920 21480
rect 15568 21360 15620 21412
rect 4620 21292 4672 21344
rect 11244 21292 11296 21344
rect 15108 21292 15160 21344
rect 38200 21335 38252 21344
rect 38200 21301 38209 21335
rect 38209 21301 38243 21335
rect 38243 21301 38252 21335
rect 38200 21292 38252 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 1584 21131 1636 21140
rect 1584 21097 1593 21131
rect 1593 21097 1627 21131
rect 1627 21097 1636 21131
rect 1584 21088 1636 21097
rect 2596 21088 2648 21140
rect 2872 21088 2924 21140
rect 4620 21131 4672 21140
rect 4620 21097 4629 21131
rect 4629 21097 4663 21131
rect 4663 21097 4672 21131
rect 4620 21088 4672 21097
rect 5264 21088 5316 21140
rect 11612 21131 11664 21140
rect 11612 21097 11621 21131
rect 11621 21097 11655 21131
rect 11655 21097 11664 21131
rect 11612 21088 11664 21097
rect 16672 21131 16724 21140
rect 16672 21097 16681 21131
rect 16681 21097 16715 21131
rect 16715 21097 16724 21131
rect 16672 21088 16724 21097
rect 18052 21088 18104 21140
rect 2688 21063 2740 21072
rect 2688 21029 2697 21063
rect 2697 21029 2731 21063
rect 2731 21029 2740 21063
rect 2688 21020 2740 21029
rect 26516 21020 26568 21072
rect 12808 20952 12860 21004
rect 13912 20952 13964 21004
rect 15476 20952 15528 21004
rect 11244 20884 11296 20936
rect 11520 20927 11572 20936
rect 11520 20893 11529 20927
rect 11529 20893 11563 20927
rect 11563 20893 11572 20927
rect 11520 20884 11572 20893
rect 13084 20927 13136 20936
rect 13084 20893 13093 20927
rect 13093 20893 13127 20927
rect 13127 20893 13136 20927
rect 13084 20884 13136 20893
rect 16948 20884 17000 20936
rect 18052 20884 18104 20936
rect 14832 20859 14884 20868
rect 14832 20825 14841 20859
rect 14841 20825 14875 20859
rect 14875 20825 14884 20859
rect 14832 20816 14884 20825
rect 15384 20816 15436 20868
rect 16672 20816 16724 20868
rect 20812 20816 20864 20868
rect 4896 20748 4948 20800
rect 10508 20748 10560 20800
rect 12072 20748 12124 20800
rect 12716 20748 12768 20800
rect 13544 20791 13596 20800
rect 13544 20757 13553 20791
rect 13553 20757 13587 20791
rect 13587 20757 13596 20791
rect 13544 20748 13596 20757
rect 15568 20791 15620 20800
rect 15568 20757 15577 20791
rect 15577 20757 15611 20791
rect 15611 20757 15620 20791
rect 15568 20748 15620 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 1584 20587 1636 20596
rect 1584 20553 1593 20587
rect 1593 20553 1627 20587
rect 1627 20553 1636 20587
rect 1584 20544 1636 20553
rect 2964 20544 3016 20596
rect 4068 20544 4120 20596
rect 5264 20587 5316 20596
rect 5264 20553 5273 20587
rect 5273 20553 5307 20587
rect 5307 20553 5316 20587
rect 5264 20544 5316 20553
rect 10324 20544 10376 20596
rect 11060 20587 11112 20596
rect 11060 20553 11069 20587
rect 11069 20553 11103 20587
rect 11103 20553 11112 20587
rect 11060 20544 11112 20553
rect 11520 20544 11572 20596
rect 12348 20544 12400 20596
rect 2780 20519 2832 20528
rect 2780 20485 2789 20519
rect 2789 20485 2823 20519
rect 2823 20485 2832 20519
rect 2780 20476 2832 20485
rect 3884 20476 3936 20528
rect 4896 20476 4948 20528
rect 6276 20476 6328 20528
rect 10508 20451 10560 20460
rect 10508 20417 10517 20451
rect 10517 20417 10551 20451
rect 10551 20417 10560 20451
rect 10508 20408 10560 20417
rect 10600 20408 10652 20460
rect 14832 20544 14884 20596
rect 16948 20587 17000 20596
rect 16948 20553 16957 20587
rect 16957 20553 16991 20587
rect 16991 20553 17000 20587
rect 16948 20544 17000 20553
rect 17868 20476 17920 20528
rect 10324 20340 10376 20392
rect 12164 20340 12216 20392
rect 15476 20408 15528 20460
rect 13544 20340 13596 20392
rect 15016 20383 15068 20392
rect 15016 20349 15025 20383
rect 15025 20349 15059 20383
rect 15059 20349 15068 20383
rect 15016 20340 15068 20349
rect 12440 20272 12492 20324
rect 13912 20272 13964 20324
rect 14832 20272 14884 20324
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 1676 20043 1728 20052
rect 1676 20009 1685 20043
rect 1685 20009 1719 20043
rect 1719 20009 1728 20043
rect 1676 20000 1728 20009
rect 2136 20000 2188 20052
rect 2872 20043 2924 20052
rect 2872 20009 2881 20043
rect 2881 20009 2915 20043
rect 2915 20009 2924 20043
rect 2872 20000 2924 20009
rect 3148 20000 3200 20052
rect 3332 20043 3384 20052
rect 3332 20009 3341 20043
rect 3341 20009 3375 20043
rect 3375 20009 3384 20043
rect 3332 20000 3384 20009
rect 4068 20043 4120 20052
rect 4068 20009 4077 20043
rect 4077 20009 4111 20043
rect 4111 20009 4120 20043
rect 4068 20000 4120 20009
rect 10876 20000 10928 20052
rect 12532 20000 12584 20052
rect 13084 20000 13136 20052
rect 16672 20043 16724 20052
rect 16672 20009 16681 20043
rect 16681 20009 16715 20043
rect 16715 20009 16724 20043
rect 16672 20000 16724 20009
rect 12348 19932 12400 19984
rect 12440 19796 12492 19848
rect 14832 19864 14884 19916
rect 16580 19864 16632 19916
rect 38108 19864 38160 19916
rect 3332 19728 3384 19780
rect 10968 19728 11020 19780
rect 12716 19728 12768 19780
rect 14740 19796 14792 19848
rect 38292 19839 38344 19848
rect 38292 19805 38301 19839
rect 38301 19805 38335 19839
rect 38335 19805 38344 19839
rect 38292 19796 38344 19805
rect 6184 19660 6236 19712
rect 10600 19703 10652 19712
rect 10600 19669 10609 19703
rect 10609 19669 10643 19703
rect 10643 19669 10652 19703
rect 10600 19660 10652 19669
rect 11244 19703 11296 19712
rect 11244 19669 11253 19703
rect 11253 19669 11287 19703
rect 11287 19669 11296 19703
rect 11244 19660 11296 19669
rect 14280 19703 14332 19712
rect 14280 19669 14289 19703
rect 14289 19669 14323 19703
rect 14323 19669 14332 19703
rect 14280 19660 14332 19669
rect 15108 19660 15160 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 10600 19456 10652 19508
rect 12440 19456 12492 19508
rect 12716 19499 12768 19508
rect 12716 19465 12725 19499
rect 12725 19465 12759 19499
rect 12759 19465 12768 19499
rect 12716 19456 12768 19465
rect 15016 19456 15068 19508
rect 11244 19388 11296 19440
rect 28540 19456 28592 19508
rect 38292 19499 38344 19508
rect 38292 19465 38301 19499
rect 38301 19465 38335 19499
rect 38335 19465 38344 19499
rect 38292 19456 38344 19465
rect 1584 19320 1636 19372
rect 14740 19320 14792 19372
rect 2320 19295 2372 19304
rect 2320 19261 2329 19295
rect 2329 19261 2363 19295
rect 2363 19261 2372 19295
rect 2320 19252 2372 19261
rect 13268 19295 13320 19304
rect 13268 19261 13277 19295
rect 13277 19261 13311 19295
rect 13311 19261 13320 19295
rect 13268 19252 13320 19261
rect 15200 19295 15252 19304
rect 15200 19261 15209 19295
rect 15209 19261 15243 19295
rect 15243 19261 15252 19295
rect 15200 19252 15252 19261
rect 15292 19184 15344 19236
rect 16028 19184 16080 19236
rect 1032 19116 1084 19168
rect 16580 19116 16632 19168
rect 17776 19116 17828 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1584 18955 1636 18964
rect 1584 18921 1593 18955
rect 1593 18921 1627 18955
rect 1627 18921 1636 18955
rect 1584 18912 1636 18921
rect 2228 18955 2280 18964
rect 2228 18921 2237 18955
rect 2237 18921 2271 18955
rect 2271 18921 2280 18955
rect 2228 18912 2280 18921
rect 5172 18912 5224 18964
rect 12440 18912 12492 18964
rect 19432 18912 19484 18964
rect 2780 18572 2832 18624
rect 22376 18572 22428 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 14280 18232 14332 18284
rect 38016 18232 38068 18284
rect 1676 18071 1728 18080
rect 1676 18037 1685 18071
rect 1685 18037 1719 18071
rect 1719 18037 1728 18071
rect 1676 18028 1728 18037
rect 17776 18028 17828 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 17868 17280 17920 17332
rect 7564 17144 7616 17196
rect 6736 16983 6788 16992
rect 6736 16949 6745 16983
rect 6745 16949 6779 16983
rect 6779 16949 6788 16983
rect 6736 16940 6788 16949
rect 24400 16940 24452 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 2780 16056 2832 16108
rect 37648 16056 37700 16108
rect 38292 16031 38344 16040
rect 38292 15997 38301 16031
rect 38301 15997 38335 16031
rect 38335 15997 38344 16031
rect 38292 15988 38344 15997
rect 1676 15895 1728 15904
rect 1676 15861 1685 15895
rect 1685 15861 1719 15895
rect 1719 15861 1728 15895
rect 1676 15852 1728 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 38292 15691 38344 15700
rect 38292 15657 38301 15691
rect 38301 15657 38335 15691
rect 38335 15657 38344 15691
rect 38292 15648 38344 15657
rect 10048 15444 10100 15496
rect 6828 15308 6880 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 4804 14560 4856 14612
rect 38016 14467 38068 14476
rect 38016 14433 38025 14467
rect 38025 14433 38059 14467
rect 38059 14433 38068 14467
rect 38016 14424 38068 14433
rect 38292 14399 38344 14408
rect 38292 14365 38301 14399
rect 38301 14365 38335 14399
rect 38335 14365 38344 14399
rect 38292 14356 38344 14365
rect 1952 14220 2004 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 38292 14059 38344 14068
rect 38292 14025 38301 14059
rect 38301 14025 38335 14059
rect 38335 14025 38344 14059
rect 38292 14016 38344 14025
rect 4712 13948 4764 14000
rect 1584 13880 1636 13932
rect 10324 13880 10376 13932
rect 2412 13855 2464 13864
rect 2412 13821 2421 13855
rect 2421 13821 2455 13855
rect 2455 13821 2464 13855
rect 2412 13812 2464 13821
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 1584 13515 1636 13524
rect 1584 13481 1593 13515
rect 1593 13481 1627 13515
rect 1627 13481 1636 13515
rect 1584 13472 1636 13481
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 6736 12792 6788 12844
rect 38200 12835 38252 12844
rect 38200 12801 38209 12835
rect 38209 12801 38243 12835
rect 38243 12801 38252 12835
rect 38200 12792 38252 12801
rect 37280 12656 37332 12708
rect 1676 12631 1728 12640
rect 1676 12597 1685 12631
rect 1685 12597 1719 12631
rect 1719 12597 1728 12631
rect 1676 12588 1728 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 15384 12384 15436 12436
rect 38016 12180 38068 12232
rect 16120 12087 16172 12096
rect 16120 12053 16129 12087
rect 16129 12053 16163 12087
rect 16163 12053 16172 12087
rect 16120 12044 16172 12053
rect 38016 12087 38068 12096
rect 38016 12053 38025 12087
rect 38025 12053 38059 12087
rect 38059 12053 38068 12087
rect 38016 12044 38068 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 8392 11092 8444 11144
rect 37832 11092 37884 11144
rect 10876 11067 10928 11076
rect 10876 11033 10885 11067
rect 10885 11033 10919 11067
rect 10919 11033 10928 11067
rect 10876 11024 10928 11033
rect 38200 11067 38252 11076
rect 38200 11033 38209 11067
rect 38209 11033 38243 11067
rect 38243 11033 38252 11067
rect 38200 11024 38252 11033
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 8944 10795 8996 10804
rect 8944 10761 8953 10795
rect 8953 10761 8987 10795
rect 8987 10761 8996 10795
rect 8944 10752 8996 10761
rect 12624 10752 12676 10804
rect 19984 10752 20036 10804
rect 2412 10616 2464 10668
rect 8668 10616 8720 10668
rect 1676 10455 1728 10464
rect 1676 10421 1685 10455
rect 1685 10421 1719 10455
rect 1719 10421 1728 10455
rect 1676 10412 1728 10421
rect 14372 10616 14424 10668
rect 29000 10616 29052 10668
rect 22008 10480 22060 10532
rect 12716 10412 12768 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 16856 10251 16908 10260
rect 16856 10217 16865 10251
rect 16865 10217 16899 10251
rect 16899 10217 16908 10251
rect 16856 10208 16908 10217
rect 16856 10004 16908 10056
rect 18604 9936 18656 9988
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 18144 9052 18196 9104
rect 13360 8916 13412 8968
rect 16028 8916 16080 8968
rect 38016 8959 38068 8968
rect 38016 8925 38025 8959
rect 38025 8925 38059 8959
rect 38059 8925 38068 8959
rect 38016 8916 38068 8925
rect 1676 8891 1728 8900
rect 1676 8857 1685 8891
rect 1685 8857 1719 8891
rect 1719 8857 1728 8891
rect 1676 8848 1728 8857
rect 13636 8780 13688 8832
rect 16856 8848 16908 8900
rect 38200 8823 38252 8832
rect 38200 8789 38209 8823
rect 38209 8789 38243 8823
rect 38243 8789 38252 8823
rect 38200 8780 38252 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 1676 8619 1728 8628
rect 1676 8585 1685 8619
rect 1685 8585 1719 8619
rect 1719 8585 1728 8619
rect 1676 8576 1728 8585
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 22376 7395 22428 7404
rect 22376 7361 22385 7395
rect 22385 7361 22419 7395
rect 22419 7361 22428 7395
rect 22376 7352 22428 7361
rect 37280 7488 37332 7540
rect 37924 7420 37976 7472
rect 38200 7395 38252 7404
rect 38200 7361 38209 7395
rect 38209 7361 38243 7395
rect 38243 7361 38252 7395
rect 38200 7352 38252 7361
rect 1584 7327 1636 7336
rect 1584 7293 1593 7327
rect 1593 7293 1627 7327
rect 1627 7293 1636 7327
rect 1584 7284 1636 7293
rect 10508 7284 10560 7336
rect 22560 7191 22612 7200
rect 22560 7157 22569 7191
rect 22569 7157 22603 7191
rect 22603 7157 22612 7191
rect 22560 7148 22612 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 1584 6987 1636 6996
rect 1584 6953 1593 6987
rect 1593 6953 1627 6987
rect 1627 6953 1636 6987
rect 1584 6944 1636 6953
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 24400 6307 24452 6316
rect 24400 6273 24409 6307
rect 24409 6273 24443 6307
rect 24443 6273 24452 6307
rect 24400 6264 24452 6273
rect 24952 6060 25004 6112
rect 37832 6060 37884 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 38384 5856 38436 5908
rect 38200 5627 38252 5636
rect 38200 5593 38209 5627
rect 38209 5593 38243 5627
rect 38243 5593 38252 5627
rect 38200 5584 38252 5593
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 1768 5355 1820 5364
rect 1768 5321 1777 5355
rect 1777 5321 1811 5355
rect 1811 5321 1820 5355
rect 1768 5312 1820 5321
rect 1584 5176 1636 5228
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 1584 4811 1636 4820
rect 1584 4777 1593 4811
rect 1593 4777 1627 4811
rect 1627 4777 1636 4811
rect 1584 4768 1636 4777
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 1676 3927 1728 3936
rect 1676 3893 1685 3927
rect 1685 3893 1719 3927
rect 1719 3893 1728 3927
rect 1676 3884 1728 3893
rect 38108 3884 38160 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 2872 3612 2924 3664
rect 1676 3519 1728 3528
rect 1676 3485 1685 3519
rect 1685 3485 1719 3519
rect 1719 3485 1728 3519
rect 1676 3476 1728 3485
rect 37372 3340 37424 3392
rect 38200 3383 38252 3392
rect 38200 3349 38209 3383
rect 38209 3349 38243 3383
rect 38243 3349 38252 3383
rect 38200 3340 38252 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 12716 3179 12768 3188
rect 12716 3145 12725 3179
rect 12725 3145 12759 3179
rect 12759 3145 12768 3179
rect 12716 3136 12768 3145
rect 15936 3136 15988 3188
rect 34704 3179 34756 3188
rect 1952 3000 2004 3052
rect 8668 3043 8720 3052
rect 8668 3009 8677 3043
rect 8677 3009 8711 3043
rect 8711 3009 8720 3043
rect 8668 3000 8720 3009
rect 14924 3068 14976 3120
rect 20628 3068 20680 3120
rect 2412 2975 2464 2984
rect 2412 2941 2421 2975
rect 2421 2941 2455 2975
rect 2455 2941 2464 2975
rect 2412 2932 2464 2941
rect 15568 2932 15620 2984
rect 15752 3000 15804 3052
rect 16120 3000 16172 3052
rect 20812 3068 20864 3120
rect 34704 3145 34713 3179
rect 34713 3145 34747 3179
rect 34747 3145 34756 3179
rect 34704 3136 34756 3145
rect 29000 3043 29052 3052
rect 29000 3009 29009 3043
rect 29009 3009 29043 3043
rect 29043 3009 29052 3043
rect 37280 3068 37332 3120
rect 37740 3068 37792 3120
rect 29000 3000 29052 3009
rect 38200 3043 38252 3052
rect 38200 3009 38209 3043
rect 38209 3009 38243 3043
rect 38243 3009 38252 3043
rect 38200 3000 38252 3009
rect 30288 2932 30340 2984
rect 36728 2932 36780 2984
rect 4712 2864 4764 2916
rect 37372 2864 37424 2916
rect 1676 2839 1728 2848
rect 1676 2805 1685 2839
rect 1685 2805 1719 2839
rect 1719 2805 1728 2839
rect 1676 2796 1728 2805
rect 4620 2796 4672 2848
rect 8576 2796 8628 2848
rect 23388 2796 23440 2848
rect 29184 2839 29236 2848
rect 29184 2805 29193 2839
rect 29193 2805 29227 2839
rect 29227 2805 29236 2839
rect 29184 2796 29236 2805
rect 36360 2839 36412 2848
rect 36360 2805 36369 2839
rect 36369 2805 36403 2839
rect 36403 2805 36412 2839
rect 36360 2796 36412 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 8668 2592 8720 2644
rect 20 2524 72 2576
rect 2964 2524 3016 2576
rect 2412 2388 2464 2440
rect 4712 2456 4764 2508
rect 15752 2592 15804 2644
rect 28540 2635 28592 2644
rect 28540 2601 28549 2635
rect 28549 2601 28583 2635
rect 28583 2601 28592 2635
rect 28540 2592 28592 2601
rect 33692 2635 33744 2644
rect 33692 2601 33701 2635
rect 33701 2601 33735 2635
rect 33735 2601 33744 2635
rect 33692 2592 33744 2601
rect 11980 2567 12032 2576
rect 11980 2533 11989 2567
rect 11989 2533 12023 2567
rect 12023 2533 12032 2567
rect 11980 2524 12032 2533
rect 15660 2524 15712 2576
rect 30288 2524 30340 2576
rect 15384 2456 15436 2508
rect 34796 2524 34848 2576
rect 37280 2456 37332 2508
rect 1308 2252 1360 2304
rect 3240 2252 3292 2304
rect 6828 2431 6880 2440
rect 6828 2397 6837 2431
rect 6837 2397 6871 2431
rect 6871 2397 6880 2431
rect 6828 2388 6880 2397
rect 8576 2431 8628 2440
rect 8576 2397 8585 2431
rect 8585 2397 8619 2431
rect 8619 2397 8628 2431
rect 8576 2388 8628 2397
rect 9680 2388 9732 2440
rect 10876 2388 10928 2440
rect 16856 2431 16908 2440
rect 16856 2397 16865 2431
rect 16865 2397 16899 2431
rect 16899 2397 16908 2431
rect 16856 2388 16908 2397
rect 18144 2431 18196 2440
rect 18144 2397 18153 2431
rect 18153 2397 18187 2431
rect 18187 2397 18196 2431
rect 18144 2388 18196 2397
rect 18604 2388 18656 2440
rect 22008 2431 22060 2440
rect 22008 2397 22017 2431
rect 22017 2397 22051 2431
rect 22051 2397 22060 2431
rect 22008 2388 22060 2397
rect 22560 2388 22612 2440
rect 24952 2388 25004 2440
rect 4528 2320 4580 2372
rect 11612 2320 11664 2372
rect 14832 2320 14884 2372
rect 23388 2320 23440 2372
rect 29184 2388 29236 2440
rect 34704 2388 34756 2440
rect 36360 2388 36412 2440
rect 37188 2388 37240 2440
rect 38108 2388 38160 2440
rect 28356 2320 28408 2372
rect 33508 2320 33560 2372
rect 36728 2320 36780 2372
rect 6460 2252 6512 2304
rect 8392 2295 8444 2304
rect 8392 2261 8401 2295
rect 8401 2261 8435 2295
rect 8435 2261 8444 2295
rect 8392 2252 8444 2261
rect 12900 2252 12952 2304
rect 16764 2252 16816 2304
rect 18052 2252 18104 2304
rect 19984 2252 20036 2304
rect 21272 2252 21324 2304
rect 23204 2252 23256 2304
rect 25136 2252 25188 2304
rect 26424 2252 26476 2304
rect 29644 2252 29696 2304
rect 31760 2295 31812 2304
rect 31760 2261 31769 2295
rect 31769 2261 31803 2295
rect 31803 2261 31812 2295
rect 31760 2252 31812 2261
rect 34796 2252 34848 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 18 39200 74 39800
rect 1950 39200 2006 39800
rect 3882 39200 3938 39800
rect 5170 39200 5226 39800
rect 7102 39200 7158 39800
rect 7208 39222 7420 39250
rect 32 37330 60 39200
rect 20 37324 72 37330
rect 20 37266 72 37272
rect 1676 37256 1728 37262
rect 1676 37198 1728 37204
rect 1688 36922 1716 37198
rect 1860 37188 1912 37194
rect 1860 37130 1912 37136
rect 1676 36916 1728 36922
rect 1676 36858 1728 36864
rect 940 36848 992 36854
rect 940 36790 992 36796
rect 848 29028 900 29034
rect 848 28970 900 28976
rect 860 26450 888 28970
rect 848 26444 900 26450
rect 848 26386 900 26392
rect 952 23866 980 36790
rect 1688 36174 1716 36858
rect 1676 36168 1728 36174
rect 1676 36110 1728 36116
rect 1308 35760 1360 35766
rect 1308 35702 1360 35708
rect 1124 33856 1176 33862
rect 1124 33798 1176 33804
rect 1032 33516 1084 33522
rect 1032 33458 1084 33464
rect 940 23860 992 23866
rect 940 23802 992 23808
rect 1044 19174 1072 33458
rect 1136 24682 1164 33798
rect 1216 32768 1268 32774
rect 1216 32710 1268 32716
rect 1228 25498 1256 32710
rect 1320 26518 1348 35702
rect 1688 35698 1716 36110
rect 1872 35894 1900 37130
rect 1780 35866 1900 35894
rect 1676 35692 1728 35698
rect 1676 35634 1728 35640
rect 1676 32428 1728 32434
rect 1676 32370 1728 32376
rect 1688 32337 1716 32370
rect 1674 32328 1730 32337
rect 1674 32263 1730 32272
rect 1674 31376 1730 31385
rect 1674 31311 1676 31320
rect 1728 31311 1730 31320
rect 1676 31282 1728 31288
rect 1780 30598 1808 35866
rect 1964 34542 1992 39200
rect 3054 38856 3110 38865
rect 3054 38791 3110 38800
rect 2320 37324 2372 37330
rect 2320 37266 2372 37272
rect 2044 35080 2096 35086
rect 2044 35022 2096 35028
rect 1952 34536 2004 34542
rect 1952 34478 2004 34484
rect 1858 31240 1914 31249
rect 1858 31175 1860 31184
rect 1912 31175 1914 31184
rect 1860 31146 1912 31152
rect 1768 30592 1820 30598
rect 1768 30534 1820 30540
rect 2056 30410 2084 35022
rect 2332 32298 2360 37266
rect 2688 37188 2740 37194
rect 2688 37130 2740 37136
rect 2412 35624 2464 35630
rect 2412 35566 2464 35572
rect 2424 34950 2452 35566
rect 2412 34944 2464 34950
rect 2412 34886 2464 34892
rect 2320 32292 2372 32298
rect 2320 32234 2372 32240
rect 2136 31748 2188 31754
rect 2136 31690 2188 31696
rect 1964 30382 2084 30410
rect 1674 30152 1730 30161
rect 1730 30110 1808 30138
rect 1674 30087 1676 30096
rect 1728 30087 1730 30096
rect 1676 30058 1728 30064
rect 1674 30016 1730 30025
rect 1674 29951 1730 29960
rect 1688 29238 1716 29951
rect 1676 29232 1728 29238
rect 1676 29174 1728 29180
rect 1688 28506 1716 29174
rect 1780 29170 1808 30110
rect 1768 29164 1820 29170
rect 1768 29106 1820 29112
rect 1780 29073 1808 29106
rect 1766 29064 1822 29073
rect 1766 28999 1822 29008
rect 1596 28478 1716 28506
rect 1860 28484 1912 28490
rect 1308 26512 1360 26518
rect 1308 26454 1360 26460
rect 1216 25492 1268 25498
rect 1216 25434 1268 25440
rect 1124 24676 1176 24682
rect 1124 24618 1176 24624
rect 1596 22386 1624 28478
rect 1860 28426 1912 28432
rect 1674 27976 1730 27985
rect 1674 27911 1676 27920
rect 1728 27911 1730 27920
rect 1676 27882 1728 27888
rect 1768 26988 1820 26994
rect 1768 26930 1820 26936
rect 1676 26784 1728 26790
rect 1676 26726 1728 26732
rect 1688 26625 1716 26726
rect 1674 26616 1730 26625
rect 1674 26551 1730 26560
rect 1676 24608 1728 24614
rect 1674 24576 1676 24585
rect 1728 24576 1730 24585
rect 1674 24511 1730 24520
rect 1780 24342 1808 26930
rect 1872 26330 1900 28426
rect 1964 27452 1992 30382
rect 2044 30252 2096 30258
rect 2044 30194 2096 30200
rect 2056 27606 2084 30194
rect 2044 27600 2096 27606
rect 2044 27542 2096 27548
rect 1964 27424 2084 27452
rect 1872 26314 1992 26330
rect 1872 26308 2004 26314
rect 1872 26302 1952 26308
rect 1952 26250 2004 26256
rect 2056 26042 2084 27424
rect 2148 26586 2176 31690
rect 2228 31340 2280 31346
rect 2228 31282 2280 31288
rect 2136 26580 2188 26586
rect 2136 26522 2188 26528
rect 2136 26308 2188 26314
rect 2136 26250 2188 26256
rect 2044 26036 2096 26042
rect 2044 25978 2096 25984
rect 1950 24712 2006 24721
rect 1950 24647 2006 24656
rect 1964 24410 1992 24647
rect 1952 24404 2004 24410
rect 1952 24346 2004 24352
rect 1768 24336 1820 24342
rect 1768 24278 1820 24284
rect 2148 23798 2176 26250
rect 2240 26234 2268 31282
rect 2320 31136 2372 31142
rect 2320 31078 2372 31084
rect 2332 28082 2360 31078
rect 2320 28076 2372 28082
rect 2320 28018 2372 28024
rect 2320 26920 2372 26926
rect 2320 26862 2372 26868
rect 2332 26382 2360 26862
rect 2424 26586 2452 34886
rect 2504 34196 2556 34202
rect 2504 34138 2556 34144
rect 2516 33289 2544 34138
rect 2502 33280 2558 33289
rect 2502 33215 2558 33224
rect 2596 32428 2648 32434
rect 2596 32370 2648 32376
rect 2608 31793 2636 32370
rect 2594 31784 2650 31793
rect 2594 31719 2650 31728
rect 2596 31340 2648 31346
rect 2596 31282 2648 31288
rect 2504 30660 2556 30666
rect 2504 30602 2556 30608
rect 2516 27130 2544 30602
rect 2608 28558 2636 31282
rect 2596 28552 2648 28558
rect 2596 28494 2648 28500
rect 2504 27124 2556 27130
rect 2504 27066 2556 27072
rect 2504 26988 2556 26994
rect 2504 26930 2556 26936
rect 2412 26580 2464 26586
rect 2412 26522 2464 26528
rect 2320 26376 2372 26382
rect 2320 26318 2372 26324
rect 2412 26240 2464 26246
rect 2240 26206 2360 26234
rect 2136 23792 2188 23798
rect 2136 23734 2188 23740
rect 1768 23112 1820 23118
rect 1768 23054 1820 23060
rect 1674 22536 1730 22545
rect 1674 22471 1676 22480
rect 1728 22471 1730 22480
rect 1676 22442 1728 22448
rect 1596 22358 1716 22386
rect 1584 21548 1636 21554
rect 1584 21490 1636 21496
rect 1596 21185 1624 21490
rect 1582 21176 1638 21185
rect 1582 21111 1584 21120
rect 1636 21111 1638 21120
rect 1584 21082 1636 21088
rect 1582 20632 1638 20641
rect 1582 20567 1584 20576
rect 1636 20567 1638 20576
rect 1584 20538 1636 20544
rect 1688 20058 1716 22358
rect 1676 20052 1728 20058
rect 1676 19994 1728 20000
rect 1584 19372 1636 19378
rect 1584 19314 1636 19320
rect 1032 19168 1084 19174
rect 1596 19145 1624 19314
rect 1032 19110 1084 19116
rect 1582 19136 1638 19145
rect 1582 19071 1638 19080
rect 1596 18970 1624 19071
rect 1584 18964 1636 18970
rect 1584 18906 1636 18912
rect 1676 18080 1728 18086
rect 1676 18022 1728 18028
rect 1688 17785 1716 18022
rect 1674 17776 1730 17785
rect 1674 17711 1730 17720
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 1688 15745 1716 15846
rect 1674 15736 1730 15745
rect 1674 15671 1730 15680
rect 1584 13932 1636 13938
rect 1584 13874 1636 13880
rect 1596 13705 1624 13874
rect 1582 13696 1638 13705
rect 1582 13631 1638 13640
rect 1596 13530 1624 13631
rect 1584 13524 1636 13530
rect 1584 13466 1636 13472
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 1688 12345 1716 12582
rect 1674 12336 1730 12345
rect 1674 12271 1730 12280
rect 1676 10464 1728 10470
rect 1676 10406 1728 10412
rect 1688 10305 1716 10406
rect 1674 10296 1730 10305
rect 1674 10231 1730 10240
rect 1674 8936 1730 8945
rect 1674 8871 1676 8880
rect 1728 8871 1730 8880
rect 1676 8842 1728 8848
rect 1688 8634 1716 8842
rect 1676 8628 1728 8634
rect 1676 8570 1728 8576
rect 1584 7336 1636 7342
rect 1584 7278 1636 7284
rect 1596 7002 1624 7278
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1596 6905 1624 6938
rect 1582 6896 1638 6905
rect 1582 6831 1638 6840
rect 1780 5370 1808 23054
rect 1860 22976 1912 22982
rect 1860 22918 1912 22924
rect 1872 22642 1900 22918
rect 1860 22636 1912 22642
rect 1860 22578 1912 22584
rect 2148 20058 2176 23734
rect 2136 20052 2188 20058
rect 2136 19994 2188 20000
rect 2332 19310 2360 26206
rect 2412 26182 2464 26188
rect 2424 25702 2452 26182
rect 2412 25696 2464 25702
rect 2412 25638 2464 25644
rect 2516 25294 2544 26930
rect 2504 25288 2556 25294
rect 2504 25230 2556 25236
rect 2516 24614 2544 25230
rect 2504 24608 2556 24614
rect 2504 24550 2556 24556
rect 2516 24206 2544 24550
rect 2504 24200 2556 24206
rect 2504 24142 2556 24148
rect 2516 23730 2544 24142
rect 2504 23724 2556 23730
rect 2504 23666 2556 23672
rect 2608 21146 2636 28494
rect 2700 24410 2728 37130
rect 2778 36816 2834 36825
rect 2778 36751 2834 36760
rect 2792 33590 2820 36751
rect 2964 36100 3016 36106
rect 2964 36042 3016 36048
rect 2976 36009 3004 36042
rect 2962 36000 3018 36009
rect 2962 35935 3018 35944
rect 2964 34060 3016 34066
rect 2964 34002 3016 34008
rect 2780 33584 2832 33590
rect 2780 33526 2832 33532
rect 2870 33552 2926 33561
rect 2870 33487 2872 33496
rect 2924 33487 2926 33496
rect 2872 33458 2924 33464
rect 2976 32978 3004 34002
rect 2964 32972 3016 32978
rect 2964 32914 3016 32920
rect 2976 32570 3004 32914
rect 2964 32564 3016 32570
rect 2964 32506 3016 32512
rect 2872 32496 2924 32502
rect 2872 32438 2924 32444
rect 2780 32020 2832 32026
rect 2884 32008 2912 32438
rect 2976 32026 3004 32506
rect 3068 32337 3096 38791
rect 3896 37194 3924 39200
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 5184 37312 5212 39200
rect 7116 39114 7144 39200
rect 7208 39114 7236 39222
rect 7116 39086 7236 39114
rect 5092 37284 5212 37312
rect 6552 37324 6604 37330
rect 4620 37256 4672 37262
rect 4620 37198 4672 37204
rect 3884 37188 3936 37194
rect 3884 37130 3936 37136
rect 3332 37120 3384 37126
rect 3332 37062 3384 37068
rect 3148 34672 3200 34678
rect 3148 34614 3200 34620
rect 3054 32328 3110 32337
rect 3054 32263 3110 32272
rect 2832 31980 2912 32008
rect 2964 32020 3016 32026
rect 2780 31962 2832 31968
rect 2964 31962 3016 31968
rect 3160 31754 3188 34614
rect 3344 33114 3372 37062
rect 3896 36922 3924 37130
rect 4252 37120 4304 37126
rect 4252 37062 4304 37068
rect 3884 36916 3936 36922
rect 3884 36858 3936 36864
rect 3896 36786 3924 36858
rect 3884 36780 3936 36786
rect 3884 36722 3936 36728
rect 3896 36242 3924 36722
rect 4068 36712 4120 36718
rect 4068 36654 4120 36660
rect 3700 36236 3752 36242
rect 3700 36178 3752 36184
rect 3884 36236 3936 36242
rect 3884 36178 3936 36184
rect 3712 35494 3740 36178
rect 3896 35834 3924 36178
rect 3976 36168 4028 36174
rect 3976 36110 4028 36116
rect 3884 35828 3936 35834
rect 3884 35770 3936 35776
rect 3700 35488 3752 35494
rect 3700 35430 3752 35436
rect 3792 35216 3844 35222
rect 3792 35158 3844 35164
rect 3424 35148 3476 35154
rect 3424 35090 3476 35096
rect 3436 34066 3464 35090
rect 3700 35080 3752 35086
rect 3700 35022 3752 35028
rect 3712 34678 3740 35022
rect 3804 34746 3832 35158
rect 3896 35154 3924 35770
rect 3988 35290 4016 36110
rect 4080 36038 4108 36654
rect 4264 36582 4292 37062
rect 4252 36576 4304 36582
rect 4252 36518 4304 36524
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4632 36378 4660 37198
rect 4988 36576 5040 36582
rect 4988 36518 5040 36524
rect 4620 36372 4672 36378
rect 4620 36314 4672 36320
rect 5000 36106 5028 36518
rect 4988 36100 5040 36106
rect 4988 36042 5040 36048
rect 4068 36032 4120 36038
rect 4068 35974 4120 35980
rect 5000 35630 5028 36042
rect 4988 35624 5040 35630
rect 4988 35566 5040 35572
rect 4712 35556 4764 35562
rect 4712 35498 4764 35504
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 3976 35284 4028 35290
rect 3976 35226 4028 35232
rect 3884 35148 3936 35154
rect 3884 35090 3936 35096
rect 3896 34746 3924 35090
rect 3988 35086 4016 35226
rect 3976 35080 4028 35086
rect 3976 35022 4028 35028
rect 3976 34944 4028 34950
rect 3976 34886 4028 34892
rect 3792 34740 3844 34746
rect 3792 34682 3844 34688
rect 3884 34740 3936 34746
rect 3884 34682 3936 34688
rect 3700 34672 3752 34678
rect 3700 34614 3752 34620
rect 3700 34536 3752 34542
rect 3700 34478 3752 34484
rect 3424 34060 3476 34066
rect 3424 34002 3476 34008
rect 3424 33856 3476 33862
rect 3424 33798 3476 33804
rect 3436 33522 3464 33798
rect 3424 33516 3476 33522
rect 3424 33458 3476 33464
rect 3332 33108 3384 33114
rect 3332 33050 3384 33056
rect 3344 33017 3372 33050
rect 3330 33008 3386 33017
rect 3330 32943 3386 32952
rect 3436 32178 3464 33458
rect 3712 32881 3740 34478
rect 3792 33312 3844 33318
rect 3792 33254 3844 33260
rect 3698 32872 3754 32881
rect 3698 32807 3754 32816
rect 3698 32600 3754 32609
rect 3698 32535 3754 32544
rect 3516 32496 3568 32502
rect 3516 32438 3568 32444
rect 2976 31726 3188 31754
rect 3344 32150 3464 32178
rect 2872 28484 2924 28490
rect 2872 28426 2924 28432
rect 2884 27674 2912 28426
rect 2872 27668 2924 27674
rect 2872 27610 2924 27616
rect 2872 27532 2924 27538
rect 2872 27474 2924 27480
rect 2884 27441 2912 27474
rect 2870 27432 2926 27441
rect 2870 27367 2926 27376
rect 2780 26376 2832 26382
rect 2780 26318 2832 26324
rect 2792 25906 2820 26318
rect 2780 25900 2832 25906
rect 2780 25842 2832 25848
rect 2792 25294 2820 25842
rect 2780 25288 2832 25294
rect 2780 25230 2832 25236
rect 2792 24818 2820 25230
rect 2780 24812 2832 24818
rect 2780 24754 2832 24760
rect 2688 24404 2740 24410
rect 2688 24346 2740 24352
rect 2792 24138 2820 24754
rect 2780 24132 2832 24138
rect 2780 24074 2832 24080
rect 2792 23866 2820 24074
rect 2780 23860 2832 23866
rect 2780 23802 2832 23808
rect 2688 23520 2740 23526
rect 2688 23462 2740 23468
rect 2596 21140 2648 21146
rect 2596 21082 2648 21088
rect 2700 21078 2728 23462
rect 2792 23322 2820 23802
rect 2780 23316 2832 23322
rect 2780 23258 2832 23264
rect 2792 22438 2820 23258
rect 2780 22432 2832 22438
rect 2780 22374 2832 22380
rect 2780 22092 2832 22098
rect 2780 22034 2832 22040
rect 2792 21690 2820 22034
rect 2884 21690 2912 27367
rect 2976 26994 3004 31726
rect 3148 31408 3200 31414
rect 3148 31350 3200 31356
rect 3056 29232 3108 29238
rect 3056 29174 3108 29180
rect 3068 27130 3096 29174
rect 3160 29102 3188 31350
rect 3240 30592 3292 30598
rect 3240 30534 3292 30540
rect 3148 29096 3200 29102
rect 3148 29038 3200 29044
rect 3148 28008 3200 28014
rect 3148 27950 3200 27956
rect 3056 27124 3108 27130
rect 3056 27066 3108 27072
rect 2964 26988 3016 26994
rect 2964 26930 3016 26936
rect 2976 25838 3004 26930
rect 3056 26784 3108 26790
rect 3056 26726 3108 26732
rect 3068 26450 3096 26726
rect 3160 26450 3188 27950
rect 3252 26994 3280 30534
rect 3344 28082 3372 32150
rect 3424 32020 3476 32026
rect 3424 31962 3476 31968
rect 3436 31822 3464 31962
rect 3424 31816 3476 31822
rect 3424 31758 3476 31764
rect 3436 30734 3464 31758
rect 3424 30728 3476 30734
rect 3424 30670 3476 30676
rect 3424 30184 3476 30190
rect 3424 30126 3476 30132
rect 3436 29714 3464 30126
rect 3424 29708 3476 29714
rect 3424 29650 3476 29656
rect 3424 28960 3476 28966
rect 3424 28902 3476 28908
rect 3436 28558 3464 28902
rect 3424 28552 3476 28558
rect 3424 28494 3476 28500
rect 3332 28076 3384 28082
rect 3332 28018 3384 28024
rect 3240 26988 3292 26994
rect 3240 26930 3292 26936
rect 3056 26444 3108 26450
rect 3056 26386 3108 26392
rect 3148 26444 3200 26450
rect 3148 26386 3200 26392
rect 3148 26240 3200 26246
rect 3148 26182 3200 26188
rect 3160 25906 3188 26182
rect 3148 25900 3200 25906
rect 3148 25842 3200 25848
rect 2964 25832 3016 25838
rect 2964 25774 3016 25780
rect 2976 25362 3004 25774
rect 3160 25702 3188 25842
rect 3148 25696 3200 25702
rect 3148 25638 3200 25644
rect 2964 25356 3016 25362
rect 2964 25298 3016 25304
rect 3160 22778 3188 25638
rect 3148 22772 3200 22778
rect 3148 22714 3200 22720
rect 3436 22642 3464 28494
rect 3528 25498 3556 32438
rect 3712 32298 3740 32535
rect 3804 32348 3832 33254
rect 3884 32360 3936 32366
rect 3804 32320 3884 32348
rect 3700 32292 3752 32298
rect 3700 32234 3752 32240
rect 3608 31884 3660 31890
rect 3608 31826 3660 31832
rect 3620 30054 3648 31826
rect 3712 30326 3740 32234
rect 3700 30320 3752 30326
rect 3700 30262 3752 30268
rect 3608 30048 3660 30054
rect 3608 29990 3660 29996
rect 3608 29640 3660 29646
rect 3608 29582 3660 29588
rect 3620 27334 3648 29582
rect 3712 27470 3740 30262
rect 3804 30258 3832 32320
rect 3884 32302 3936 32308
rect 3882 31920 3938 31929
rect 3988 31906 4016 34886
rect 4620 34672 4672 34678
rect 4618 34640 4620 34649
rect 4672 34640 4674 34649
rect 4618 34575 4674 34584
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4620 33584 4672 33590
rect 4620 33526 4672 33532
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 3938 31878 4016 31906
rect 3882 31855 3938 31864
rect 3792 30252 3844 30258
rect 3792 30194 3844 30200
rect 3792 30048 3844 30054
rect 3792 29990 3844 29996
rect 3700 27464 3752 27470
rect 3700 27406 3752 27412
rect 3608 27328 3660 27334
rect 3608 27270 3660 27276
rect 3620 26382 3648 27270
rect 3608 26376 3660 26382
rect 3608 26318 3660 26324
rect 3516 25492 3568 25498
rect 3516 25434 3568 25440
rect 3712 25362 3740 27406
rect 3804 25838 3832 29990
rect 3896 29850 3924 31855
rect 4252 31680 4304 31686
rect 4252 31622 4304 31628
rect 4264 31414 4292 31622
rect 4252 31408 4304 31414
rect 4252 31350 4304 31356
rect 3976 31272 4028 31278
rect 3976 31214 4028 31220
rect 3988 30734 4016 31214
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 3976 30728 4028 30734
rect 3976 30670 4028 30676
rect 3988 30190 4016 30670
rect 4068 30252 4120 30258
rect 4068 30194 4120 30200
rect 3976 30184 4028 30190
rect 3976 30126 4028 30132
rect 3884 29844 3936 29850
rect 3884 29786 3936 29792
rect 3884 29708 3936 29714
rect 3884 29650 3936 29656
rect 3896 27334 3924 29650
rect 3976 29572 4028 29578
rect 3976 29514 4028 29520
rect 3884 27328 3936 27334
rect 3884 27270 3936 27276
rect 3896 27130 3924 27270
rect 3884 27124 3936 27130
rect 3884 27066 3936 27072
rect 3884 26444 3936 26450
rect 3884 26386 3936 26392
rect 3792 25832 3844 25838
rect 3792 25774 3844 25780
rect 3700 25356 3752 25362
rect 3700 25298 3752 25304
rect 3698 24984 3754 24993
rect 3698 24919 3754 24928
rect 3712 24818 3740 24919
rect 3700 24812 3752 24818
rect 3700 24754 3752 24760
rect 3896 22778 3924 26386
rect 3988 25498 4016 29514
rect 4080 28966 4108 30194
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4632 29730 4660 33526
rect 4724 30802 4752 35498
rect 5092 34202 5120 37284
rect 6552 37266 6604 37272
rect 6000 37120 6052 37126
rect 5920 37080 6000 37108
rect 5920 36922 5948 37080
rect 6000 37062 6052 37068
rect 5908 36916 5960 36922
rect 5908 36858 5960 36864
rect 6276 36848 6328 36854
rect 6276 36790 6328 36796
rect 6288 36582 6316 36790
rect 6368 36712 6420 36718
rect 6368 36654 6420 36660
rect 6276 36576 6328 36582
rect 6276 36518 6328 36524
rect 5722 35864 5778 35873
rect 5722 35799 5778 35808
rect 5736 35766 5764 35799
rect 5264 35760 5316 35766
rect 5262 35728 5264 35737
rect 5724 35760 5776 35766
rect 5316 35728 5318 35737
rect 5724 35702 5776 35708
rect 5262 35663 5318 35672
rect 5172 35012 5224 35018
rect 5172 34954 5224 34960
rect 5080 34196 5132 34202
rect 5080 34138 5132 34144
rect 4804 33992 4856 33998
rect 4804 33934 4856 33940
rect 4988 33992 5040 33998
rect 4988 33934 5040 33940
rect 4816 31754 4844 33934
rect 5000 32910 5028 33934
rect 5184 33153 5212 34954
rect 5632 34944 5684 34950
rect 5632 34886 5684 34892
rect 5540 34604 5592 34610
rect 5540 34546 5592 34552
rect 5264 34400 5316 34406
rect 5264 34342 5316 34348
rect 5448 34400 5500 34406
rect 5448 34342 5500 34348
rect 5276 34202 5304 34342
rect 5264 34196 5316 34202
rect 5264 34138 5316 34144
rect 5460 33998 5488 34342
rect 5552 34066 5580 34546
rect 5540 34060 5592 34066
rect 5540 34002 5592 34008
rect 5448 33992 5500 33998
rect 5448 33934 5500 33940
rect 5552 33522 5580 34002
rect 5644 33998 5672 34886
rect 5816 34604 5868 34610
rect 5816 34546 5868 34552
rect 5632 33992 5684 33998
rect 5632 33934 5684 33940
rect 5632 33856 5684 33862
rect 5632 33798 5684 33804
rect 5540 33516 5592 33522
rect 5540 33458 5592 33464
rect 5170 33144 5226 33153
rect 5170 33079 5226 33088
rect 5552 33046 5580 33458
rect 5540 33040 5592 33046
rect 5540 32982 5592 32988
rect 5448 32972 5500 32978
rect 5448 32914 5500 32920
rect 4988 32904 5040 32910
rect 5040 32852 5212 32858
rect 4988 32846 5212 32852
rect 5000 32830 5212 32846
rect 5080 32564 5132 32570
rect 5080 32506 5132 32512
rect 4816 31726 5028 31754
rect 4804 30932 4856 30938
rect 4804 30874 4856 30880
rect 4712 30796 4764 30802
rect 4712 30738 4764 30744
rect 4816 29850 4844 30874
rect 4896 30796 4948 30802
rect 4896 30738 4948 30744
rect 4804 29844 4856 29850
rect 4804 29786 4856 29792
rect 4632 29702 4844 29730
rect 4712 29572 4764 29578
rect 4712 29514 4764 29520
rect 4068 28960 4120 28966
rect 4068 28902 4120 28908
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4160 28620 4212 28626
rect 4160 28562 4212 28568
rect 4068 28484 4120 28490
rect 4068 28426 4120 28432
rect 4080 28218 4108 28426
rect 4068 28212 4120 28218
rect 4068 28154 4120 28160
rect 4068 28076 4120 28082
rect 4172 28064 4200 28562
rect 4620 28416 4672 28422
rect 4620 28358 4672 28364
rect 4120 28036 4200 28064
rect 4526 28112 4582 28121
rect 4526 28047 4528 28056
rect 4068 28018 4120 28024
rect 4580 28047 4582 28056
rect 4528 28018 4580 28024
rect 4080 27554 4108 28018
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4632 27606 4660 28358
rect 4620 27600 4672 27606
rect 4080 27526 4200 27554
rect 4620 27542 4672 27548
rect 4172 27418 4200 27526
rect 4172 27390 4660 27418
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4528 26376 4580 26382
rect 4066 26344 4122 26353
rect 4528 26318 4580 26324
rect 4066 26279 4122 26288
rect 4080 26042 4108 26279
rect 4068 26036 4120 26042
rect 4068 25978 4120 25984
rect 4540 25945 4568 26318
rect 4526 25936 4582 25945
rect 4068 25900 4120 25906
rect 4632 25906 4660 27390
rect 4724 25974 4752 29514
rect 4816 26314 4844 29702
rect 4908 27334 4936 30738
rect 5000 28150 5028 31726
rect 5092 28966 5120 32506
rect 5184 31142 5212 32830
rect 5460 32298 5488 32914
rect 5552 32570 5580 32982
rect 5644 32842 5672 33798
rect 5632 32836 5684 32842
rect 5632 32778 5684 32784
rect 5540 32564 5592 32570
rect 5540 32506 5592 32512
rect 5448 32292 5500 32298
rect 5368 32252 5448 32280
rect 5368 31754 5396 32252
rect 5448 32234 5500 32240
rect 5552 31890 5580 32506
rect 5540 31884 5592 31890
rect 5540 31826 5592 31832
rect 5448 31816 5500 31822
rect 5448 31758 5500 31764
rect 5276 31726 5396 31754
rect 5172 31136 5224 31142
rect 5172 31078 5224 31084
rect 5276 30938 5304 31726
rect 5460 31346 5488 31758
rect 5632 31748 5684 31754
rect 5632 31690 5684 31696
rect 5448 31340 5500 31346
rect 5368 31300 5448 31328
rect 5264 30932 5316 30938
rect 5264 30874 5316 30880
rect 5264 30660 5316 30666
rect 5184 30620 5264 30648
rect 5080 28960 5132 28966
rect 5080 28902 5132 28908
rect 5078 28520 5134 28529
rect 5078 28455 5080 28464
rect 5132 28455 5134 28464
rect 5080 28426 5132 28432
rect 5078 28384 5134 28393
rect 5078 28319 5134 28328
rect 4988 28144 5040 28150
rect 4988 28086 5040 28092
rect 4896 27328 4948 27334
rect 4896 27270 4948 27276
rect 5092 27112 5120 28319
rect 5000 27084 5120 27112
rect 4896 27056 4948 27062
rect 4894 27024 4896 27033
rect 4948 27024 4950 27033
rect 4894 26959 4950 26968
rect 4896 26784 4948 26790
rect 4896 26726 4948 26732
rect 4908 26382 4936 26726
rect 4896 26376 4948 26382
rect 4896 26318 4948 26324
rect 4804 26308 4856 26314
rect 4804 26250 4856 26256
rect 4802 26208 4858 26217
rect 4802 26143 4858 26152
rect 4712 25968 4764 25974
rect 4712 25910 4764 25916
rect 4526 25871 4582 25880
rect 4620 25900 4672 25906
rect 4068 25842 4120 25848
rect 4620 25842 4672 25848
rect 3976 25492 4028 25498
rect 3976 25434 4028 25440
rect 3976 24812 4028 24818
rect 3976 24754 4028 24760
rect 3988 24410 4016 24754
rect 3976 24404 4028 24410
rect 3976 24346 4028 24352
rect 4080 23866 4108 25842
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4618 25528 4674 25537
rect 4618 25463 4674 25472
rect 4160 25288 4212 25294
rect 4160 25230 4212 25236
rect 4172 24614 4200 25230
rect 4632 24750 4660 25463
rect 4816 25294 4844 26143
rect 4804 25288 4856 25294
rect 4804 25230 4856 25236
rect 4908 25106 4936 26318
rect 5000 26042 5028 27084
rect 5080 26988 5132 26994
rect 5080 26930 5132 26936
rect 5092 26586 5120 26930
rect 5080 26580 5132 26586
rect 5080 26522 5132 26528
rect 5078 26480 5134 26489
rect 5078 26415 5134 26424
rect 5092 26246 5120 26415
rect 5080 26240 5132 26246
rect 5080 26182 5132 26188
rect 4988 26036 5040 26042
rect 4988 25978 5040 25984
rect 5000 25226 5028 25978
rect 5080 25900 5132 25906
rect 5080 25842 5132 25848
rect 4988 25220 5040 25226
rect 4988 25162 5040 25168
rect 4816 25078 4936 25106
rect 4712 24812 4764 24818
rect 4712 24754 4764 24760
rect 4620 24744 4672 24750
rect 4620 24686 4672 24692
rect 4160 24608 4212 24614
rect 4160 24550 4212 24556
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4068 23860 4120 23866
rect 4068 23802 4120 23808
rect 3516 22772 3568 22778
rect 3516 22714 3568 22720
rect 3884 22772 3936 22778
rect 3884 22714 3936 22720
rect 3424 22636 3476 22642
rect 3424 22578 3476 22584
rect 2964 22432 3016 22438
rect 2964 22374 3016 22380
rect 2976 21894 3004 22374
rect 3528 22030 3556 22714
rect 3516 22024 3568 22030
rect 3516 21966 3568 21972
rect 2964 21888 3016 21894
rect 2964 21830 3016 21836
rect 2780 21684 2832 21690
rect 2780 21626 2832 21632
rect 2872 21684 2924 21690
rect 2872 21626 2924 21632
rect 2872 21140 2924 21146
rect 2872 21082 2924 21088
rect 2688 21072 2740 21078
rect 2688 21014 2740 21020
rect 2780 20528 2832 20534
rect 2780 20470 2832 20476
rect 2792 19938 2820 20470
rect 2884 20058 2912 21082
rect 2976 20602 3004 21830
rect 2964 20596 3016 20602
rect 2964 20538 3016 20544
rect 3896 20534 3924 22714
rect 4080 22098 4108 23802
rect 4620 23588 4672 23594
rect 4620 23530 4672 23536
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4632 23322 4660 23530
rect 4620 23316 4672 23322
rect 4620 23258 4672 23264
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4068 22092 4120 22098
rect 4068 22034 4120 22040
rect 4620 21344 4672 21350
rect 4620 21286 4672 21292
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4632 21146 4660 21286
rect 4620 21140 4672 21146
rect 4620 21082 4672 21088
rect 4068 20596 4120 20602
rect 4068 20538 4120 20544
rect 3884 20528 3936 20534
rect 3884 20470 3936 20476
rect 3330 20088 3386 20097
rect 2872 20052 2924 20058
rect 2872 19994 2924 20000
rect 3148 20052 3200 20058
rect 4080 20058 4108 20538
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 3330 20023 3332 20032
rect 3148 19994 3200 20000
rect 3384 20023 3386 20032
rect 4068 20052 4120 20058
rect 3332 19994 3384 20000
rect 4068 19994 4120 20000
rect 2792 19910 2912 19938
rect 2320 19304 2372 19310
rect 2320 19246 2372 19252
rect 2226 19000 2282 19009
rect 2226 18935 2228 18944
rect 2280 18935 2282 18944
rect 2228 18906 2280 18912
rect 2780 18624 2832 18630
rect 2780 18566 2832 18572
rect 2792 16114 2820 18566
rect 2780 16108 2832 16114
rect 2780 16050 2832 16056
rect 1952 14272 2004 14278
rect 1952 14214 2004 14220
rect 1768 5364 1820 5370
rect 1768 5306 1820 5312
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1596 4865 1624 5170
rect 1582 4856 1638 4865
rect 1582 4791 1584 4800
rect 1636 4791 1638 4800
rect 1584 4762 1636 4768
rect 1676 3936 1728 3942
rect 1676 3878 1728 3884
rect 1688 3534 1716 3878
rect 1676 3528 1728 3534
rect 1674 3496 1676 3505
rect 1728 3496 1730 3505
rect 1674 3431 1730 3440
rect 1964 3058 1992 14214
rect 2412 13864 2464 13870
rect 2412 13806 2464 13812
rect 2424 10674 2452 13806
rect 2412 10668 2464 10674
rect 2412 10610 2464 10616
rect 2884 3670 2912 19910
rect 3160 6914 3188 19994
rect 3344 19786 3372 19994
rect 3332 19780 3384 19786
rect 3332 19722 3384 19728
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4724 14006 4752 24754
rect 4816 24070 4844 25078
rect 4804 24064 4856 24070
rect 4804 24006 4856 24012
rect 4816 14618 4844 24006
rect 4988 23860 5040 23866
rect 4988 23802 5040 23808
rect 4896 22024 4948 22030
rect 4896 21966 4948 21972
rect 4908 20806 4936 21966
rect 5000 21690 5028 23802
rect 5092 22098 5120 25842
rect 5184 25770 5212 30620
rect 5264 30602 5316 30608
rect 5264 30320 5316 30326
rect 5264 30262 5316 30268
rect 5172 25764 5224 25770
rect 5172 25706 5224 25712
rect 5276 25498 5304 30262
rect 5368 26489 5396 31300
rect 5448 31282 5500 31288
rect 5448 31136 5500 31142
rect 5448 31078 5500 31084
rect 5460 28393 5488 31078
rect 5538 30968 5594 30977
rect 5538 30903 5594 30912
rect 5552 29510 5580 30903
rect 5644 30802 5672 31690
rect 5632 30796 5684 30802
rect 5632 30738 5684 30744
rect 5644 30598 5672 30738
rect 5632 30592 5684 30598
rect 5632 30534 5684 30540
rect 5828 29714 5856 34546
rect 5908 33584 5960 33590
rect 5908 33526 5960 33532
rect 5920 31668 5948 33526
rect 6000 32768 6052 32774
rect 6380 32745 6408 36654
rect 6460 35488 6512 35494
rect 6460 35430 6512 35436
rect 6000 32710 6052 32716
rect 6366 32736 6422 32745
rect 6012 31822 6040 32710
rect 6366 32671 6422 32680
rect 6274 32056 6330 32065
rect 6274 31991 6330 32000
rect 6000 31816 6052 31822
rect 6000 31758 6052 31764
rect 6092 31680 6144 31686
rect 5920 31640 6092 31668
rect 5920 30734 5948 31640
rect 6092 31622 6144 31628
rect 6000 31272 6052 31278
rect 6000 31214 6052 31220
rect 5908 30728 5960 30734
rect 5908 30670 5960 30676
rect 6012 30326 6040 31214
rect 6184 30728 6236 30734
rect 6184 30670 6236 30676
rect 6000 30320 6052 30326
rect 6000 30262 6052 30268
rect 5908 30184 5960 30190
rect 5908 30126 5960 30132
rect 5816 29708 5868 29714
rect 5816 29650 5868 29656
rect 5920 29646 5948 30126
rect 5908 29640 5960 29646
rect 5908 29582 5960 29588
rect 5540 29504 5592 29510
rect 5540 29446 5592 29452
rect 5540 29164 5592 29170
rect 5540 29106 5592 29112
rect 5446 28384 5502 28393
rect 5446 28319 5502 28328
rect 5552 28234 5580 29106
rect 5920 29102 5948 29582
rect 5908 29096 5960 29102
rect 5908 29038 5960 29044
rect 5632 28960 5684 28966
rect 5632 28902 5684 28908
rect 5816 28960 5868 28966
rect 5816 28902 5868 28908
rect 5460 28206 5580 28234
rect 5460 28082 5488 28206
rect 5540 28144 5592 28150
rect 5540 28086 5592 28092
rect 5448 28076 5500 28082
rect 5448 28018 5500 28024
rect 5460 27282 5488 28018
rect 5552 27470 5580 28086
rect 5540 27464 5592 27470
rect 5540 27406 5592 27412
rect 5460 27254 5580 27282
rect 5448 27124 5500 27130
rect 5448 27066 5500 27072
rect 5354 26480 5410 26489
rect 5354 26415 5410 26424
rect 5460 26194 5488 27066
rect 5368 26166 5488 26194
rect 5264 25492 5316 25498
rect 5264 25434 5316 25440
rect 5172 25220 5224 25226
rect 5172 25162 5224 25168
rect 5184 23746 5212 25162
rect 5368 24698 5396 26166
rect 5446 26072 5502 26081
rect 5446 26007 5502 26016
rect 5276 24670 5396 24698
rect 5276 23866 5304 24670
rect 5356 24608 5408 24614
rect 5354 24576 5356 24585
rect 5408 24576 5410 24585
rect 5354 24511 5410 24520
rect 5264 23860 5316 23866
rect 5264 23802 5316 23808
rect 5184 23718 5304 23746
rect 5172 22772 5224 22778
rect 5172 22714 5224 22720
rect 5080 22092 5132 22098
rect 5080 22034 5132 22040
rect 4988 21684 5040 21690
rect 4988 21626 5040 21632
rect 4896 20800 4948 20806
rect 4896 20742 4948 20748
rect 4908 20534 4936 20742
rect 4896 20528 4948 20534
rect 4896 20470 4948 20476
rect 5184 18970 5212 22714
rect 5276 22710 5304 23718
rect 5460 22778 5488 26007
rect 5552 23322 5580 27254
rect 5644 26382 5672 28902
rect 5724 28416 5776 28422
rect 5724 28358 5776 28364
rect 5736 28014 5764 28358
rect 5724 28008 5776 28014
rect 5724 27950 5776 27956
rect 5828 27826 5856 28902
rect 5920 27878 5948 29038
rect 5736 27798 5856 27826
rect 5908 27872 5960 27878
rect 5908 27814 5960 27820
rect 5632 26376 5684 26382
rect 5632 26318 5684 26324
rect 5736 25906 5764 27798
rect 5814 27432 5870 27441
rect 5814 27367 5870 27376
rect 5828 27010 5856 27367
rect 6012 27282 6040 30262
rect 6092 29164 6144 29170
rect 6092 29106 6144 29112
rect 6104 27402 6132 29106
rect 6196 28626 6224 30670
rect 6288 29102 6316 31991
rect 6368 29572 6420 29578
rect 6368 29514 6420 29520
rect 6276 29096 6328 29102
rect 6276 29038 6328 29044
rect 6276 28960 6328 28966
rect 6276 28902 6328 28908
rect 6184 28620 6236 28626
rect 6184 28562 6236 28568
rect 6288 28422 6316 28902
rect 6276 28416 6328 28422
rect 6276 28358 6328 28364
rect 6184 28008 6236 28014
rect 6182 27976 6184 27985
rect 6236 27976 6238 27985
rect 6182 27911 6238 27920
rect 6092 27396 6144 27402
rect 6092 27338 6144 27344
rect 6012 27254 6132 27282
rect 5828 27000 5864 27010
rect 5824 26994 5876 27000
rect 5824 26936 5876 26942
rect 5836 26874 5864 26936
rect 5828 26846 5864 26874
rect 5724 25900 5776 25906
rect 5724 25842 5776 25848
rect 5632 25832 5684 25838
rect 5632 25774 5684 25780
rect 5644 25362 5672 25774
rect 5632 25356 5684 25362
rect 5632 25298 5684 25304
rect 5632 25152 5684 25158
rect 5828 25129 5856 26846
rect 6000 25356 6052 25362
rect 6000 25298 6052 25304
rect 5632 25094 5684 25100
rect 5814 25120 5870 25129
rect 5644 24818 5672 25094
rect 5814 25055 5870 25064
rect 5632 24812 5684 24818
rect 5632 24754 5684 24760
rect 5828 24410 5856 25055
rect 6012 24818 6040 25298
rect 6000 24812 6052 24818
rect 6000 24754 6052 24760
rect 5816 24404 5868 24410
rect 5816 24346 5868 24352
rect 5722 23352 5778 23361
rect 5540 23316 5592 23322
rect 5722 23287 5724 23296
rect 5540 23258 5592 23264
rect 5776 23287 5778 23296
rect 5724 23258 5776 23264
rect 5552 22778 5580 23258
rect 5448 22772 5500 22778
rect 5448 22714 5500 22720
rect 5540 22772 5592 22778
rect 5540 22714 5592 22720
rect 5264 22704 5316 22710
rect 5264 22646 5316 22652
rect 5264 22228 5316 22234
rect 5264 22170 5316 22176
rect 5276 21146 5304 22170
rect 5736 21554 5764 23258
rect 6000 22568 6052 22574
rect 6000 22510 6052 22516
rect 6012 22234 6040 22510
rect 6000 22228 6052 22234
rect 6000 22170 6052 22176
rect 6104 22094 6132 27254
rect 6184 27124 6236 27130
rect 6184 27066 6236 27072
rect 6196 26790 6224 27066
rect 6184 26784 6236 26790
rect 6184 26726 6236 26732
rect 6184 25968 6236 25974
rect 6184 25910 6236 25916
rect 6196 25498 6224 25910
rect 6276 25696 6328 25702
rect 6276 25638 6328 25644
rect 6184 25492 6236 25498
rect 6184 25434 6236 25440
rect 6104 22066 6224 22094
rect 6196 21690 6224 22066
rect 6184 21684 6236 21690
rect 6184 21626 6236 21632
rect 5724 21548 5776 21554
rect 5724 21490 5776 21496
rect 5264 21140 5316 21146
rect 5264 21082 5316 21088
rect 5276 20602 5304 21082
rect 5264 20596 5316 20602
rect 5264 20538 5316 20544
rect 6196 19718 6224 21626
rect 6288 20534 6316 25638
rect 6380 25226 6408 29514
rect 6472 27470 6500 35430
rect 6564 34950 6592 37266
rect 6828 36712 6880 36718
rect 6828 36654 6880 36660
rect 7196 36712 7248 36718
rect 7196 36654 7248 36660
rect 6840 36242 6868 36654
rect 7102 36544 7158 36553
rect 7102 36479 7158 36488
rect 6828 36236 6880 36242
rect 6828 36178 6880 36184
rect 6920 36032 6972 36038
rect 6920 35974 6972 35980
rect 6552 34944 6604 34950
rect 6552 34886 6604 34892
rect 6564 32473 6592 34886
rect 6932 34626 6960 35974
rect 7116 35698 7144 36479
rect 7208 36378 7236 36654
rect 7196 36372 7248 36378
rect 7196 36314 7248 36320
rect 7196 36100 7248 36106
rect 7196 36042 7248 36048
rect 7104 35692 7156 35698
rect 7104 35634 7156 35640
rect 7208 35494 7236 36042
rect 7196 35488 7248 35494
rect 7196 35430 7248 35436
rect 7208 35290 7236 35430
rect 7196 35284 7248 35290
rect 7196 35226 7248 35232
rect 7392 35193 7420 39222
rect 8390 39200 8446 39800
rect 10322 39200 10378 39800
rect 12254 39200 12310 39800
rect 13542 39200 13598 39800
rect 15474 39200 15530 39800
rect 15580 39222 15792 39250
rect 8208 37460 8260 37466
rect 8208 37402 8260 37408
rect 8220 37262 8248 37402
rect 8208 37256 8260 37262
rect 8208 37198 8260 37204
rect 8116 36712 8168 36718
rect 8116 36654 8168 36660
rect 7748 36236 7800 36242
rect 7748 36178 7800 36184
rect 7654 35320 7710 35329
rect 7654 35255 7656 35264
rect 7708 35255 7710 35264
rect 7656 35226 7708 35232
rect 7378 35184 7434 35193
rect 7378 35119 7434 35128
rect 7196 34672 7248 34678
rect 6932 34598 7052 34626
rect 7196 34614 7248 34620
rect 6920 34536 6972 34542
rect 6920 34478 6972 34484
rect 6644 32836 6696 32842
rect 6644 32778 6696 32784
rect 6550 32464 6606 32473
rect 6550 32399 6606 32408
rect 6656 31770 6684 32778
rect 6734 31784 6790 31793
rect 6656 31742 6734 31770
rect 6734 31719 6790 31728
rect 6644 28484 6696 28490
rect 6644 28426 6696 28432
rect 6656 28082 6684 28426
rect 6644 28076 6696 28082
rect 6644 28018 6696 28024
rect 6552 27872 6604 27878
rect 6552 27814 6604 27820
rect 6460 27464 6512 27470
rect 6460 27406 6512 27412
rect 6460 27328 6512 27334
rect 6460 27270 6512 27276
rect 6472 27169 6500 27270
rect 6458 27160 6514 27169
rect 6458 27095 6514 27104
rect 6460 26308 6512 26314
rect 6460 26250 6512 26256
rect 6368 25220 6420 25226
rect 6368 25162 6420 25168
rect 6472 21622 6500 26250
rect 6564 22574 6592 27814
rect 6644 26376 6696 26382
rect 6642 26344 6644 26353
rect 6696 26344 6698 26353
rect 6642 26279 6698 26288
rect 6748 25906 6776 31719
rect 6932 30666 6960 34478
rect 7024 34406 7052 34598
rect 7012 34400 7064 34406
rect 7012 34342 7064 34348
rect 7024 33930 7052 34342
rect 7012 33924 7064 33930
rect 7012 33866 7064 33872
rect 7012 33108 7064 33114
rect 7012 33050 7064 33056
rect 7024 32570 7052 33050
rect 7104 33040 7156 33046
rect 7104 32982 7156 32988
rect 7012 32564 7064 32570
rect 7012 32506 7064 32512
rect 6920 30660 6972 30666
rect 6920 30602 6972 30608
rect 6920 29504 6972 29510
rect 6920 29446 6972 29452
rect 6932 29102 6960 29446
rect 6920 29096 6972 29102
rect 6920 29038 6972 29044
rect 6932 28762 6960 29038
rect 6920 28756 6972 28762
rect 6920 28698 6972 28704
rect 6826 28520 6882 28529
rect 6826 28455 6882 28464
rect 6736 25900 6788 25906
rect 6736 25842 6788 25848
rect 6840 23322 6868 28455
rect 6920 28076 6972 28082
rect 6920 28018 6972 28024
rect 6932 27402 6960 28018
rect 6920 27396 6972 27402
rect 6920 27338 6972 27344
rect 7024 26586 7052 32506
rect 7116 32298 7144 32982
rect 7104 32292 7156 32298
rect 7104 32234 7156 32240
rect 7104 32020 7156 32026
rect 7104 31962 7156 31968
rect 7116 29646 7144 31962
rect 7208 31754 7236 34614
rect 7288 34536 7340 34542
rect 7288 34478 7340 34484
rect 7300 33590 7328 34478
rect 7564 34400 7616 34406
rect 7564 34342 7616 34348
rect 7472 33992 7524 33998
rect 7472 33934 7524 33940
rect 7288 33584 7340 33590
rect 7288 33526 7340 33532
rect 7286 33144 7342 33153
rect 7286 33079 7288 33088
rect 7340 33079 7342 33088
rect 7288 33050 7340 33056
rect 7484 32994 7512 33934
rect 7288 32972 7340 32978
rect 7288 32914 7340 32920
rect 7392 32966 7512 32994
rect 7300 32609 7328 32914
rect 7286 32600 7342 32609
rect 7286 32535 7342 32544
rect 7288 32020 7340 32026
rect 7288 31962 7340 31968
rect 7300 31929 7328 31962
rect 7286 31920 7342 31929
rect 7286 31855 7342 31864
rect 7196 31748 7248 31754
rect 7196 31690 7248 31696
rect 7104 29640 7156 29646
rect 7104 29582 7156 29588
rect 7208 29492 7236 31690
rect 7288 30388 7340 30394
rect 7288 30330 7340 30336
rect 7116 29464 7236 29492
rect 7116 27470 7144 29464
rect 7104 27464 7156 27470
rect 7104 27406 7156 27412
rect 7012 26580 7064 26586
rect 7012 26522 7064 26528
rect 7012 26376 7064 26382
rect 7012 26318 7064 26324
rect 7024 24750 7052 26318
rect 7012 24744 7064 24750
rect 7012 24686 7064 24692
rect 7116 23730 7144 27406
rect 7300 26382 7328 30330
rect 7392 27470 7420 32966
rect 7472 32904 7524 32910
rect 7472 32846 7524 32852
rect 7484 31346 7512 32846
rect 7576 31958 7604 34342
rect 7656 34196 7708 34202
rect 7656 34138 7708 34144
rect 7564 31952 7616 31958
rect 7564 31894 7616 31900
rect 7472 31340 7524 31346
rect 7472 31282 7524 31288
rect 7668 30938 7696 34138
rect 7760 33998 7788 36178
rect 7840 35284 7892 35290
rect 7840 35226 7892 35232
rect 7852 35018 7880 35226
rect 7840 35012 7892 35018
rect 7840 34954 7892 34960
rect 7932 34468 7984 34474
rect 7932 34410 7984 34416
rect 7840 34400 7892 34406
rect 7840 34342 7892 34348
rect 7852 34202 7880 34342
rect 7840 34196 7892 34202
rect 7840 34138 7892 34144
rect 7944 33998 7972 34410
rect 7748 33992 7800 33998
rect 7748 33934 7800 33940
rect 7932 33992 7984 33998
rect 7932 33934 7984 33940
rect 7932 33856 7984 33862
rect 7932 33798 7984 33804
rect 7944 33590 7972 33798
rect 7932 33584 7984 33590
rect 7932 33526 7984 33532
rect 7840 33312 7892 33318
rect 7840 33254 7892 33260
rect 7932 33312 7984 33318
rect 7932 33254 7984 33260
rect 7748 32768 7800 32774
rect 7748 32710 7800 32716
rect 7760 32502 7788 32710
rect 7748 32496 7800 32502
rect 7748 32438 7800 32444
rect 7748 31204 7800 31210
rect 7748 31146 7800 31152
rect 7656 30932 7708 30938
rect 7656 30874 7708 30880
rect 7668 30394 7696 30874
rect 7656 30388 7708 30394
rect 7656 30330 7708 30336
rect 7760 30190 7788 31146
rect 7748 30184 7800 30190
rect 7748 30126 7800 30132
rect 7472 30048 7524 30054
rect 7472 29990 7524 29996
rect 7484 28082 7512 29990
rect 7760 29850 7788 30126
rect 7748 29844 7800 29850
rect 7748 29786 7800 29792
rect 7656 28960 7708 28966
rect 7656 28902 7708 28908
rect 7748 28960 7800 28966
rect 7748 28902 7800 28908
rect 7564 28756 7616 28762
rect 7564 28698 7616 28704
rect 7576 28558 7604 28698
rect 7564 28552 7616 28558
rect 7564 28494 7616 28500
rect 7472 28076 7524 28082
rect 7472 28018 7524 28024
rect 7668 28014 7696 28902
rect 7760 28626 7788 28902
rect 7748 28620 7800 28626
rect 7748 28562 7800 28568
rect 7748 28416 7800 28422
rect 7748 28358 7800 28364
rect 7656 28008 7708 28014
rect 7656 27950 7708 27956
rect 7564 27940 7616 27946
rect 7564 27882 7616 27888
rect 7576 27577 7604 27882
rect 7562 27568 7618 27577
rect 7562 27503 7618 27512
rect 7380 27464 7432 27470
rect 7380 27406 7432 27412
rect 7564 27328 7616 27334
rect 7562 27296 7564 27305
rect 7616 27296 7618 27305
rect 7562 27231 7618 27240
rect 7380 26988 7432 26994
rect 7380 26930 7432 26936
rect 7392 26586 7420 26930
rect 7668 26586 7696 27950
rect 7380 26580 7432 26586
rect 7380 26522 7432 26528
rect 7564 26580 7616 26586
rect 7564 26522 7616 26528
rect 7656 26580 7708 26586
rect 7656 26522 7708 26528
rect 7288 26376 7340 26382
rect 7288 26318 7340 26324
rect 7378 26208 7434 26217
rect 7378 26143 7434 26152
rect 7286 25936 7342 25945
rect 7286 25871 7342 25880
rect 7300 25294 7328 25871
rect 7392 25401 7420 26143
rect 7576 25838 7604 26522
rect 7656 26308 7708 26314
rect 7656 26250 7708 26256
rect 7564 25832 7616 25838
rect 7564 25774 7616 25780
rect 7378 25392 7434 25401
rect 7378 25327 7434 25336
rect 7288 25288 7340 25294
rect 7288 25230 7340 25236
rect 7196 24064 7248 24070
rect 7196 24006 7248 24012
rect 7208 23798 7236 24006
rect 7196 23792 7248 23798
rect 7196 23734 7248 23740
rect 7104 23724 7156 23730
rect 7104 23666 7156 23672
rect 7194 23624 7250 23633
rect 7194 23559 7196 23568
rect 7248 23559 7250 23568
rect 7196 23530 7248 23536
rect 6828 23316 6880 23322
rect 6828 23258 6880 23264
rect 6552 22568 6604 22574
rect 6552 22510 6604 22516
rect 6564 21690 6592 22510
rect 7392 22098 7420 25327
rect 7380 22092 7432 22098
rect 7380 22034 7432 22040
rect 6552 21684 6604 21690
rect 6552 21626 6604 21632
rect 6460 21616 6512 21622
rect 6460 21558 6512 21564
rect 6276 20528 6328 20534
rect 6276 20470 6328 20476
rect 6184 19712 6236 19718
rect 6184 19654 6236 19660
rect 5172 18964 5224 18970
rect 5172 18906 5224 18912
rect 7576 17202 7604 25774
rect 7668 24188 7696 26250
rect 7760 24290 7788 28358
rect 7852 27441 7880 33254
rect 7944 30054 7972 33254
rect 8128 31754 8156 36654
rect 8208 36168 8260 36174
rect 8206 36136 8208 36145
rect 8260 36136 8262 36145
rect 8206 36071 8262 36080
rect 8404 35834 8432 39200
rect 9128 37256 9180 37262
rect 9128 37198 9180 37204
rect 9140 36718 9168 37198
rect 9588 37188 9640 37194
rect 9588 37130 9640 37136
rect 9036 36712 9088 36718
rect 9036 36654 9088 36660
rect 9128 36712 9180 36718
rect 9128 36654 9180 36660
rect 9048 36281 9076 36654
rect 9034 36272 9090 36281
rect 9034 36207 9090 36216
rect 8576 36168 8628 36174
rect 8576 36110 8628 36116
rect 8392 35828 8444 35834
rect 8392 35770 8444 35776
rect 8300 35556 8352 35562
rect 8300 35498 8352 35504
rect 8312 35465 8340 35498
rect 8298 35456 8354 35465
rect 8298 35391 8354 35400
rect 8588 35086 8616 36110
rect 8852 35760 8904 35766
rect 8852 35702 8904 35708
rect 8576 35080 8628 35086
rect 8576 35022 8628 35028
rect 8208 34944 8260 34950
rect 8484 34944 8536 34950
rect 8260 34904 8340 34932
rect 8208 34886 8260 34892
rect 8206 34776 8262 34785
rect 8206 34711 8208 34720
rect 8260 34711 8262 34720
rect 8208 34682 8260 34688
rect 8208 34536 8260 34542
rect 8208 34478 8260 34484
rect 8220 32065 8248 34478
rect 8312 34202 8340 34904
rect 8484 34886 8536 34892
rect 8300 34196 8352 34202
rect 8300 34138 8352 34144
rect 8300 33992 8352 33998
rect 8300 33934 8352 33940
rect 8312 32910 8340 33934
rect 8496 33402 8524 34886
rect 8588 34406 8616 35022
rect 8668 35012 8720 35018
rect 8668 34954 8720 34960
rect 8576 34400 8628 34406
rect 8576 34342 8628 34348
rect 8496 33374 8616 33402
rect 8300 32904 8352 32910
rect 8300 32846 8352 32852
rect 8484 32768 8536 32774
rect 8484 32710 8536 32716
rect 8392 32360 8444 32366
rect 8392 32302 8444 32308
rect 8206 32056 8262 32065
rect 8206 31991 8262 32000
rect 8036 31726 8156 31754
rect 8036 30190 8064 31726
rect 8300 31476 8352 31482
rect 8300 31418 8352 31424
rect 8312 30326 8340 31418
rect 8300 30320 8352 30326
rect 8300 30262 8352 30268
rect 8024 30184 8076 30190
rect 8024 30126 8076 30132
rect 7932 30048 7984 30054
rect 7932 29990 7984 29996
rect 8404 29850 8432 32302
rect 8496 31414 8524 32710
rect 8588 31686 8616 33374
rect 8576 31680 8628 31686
rect 8576 31622 8628 31628
rect 8484 31408 8536 31414
rect 8484 31350 8536 31356
rect 8576 30660 8628 30666
rect 8496 30620 8576 30648
rect 8024 29844 8076 29850
rect 8024 29786 8076 29792
rect 8392 29844 8444 29850
rect 8392 29786 8444 29792
rect 7932 29232 7984 29238
rect 7932 29174 7984 29180
rect 7944 28490 7972 29174
rect 7932 28484 7984 28490
rect 7932 28426 7984 28432
rect 7838 27432 7894 27441
rect 7838 27367 7894 27376
rect 7840 27056 7892 27062
rect 7838 27024 7840 27033
rect 7892 27024 7894 27033
rect 8036 27010 8064 29786
rect 8404 29730 8432 29786
rect 8128 29702 8432 29730
rect 8128 29578 8156 29702
rect 8116 29572 8168 29578
rect 8116 29514 8168 29520
rect 8128 27674 8156 29514
rect 8298 29336 8354 29345
rect 8298 29271 8354 29280
rect 8208 29232 8260 29238
rect 8208 29174 8260 29180
rect 8220 29034 8248 29174
rect 8208 29028 8260 29034
rect 8208 28970 8260 28976
rect 8116 27668 8168 27674
rect 8116 27610 8168 27616
rect 8312 27418 8340 29271
rect 8392 29232 8444 29238
rect 8392 29174 8444 29180
rect 8404 28490 8432 29174
rect 8392 28484 8444 28490
rect 8392 28426 8444 28432
rect 8404 28014 8432 28426
rect 8392 28008 8444 28014
rect 8392 27950 8444 27956
rect 8220 27390 8340 27418
rect 8220 27130 8248 27390
rect 8300 27328 8352 27334
rect 8298 27296 8300 27305
rect 8352 27296 8354 27305
rect 8298 27231 8354 27240
rect 8208 27124 8260 27130
rect 8208 27066 8260 27072
rect 8036 26982 8156 27010
rect 7838 26959 7894 26968
rect 8024 26920 8076 26926
rect 8024 26862 8076 26868
rect 8036 26314 8064 26862
rect 7932 26308 7984 26314
rect 7932 26250 7984 26256
rect 8024 26308 8076 26314
rect 8024 26250 8076 26256
rect 7944 25498 7972 26250
rect 8128 26217 8156 26982
rect 8300 26308 8352 26314
rect 8300 26250 8352 26256
rect 8114 26208 8170 26217
rect 8114 26143 8170 26152
rect 8312 25838 8340 26250
rect 8300 25832 8352 25838
rect 8300 25774 8352 25780
rect 8208 25696 8260 25702
rect 8208 25638 8260 25644
rect 7932 25492 7984 25498
rect 7932 25434 7984 25440
rect 8024 25492 8076 25498
rect 8024 25434 8076 25440
rect 7944 24868 7972 25434
rect 8036 25158 8064 25434
rect 8024 25152 8076 25158
rect 8024 25094 8076 25100
rect 8024 24880 8076 24886
rect 7944 24840 8024 24868
rect 8024 24822 8076 24828
rect 7760 24262 7972 24290
rect 7748 24200 7800 24206
rect 7668 24168 7748 24188
rect 7840 24200 7892 24206
rect 7800 24168 7802 24177
rect 7668 24160 7746 24168
rect 7840 24142 7892 24148
rect 7746 24103 7802 24112
rect 7746 23760 7802 23769
rect 7746 23695 7748 23704
rect 7800 23695 7802 23704
rect 7748 23666 7800 23672
rect 7760 22778 7788 23666
rect 7852 23662 7880 24142
rect 7840 23656 7892 23662
rect 7840 23598 7892 23604
rect 7748 22772 7800 22778
rect 7748 22714 7800 22720
rect 7944 22506 7972 24262
rect 7932 22500 7984 22506
rect 7932 22442 7984 22448
rect 8220 22098 8248 25638
rect 8300 25152 8352 25158
rect 8300 25094 8352 25100
rect 8312 24818 8340 25094
rect 8300 24812 8352 24818
rect 8300 24754 8352 24760
rect 8300 24268 8352 24274
rect 8300 24210 8352 24216
rect 8312 24070 8340 24210
rect 8300 24064 8352 24070
rect 8300 24006 8352 24012
rect 8208 22092 8260 22098
rect 8208 22034 8260 22040
rect 7564 17196 7616 17202
rect 7564 17138 7616 17144
rect 6736 16992 6788 16998
rect 6736 16934 6788 16940
rect 4804 14612 4856 14618
rect 4804 14554 4856 14560
rect 4712 14000 4764 14006
rect 4712 13942 4764 13948
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 6748 12850 6776 16934
rect 6828 15360 6880 15366
rect 6828 15302 6880 15308
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 2976 6886 3188 6914
rect 2872 3664 2924 3670
rect 2872 3606 2924 3612
rect 1952 3052 2004 3058
rect 1952 2994 2004 3000
rect 2412 2984 2464 2990
rect 2412 2926 2464 2932
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 20 2576 72 2582
rect 20 2518 72 2524
rect 32 800 60 2518
rect 1308 2304 1360 2310
rect 1308 2246 1360 2252
rect 1320 800 1348 2246
rect 1688 1465 1716 2790
rect 2424 2446 2452 2926
rect 2976 2582 3004 6886
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4712 2916 4764 2922
rect 4712 2858 4764 2864
rect 4620 2848 4672 2854
rect 4620 2790 4672 2796
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 2964 2576 3016 2582
rect 4632 2530 4660 2790
rect 2964 2518 3016 2524
rect 4540 2502 4660 2530
rect 4724 2514 4752 2858
rect 4712 2508 4764 2514
rect 2412 2440 2464 2446
rect 2412 2382 2464 2388
rect 4540 2378 4568 2502
rect 4712 2450 4764 2456
rect 6840 2446 6868 15302
rect 8404 11150 8432 27950
rect 8496 25158 8524 30620
rect 8576 30602 8628 30608
rect 8680 29186 8708 34954
rect 8760 34944 8812 34950
rect 8760 34886 8812 34892
rect 8772 33930 8800 34886
rect 8864 34746 8892 35702
rect 8942 35320 8998 35329
rect 8942 35255 8998 35264
rect 8852 34740 8904 34746
rect 8852 34682 8904 34688
rect 8956 34649 8984 35255
rect 8942 34640 8998 34649
rect 8864 34598 8942 34626
rect 8760 33924 8812 33930
rect 8760 33866 8812 33872
rect 8864 32910 8892 34598
rect 8942 34575 8998 34584
rect 8944 34536 8996 34542
rect 8942 34504 8944 34513
rect 8996 34504 8998 34513
rect 8942 34439 8998 34448
rect 8852 32904 8904 32910
rect 8852 32846 8904 32852
rect 9048 32502 9076 36207
rect 9140 36174 9168 36654
rect 9128 36168 9180 36174
rect 9128 36110 9180 36116
rect 9140 35834 9168 36110
rect 9496 36100 9548 36106
rect 9496 36042 9548 36048
rect 9128 35828 9180 35834
rect 9128 35770 9180 35776
rect 9220 35828 9272 35834
rect 9220 35770 9272 35776
rect 9232 35630 9260 35770
rect 9220 35624 9272 35630
rect 9220 35566 9272 35572
rect 9404 35216 9456 35222
rect 9126 35184 9182 35193
rect 9404 35158 9456 35164
rect 9126 35119 9182 35128
rect 9140 35086 9168 35119
rect 9128 35080 9180 35086
rect 9128 35022 9180 35028
rect 9416 34542 9444 35158
rect 9508 35018 9536 36042
rect 9496 35012 9548 35018
rect 9496 34954 9548 34960
rect 9404 34536 9456 34542
rect 9404 34478 9456 34484
rect 9312 34400 9364 34406
rect 9312 34342 9364 34348
rect 9324 33522 9352 34342
rect 9600 34134 9628 37130
rect 9680 36848 9732 36854
rect 9680 36790 9732 36796
rect 9692 34678 9720 36790
rect 10336 35834 10364 39200
rect 10690 37496 10746 37505
rect 10690 37431 10746 37440
rect 10704 37194 10732 37431
rect 10966 37360 11022 37369
rect 10966 37295 11022 37304
rect 11244 37324 11296 37330
rect 10782 37224 10838 37233
rect 10692 37188 10744 37194
rect 10782 37159 10838 37168
rect 10692 37130 10744 37136
rect 10692 36032 10744 36038
rect 10692 35974 10744 35980
rect 9772 35828 9824 35834
rect 9772 35770 9824 35776
rect 10324 35828 10376 35834
rect 10324 35770 10376 35776
rect 9680 34672 9732 34678
rect 9680 34614 9732 34620
rect 9680 34400 9732 34406
rect 9680 34342 9732 34348
rect 9588 34128 9640 34134
rect 9588 34070 9640 34076
rect 9312 33516 9364 33522
rect 9312 33458 9364 33464
rect 9692 33454 9720 34342
rect 9784 34202 9812 35770
rect 10598 35592 10654 35601
rect 10598 35527 10654 35536
rect 10612 35494 10640 35527
rect 10600 35488 10652 35494
rect 10600 35430 10652 35436
rect 10704 34746 10732 35974
rect 10796 35698 10824 37159
rect 10980 37126 11008 37295
rect 11244 37266 11296 37272
rect 10968 37120 11020 37126
rect 10968 37062 11020 37068
rect 11152 37120 11204 37126
rect 11152 37062 11204 37068
rect 11164 36854 11192 37062
rect 10968 36848 11020 36854
rect 10966 36816 10968 36825
rect 11152 36848 11204 36854
rect 11020 36816 11022 36825
rect 11152 36790 11204 36796
rect 10966 36751 11022 36760
rect 11060 36712 11112 36718
rect 11060 36654 11112 36660
rect 10968 36236 11020 36242
rect 10968 36178 11020 36184
rect 10980 36038 11008 36178
rect 11072 36174 11100 36654
rect 11060 36168 11112 36174
rect 11060 36110 11112 36116
rect 10876 36032 10928 36038
rect 10876 35974 10928 35980
rect 10968 36032 11020 36038
rect 10968 35974 11020 35980
rect 10888 35766 10916 35974
rect 10876 35760 10928 35766
rect 10876 35702 10928 35708
rect 10784 35692 10836 35698
rect 10784 35634 10836 35640
rect 10692 34740 10744 34746
rect 10692 34682 10744 34688
rect 10506 34640 10562 34649
rect 9864 34604 9916 34610
rect 10506 34575 10508 34584
rect 9864 34546 9916 34552
rect 10560 34575 10562 34584
rect 10508 34546 10560 34552
rect 9876 34354 9904 34546
rect 9876 34326 9996 34354
rect 9772 34196 9824 34202
rect 9824 34156 9904 34184
rect 9772 34138 9824 34144
rect 9680 33448 9732 33454
rect 9680 33390 9732 33396
rect 9312 33312 9364 33318
rect 9692 33300 9720 33390
rect 9364 33272 9720 33300
rect 9312 33254 9364 33260
rect 9312 32904 9364 32910
rect 9312 32846 9364 32852
rect 9220 32768 9272 32774
rect 9220 32710 9272 32716
rect 9036 32496 9088 32502
rect 9036 32438 9088 32444
rect 8760 32360 8812 32366
rect 8760 32302 8812 32308
rect 8772 31890 8800 32302
rect 8760 31884 8812 31890
rect 8760 31826 8812 31832
rect 8852 31408 8904 31414
rect 8852 31350 8904 31356
rect 8760 30864 8812 30870
rect 8760 30806 8812 30812
rect 8588 29158 8708 29186
rect 8588 28121 8616 29158
rect 8668 29028 8720 29034
rect 8668 28970 8720 28976
rect 8574 28112 8630 28121
rect 8574 28047 8630 28056
rect 8680 25770 8708 28970
rect 8772 27470 8800 30806
rect 8864 30598 8892 31350
rect 9128 31272 9180 31278
rect 9128 31214 9180 31220
rect 8852 30592 8904 30598
rect 8852 30534 8904 30540
rect 8760 27464 8812 27470
rect 8760 27406 8812 27412
rect 8772 26314 8800 27406
rect 8760 26308 8812 26314
rect 8760 26250 8812 26256
rect 8668 25764 8720 25770
rect 8668 25706 8720 25712
rect 8484 25152 8536 25158
rect 8484 25094 8536 25100
rect 8576 25152 8628 25158
rect 8576 25094 8628 25100
rect 8484 24812 8536 24818
rect 8484 24754 8536 24760
rect 8496 24585 8524 24754
rect 8482 24576 8538 24585
rect 8482 24511 8538 24520
rect 8496 24342 8524 24511
rect 8588 24410 8616 25094
rect 8680 24410 8708 25706
rect 8576 24404 8628 24410
rect 8576 24346 8628 24352
rect 8668 24404 8720 24410
rect 8668 24346 8720 24352
rect 8484 24336 8536 24342
rect 8484 24278 8536 24284
rect 8576 24132 8628 24138
rect 8576 24074 8628 24080
rect 8588 23526 8616 24074
rect 8772 24070 8800 26250
rect 8864 24936 8892 30534
rect 9140 30394 9168 31214
rect 9128 30388 9180 30394
rect 9128 30330 9180 30336
rect 9232 30326 9260 32710
rect 9324 32026 9352 32846
rect 9496 32768 9548 32774
rect 9496 32710 9548 32716
rect 9404 32360 9456 32366
rect 9404 32302 9456 32308
rect 9312 32020 9364 32026
rect 9312 31962 9364 31968
rect 9312 31816 9364 31822
rect 9312 31758 9364 31764
rect 9220 30320 9272 30326
rect 9220 30262 9272 30268
rect 9324 29238 9352 31758
rect 9416 31346 9444 32302
rect 9508 31754 9536 32710
rect 9588 31816 9640 31822
rect 9588 31758 9640 31764
rect 9496 31748 9548 31754
rect 9496 31690 9548 31696
rect 9404 31340 9456 31346
rect 9404 31282 9456 31288
rect 9416 30938 9444 31282
rect 9404 30932 9456 30938
rect 9404 30874 9456 30880
rect 9416 30802 9444 30874
rect 9404 30796 9456 30802
rect 9404 30738 9456 30744
rect 9600 30666 9628 31758
rect 9876 30870 9904 34156
rect 9968 33998 9996 34326
rect 10782 34232 10838 34241
rect 10782 34167 10838 34176
rect 10796 34134 10824 34167
rect 10784 34128 10836 34134
rect 10598 34096 10654 34105
rect 10784 34070 10836 34076
rect 10598 34031 10654 34040
rect 10612 33998 10640 34031
rect 9956 33992 10008 33998
rect 9956 33934 10008 33940
rect 10600 33992 10652 33998
rect 10600 33934 10652 33940
rect 9956 33448 10008 33454
rect 9956 33390 10008 33396
rect 9968 31793 9996 33390
rect 10506 33280 10562 33289
rect 10506 33215 10562 33224
rect 10520 32774 10548 33215
rect 10508 32768 10560 32774
rect 10508 32710 10560 32716
rect 10692 32768 10744 32774
rect 10692 32710 10744 32716
rect 10598 32600 10654 32609
rect 10598 32535 10654 32544
rect 10232 32020 10284 32026
rect 10232 31962 10284 31968
rect 10140 31816 10192 31822
rect 9954 31784 10010 31793
rect 10140 31758 10192 31764
rect 9954 31719 10010 31728
rect 9864 30864 9916 30870
rect 9864 30806 9916 30812
rect 9968 30734 9996 31719
rect 9956 30728 10008 30734
rect 9956 30670 10008 30676
rect 9588 30660 9640 30666
rect 9588 30602 9640 30608
rect 9586 29880 9642 29889
rect 9586 29815 9588 29824
rect 9640 29815 9642 29824
rect 9956 29844 10008 29850
rect 9588 29786 9640 29792
rect 9956 29786 10008 29792
rect 9680 29776 9732 29782
rect 9680 29718 9732 29724
rect 9404 29572 9456 29578
rect 9404 29514 9456 29520
rect 9416 29345 9444 29514
rect 9692 29481 9720 29718
rect 9678 29472 9734 29481
rect 9678 29407 9734 29416
rect 9402 29336 9458 29345
rect 9402 29271 9458 29280
rect 9496 29300 9548 29306
rect 9496 29242 9548 29248
rect 9312 29232 9364 29238
rect 9312 29174 9364 29180
rect 9404 29096 9456 29102
rect 9404 29038 9456 29044
rect 9416 28490 9444 29038
rect 9508 28490 9536 29242
rect 9864 28688 9916 28694
rect 9864 28630 9916 28636
rect 9586 28520 9642 28529
rect 9404 28484 9456 28490
rect 9404 28426 9456 28432
rect 9496 28484 9548 28490
rect 9586 28455 9642 28464
rect 9496 28426 9548 28432
rect 9600 28218 9628 28455
rect 9588 28212 9640 28218
rect 9588 28154 9640 28160
rect 9680 28144 9732 28150
rect 9680 28086 9732 28092
rect 9036 28008 9088 28014
rect 9036 27950 9088 27956
rect 9048 27470 9076 27950
rect 9494 27704 9550 27713
rect 9494 27639 9550 27648
rect 9310 27568 9366 27577
rect 9310 27503 9366 27512
rect 9324 27470 9352 27503
rect 9036 27464 9088 27470
rect 9036 27406 9088 27412
rect 9312 27464 9364 27470
rect 9312 27406 9364 27412
rect 9404 27464 9456 27470
rect 9404 27406 9456 27412
rect 9048 26858 9076 27406
rect 9140 27254 9352 27282
rect 9140 27062 9168 27254
rect 9218 27160 9274 27169
rect 9324 27130 9352 27254
rect 9218 27095 9274 27104
rect 9312 27124 9364 27130
rect 9232 27062 9260 27095
rect 9312 27066 9364 27072
rect 9128 27056 9180 27062
rect 9128 26998 9180 27004
rect 9220 27056 9272 27062
rect 9220 26998 9272 27004
rect 9128 26920 9180 26926
rect 9128 26862 9180 26868
rect 9036 26852 9088 26858
rect 9036 26794 9088 26800
rect 9048 26450 9076 26794
rect 9036 26444 9088 26450
rect 9036 26386 9088 26392
rect 9036 25968 9088 25974
rect 9140 25945 9168 26862
rect 9416 26382 9444 27406
rect 9404 26376 9456 26382
rect 9404 26318 9456 26324
rect 9312 26308 9364 26314
rect 9312 26250 9364 26256
rect 9220 26240 9272 26246
rect 9220 26182 9272 26188
rect 9036 25910 9088 25916
rect 9126 25936 9182 25945
rect 9048 25430 9076 25910
rect 9126 25871 9182 25880
rect 9232 25770 9260 26182
rect 9324 25974 9352 26250
rect 9508 26246 9536 27639
rect 9692 27334 9720 28086
rect 9876 27418 9904 28630
rect 9968 28082 9996 29786
rect 10152 29238 10180 31758
rect 10140 29232 10192 29238
rect 10140 29174 10192 29180
rect 10244 29034 10272 31962
rect 10612 31890 10640 32535
rect 10600 31884 10652 31890
rect 10600 31826 10652 31832
rect 10612 31793 10640 31826
rect 10598 31784 10654 31793
rect 10598 31719 10654 31728
rect 10704 31482 10732 32710
rect 10782 32192 10838 32201
rect 10782 32127 10838 32136
rect 10692 31476 10744 31482
rect 10692 31418 10744 31424
rect 10416 31136 10468 31142
rect 10416 31078 10468 31084
rect 10428 30802 10456 31078
rect 10508 30864 10560 30870
rect 10508 30806 10560 30812
rect 10416 30796 10468 30802
rect 10416 30738 10468 30744
rect 10416 29776 10468 29782
rect 10416 29718 10468 29724
rect 10324 29096 10376 29102
rect 10324 29038 10376 29044
rect 10232 29028 10284 29034
rect 10232 28970 10284 28976
rect 10140 28960 10192 28966
rect 10140 28902 10192 28908
rect 10152 28626 10180 28902
rect 10140 28620 10192 28626
rect 10140 28562 10192 28568
rect 9956 28076 10008 28082
rect 9956 28018 10008 28024
rect 9876 27390 9996 27418
rect 10152 27402 10180 28562
rect 10336 28422 10364 29038
rect 10324 28416 10376 28422
rect 10324 28358 10376 28364
rect 10336 28014 10364 28358
rect 10324 28008 10376 28014
rect 10324 27950 10376 27956
rect 10324 27600 10376 27606
rect 10324 27542 10376 27548
rect 9680 27328 9732 27334
rect 9680 27270 9732 27276
rect 9772 27328 9824 27334
rect 9772 27270 9824 27276
rect 9680 26852 9732 26858
rect 9680 26794 9732 26800
rect 9692 26466 9720 26794
rect 9784 26586 9812 27270
rect 9864 26852 9916 26858
rect 9864 26794 9916 26800
rect 9772 26580 9824 26586
rect 9772 26522 9824 26528
rect 9876 26466 9904 26794
rect 9692 26438 9904 26466
rect 9678 26344 9734 26353
rect 9678 26279 9680 26288
rect 9732 26279 9734 26288
rect 9680 26250 9732 26256
rect 9496 26240 9548 26246
rect 9496 26182 9548 26188
rect 9312 25968 9364 25974
rect 9312 25910 9364 25916
rect 9220 25764 9272 25770
rect 9220 25706 9272 25712
rect 9036 25424 9088 25430
rect 9036 25366 9088 25372
rect 9312 25424 9364 25430
rect 9312 25366 9364 25372
rect 9128 25220 9180 25226
rect 9128 25162 9180 25168
rect 8864 24908 8984 24936
rect 8852 24812 8904 24818
rect 8852 24754 8904 24760
rect 8864 24721 8892 24754
rect 8850 24712 8906 24721
rect 8850 24647 8906 24656
rect 8956 24256 8984 24908
rect 9140 24750 9168 25162
rect 9128 24744 9180 24750
rect 9128 24686 9180 24692
rect 9220 24744 9272 24750
rect 9220 24686 9272 24692
rect 8864 24228 8984 24256
rect 8760 24064 8812 24070
rect 8760 24006 8812 24012
rect 8864 23662 8892 24228
rect 8944 24132 8996 24138
rect 8944 24074 8996 24080
rect 8852 23656 8904 23662
rect 8852 23598 8904 23604
rect 8576 23520 8628 23526
rect 8576 23462 8628 23468
rect 8864 22234 8892 23598
rect 8852 22228 8904 22234
rect 8852 22170 8904 22176
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 8956 10810 8984 24074
rect 9036 23656 9088 23662
rect 9232 23633 9260 24686
rect 9324 24274 9352 25366
rect 9508 25362 9536 26182
rect 9772 25968 9824 25974
rect 9770 25936 9772 25945
rect 9824 25936 9826 25945
rect 9770 25871 9826 25880
rect 9772 25832 9824 25838
rect 9772 25774 9824 25780
rect 9496 25356 9548 25362
rect 9784 25344 9812 25774
rect 9876 25362 9904 26438
rect 9968 26382 9996 27390
rect 10140 27396 10192 27402
rect 10140 27338 10192 27344
rect 10048 26580 10100 26586
rect 10048 26522 10100 26528
rect 9956 26376 10008 26382
rect 9956 26318 10008 26324
rect 9496 25298 9548 25304
rect 9692 25316 9812 25344
rect 9864 25356 9916 25362
rect 9496 24880 9548 24886
rect 9692 24834 9720 25316
rect 9864 25298 9916 25304
rect 9772 25220 9824 25226
rect 9772 25162 9824 25168
rect 9496 24822 9548 24828
rect 9312 24268 9364 24274
rect 9312 24210 9364 24216
rect 9312 24132 9364 24138
rect 9312 24074 9364 24080
rect 9036 23598 9088 23604
rect 9218 23624 9274 23633
rect 9048 23186 9076 23598
rect 9218 23559 9274 23568
rect 9036 23180 9088 23186
rect 9036 23122 9088 23128
rect 9324 22710 9352 24074
rect 9508 23798 9536 24822
rect 9600 24806 9720 24834
rect 9600 24070 9628 24806
rect 9784 24698 9812 25162
rect 9692 24670 9812 24698
rect 9876 24698 9904 25298
rect 9876 24682 9996 24698
rect 9876 24676 10008 24682
rect 9876 24670 9956 24676
rect 9692 24614 9720 24670
rect 9956 24618 10008 24624
rect 9680 24608 9732 24614
rect 9680 24550 9732 24556
rect 9680 24404 9732 24410
rect 9680 24346 9732 24352
rect 9692 24274 9720 24346
rect 9680 24268 9732 24274
rect 9680 24210 9732 24216
rect 9588 24064 9640 24070
rect 9588 24006 9640 24012
rect 9496 23792 9548 23798
rect 9496 23734 9548 23740
rect 10060 23662 10088 26522
rect 10048 23656 10100 23662
rect 10048 23598 10100 23604
rect 9312 22704 9364 22710
rect 9312 22646 9364 22652
rect 9588 22636 9640 22642
rect 9588 22578 9640 22584
rect 9600 22234 9628 22578
rect 9588 22228 9640 22234
rect 9588 22170 9640 22176
rect 10152 22094 10180 27338
rect 10336 26926 10364 27542
rect 10324 26920 10376 26926
rect 10324 26862 10376 26868
rect 10324 26784 10376 26790
rect 10324 26726 10376 26732
rect 10336 26450 10364 26726
rect 10324 26444 10376 26450
rect 10324 26386 10376 26392
rect 10232 25152 10284 25158
rect 10230 25120 10232 25129
rect 10284 25120 10286 25129
rect 10230 25055 10286 25064
rect 10428 24177 10456 29718
rect 10414 24168 10470 24177
rect 10414 24103 10470 24112
rect 10324 23588 10376 23594
rect 10324 23530 10376 23536
rect 10336 23050 10364 23530
rect 10428 23497 10456 24103
rect 10414 23488 10470 23497
rect 10414 23423 10470 23432
rect 10520 23186 10548 30806
rect 10598 30696 10654 30705
rect 10598 30631 10654 30640
rect 10612 28558 10640 30631
rect 10796 30274 10824 32127
rect 10888 31346 10916 35702
rect 11072 35630 11100 36110
rect 11060 35624 11112 35630
rect 11060 35566 11112 35572
rect 11072 35154 11100 35566
rect 11060 35148 11112 35154
rect 11060 35090 11112 35096
rect 11072 34082 11100 35090
rect 11150 34912 11206 34921
rect 11150 34847 11206 34856
rect 11164 34610 11192 34847
rect 11152 34604 11204 34610
rect 11152 34546 11204 34552
rect 11072 34066 11192 34082
rect 11072 34060 11204 34066
rect 11072 34054 11152 34060
rect 11072 33522 11100 34054
rect 11152 34002 11204 34008
rect 11060 33516 11112 33522
rect 11060 33458 11112 33464
rect 11072 32978 11100 33458
rect 11152 33108 11204 33114
rect 11152 33050 11204 33056
rect 11060 32972 11112 32978
rect 11060 32914 11112 32920
rect 10968 32224 11020 32230
rect 10968 32166 11020 32172
rect 10876 31340 10928 31346
rect 10876 31282 10928 31288
rect 10980 31210 11008 32166
rect 11072 31890 11100 32914
rect 11164 32434 11192 33050
rect 11152 32428 11204 32434
rect 11152 32370 11204 32376
rect 11060 31884 11112 31890
rect 11060 31826 11112 31832
rect 10968 31204 11020 31210
rect 10968 31146 11020 31152
rect 11256 30938 11284 37266
rect 11704 37120 11756 37126
rect 11704 37062 11756 37068
rect 11716 36802 11744 37062
rect 11886 36952 11942 36961
rect 11886 36887 11888 36896
rect 11940 36887 11942 36896
rect 11888 36858 11940 36864
rect 11624 36786 11744 36802
rect 11612 36780 11744 36786
rect 11664 36774 11744 36780
rect 11612 36722 11664 36728
rect 11612 36644 11664 36650
rect 11612 36586 11664 36592
rect 11624 36378 11652 36586
rect 11612 36372 11664 36378
rect 11612 36314 11664 36320
rect 11612 36236 11664 36242
rect 11612 36178 11664 36184
rect 11624 35834 11652 36178
rect 11612 35828 11664 35834
rect 11612 35770 11664 35776
rect 11612 34400 11664 34406
rect 11612 34342 11664 34348
rect 11334 33960 11390 33969
rect 11334 33895 11390 33904
rect 11428 33924 11480 33930
rect 11348 33318 11376 33895
rect 11428 33866 11480 33872
rect 11440 33658 11468 33866
rect 11624 33862 11652 34342
rect 11520 33856 11572 33862
rect 11520 33798 11572 33804
rect 11612 33856 11664 33862
rect 11612 33798 11664 33804
rect 11428 33652 11480 33658
rect 11428 33594 11480 33600
rect 11336 33312 11388 33318
rect 11336 33254 11388 33260
rect 11532 32978 11560 33798
rect 11520 32972 11572 32978
rect 11520 32914 11572 32920
rect 11428 32836 11480 32842
rect 11428 32778 11480 32784
rect 11336 31680 11388 31686
rect 11336 31622 11388 31628
rect 11348 31278 11376 31622
rect 11336 31272 11388 31278
rect 11336 31214 11388 31220
rect 11060 30932 11112 30938
rect 11060 30874 11112 30880
rect 11244 30932 11296 30938
rect 11244 30874 11296 30880
rect 10876 30864 10928 30870
rect 10876 30806 10928 30812
rect 10704 30246 10824 30274
rect 10704 30054 10732 30246
rect 10888 30190 10916 30806
rect 10784 30184 10836 30190
rect 10784 30126 10836 30132
rect 10876 30184 10928 30190
rect 10876 30126 10928 30132
rect 10692 30048 10744 30054
rect 10692 29990 10744 29996
rect 10704 29050 10732 29990
rect 10796 29209 10824 30126
rect 10876 30048 10928 30054
rect 10876 29990 10928 29996
rect 10888 29578 10916 29990
rect 10876 29572 10928 29578
rect 10876 29514 10928 29520
rect 10888 29238 10916 29514
rect 10876 29232 10928 29238
rect 10782 29200 10838 29209
rect 10876 29174 10928 29180
rect 10782 29135 10838 29144
rect 10704 29022 10916 29050
rect 10600 28552 10652 28558
rect 10600 28494 10652 28500
rect 10612 27418 10640 28494
rect 10692 28144 10744 28150
rect 10692 28086 10744 28092
rect 10704 27674 10732 28086
rect 10784 27940 10836 27946
rect 10784 27882 10836 27888
rect 10692 27668 10744 27674
rect 10692 27610 10744 27616
rect 10612 27390 10732 27418
rect 10600 27056 10652 27062
rect 10600 26998 10652 27004
rect 10612 25770 10640 26998
rect 10704 26330 10732 27390
rect 10796 26450 10824 27882
rect 10888 26489 10916 29022
rect 10968 28688 11020 28694
rect 10968 28630 11020 28636
rect 10980 27062 11008 28630
rect 11072 28422 11100 30874
rect 11256 30734 11284 30874
rect 11244 30728 11296 30734
rect 11244 30670 11296 30676
rect 11336 30320 11388 30326
rect 11336 30262 11388 30268
rect 11150 29336 11206 29345
rect 11150 29271 11206 29280
rect 11164 29170 11192 29271
rect 11152 29164 11204 29170
rect 11152 29106 11204 29112
rect 11244 29028 11296 29034
rect 11244 28970 11296 28976
rect 11256 28626 11284 28970
rect 11244 28620 11296 28626
rect 11244 28562 11296 28568
rect 11060 28416 11112 28422
rect 11060 28358 11112 28364
rect 11060 27940 11112 27946
rect 11060 27882 11112 27888
rect 11072 27130 11100 27882
rect 11244 27396 11296 27402
rect 11244 27338 11296 27344
rect 11256 27130 11284 27338
rect 11060 27124 11112 27130
rect 11060 27066 11112 27072
rect 11244 27124 11296 27130
rect 11244 27066 11296 27072
rect 10968 27056 11020 27062
rect 10968 26998 11020 27004
rect 10874 26480 10930 26489
rect 10784 26444 10836 26450
rect 10874 26415 10930 26424
rect 10784 26386 10836 26392
rect 10704 26302 10824 26330
rect 10600 25764 10652 25770
rect 10600 25706 10652 25712
rect 10600 24880 10652 24886
rect 10600 24822 10652 24828
rect 10508 23180 10560 23186
rect 10508 23122 10560 23128
rect 10324 23044 10376 23050
rect 10324 22986 10376 22992
rect 10416 23044 10468 23050
rect 10416 22986 10468 22992
rect 10232 22636 10284 22642
rect 10232 22578 10284 22584
rect 10060 22066 10180 22094
rect 10060 15502 10088 22066
rect 10244 21486 10272 22578
rect 10232 21480 10284 21486
rect 10232 21422 10284 21428
rect 10336 20602 10364 22986
rect 10428 22778 10456 22986
rect 10416 22772 10468 22778
rect 10416 22714 10468 22720
rect 10520 22642 10548 23122
rect 10612 22710 10640 24822
rect 10692 24200 10744 24206
rect 10692 24142 10744 24148
rect 10704 23254 10732 24142
rect 10692 23248 10744 23254
rect 10692 23190 10744 23196
rect 10796 23186 10824 26302
rect 10966 25936 11022 25945
rect 10966 25871 10968 25880
rect 11020 25871 11022 25880
rect 10968 25842 11020 25848
rect 11150 24712 11206 24721
rect 11150 24647 11206 24656
rect 10876 24200 10928 24206
rect 10876 24142 10928 24148
rect 10784 23180 10836 23186
rect 10784 23122 10836 23128
rect 10600 22704 10652 22710
rect 10600 22646 10652 22652
rect 10508 22636 10560 22642
rect 10508 22578 10560 22584
rect 10416 22092 10468 22098
rect 10416 22034 10468 22040
rect 10324 20596 10376 20602
rect 10324 20538 10376 20544
rect 10428 20482 10456 22034
rect 10600 21956 10652 21962
rect 10600 21898 10652 21904
rect 10692 21956 10744 21962
rect 10692 21898 10744 21904
rect 10508 21888 10560 21894
rect 10508 21830 10560 21836
rect 10520 21554 10548 21830
rect 10612 21622 10640 21898
rect 10704 21622 10732 21898
rect 10600 21616 10652 21622
rect 10600 21558 10652 21564
rect 10692 21616 10744 21622
rect 10692 21558 10744 21564
rect 10508 21548 10560 21554
rect 10508 21490 10560 21496
rect 10508 20800 10560 20806
rect 10508 20742 10560 20748
rect 10336 20454 10456 20482
rect 10520 20466 10548 20742
rect 10508 20460 10560 20466
rect 10336 20398 10364 20454
rect 10508 20402 10560 20408
rect 10600 20460 10652 20466
rect 10600 20402 10652 20408
rect 10324 20392 10376 20398
rect 10324 20334 10376 20340
rect 10048 15496 10100 15502
rect 10048 15438 10100 15444
rect 10336 13938 10364 20334
rect 10324 13932 10376 13938
rect 10324 13874 10376 13880
rect 8944 10804 8996 10810
rect 8944 10746 8996 10752
rect 8668 10668 8720 10674
rect 8668 10610 8720 10616
rect 8680 3058 8708 10610
rect 10520 7342 10548 20402
rect 10612 19718 10640 20402
rect 10888 20058 10916 24142
rect 11060 23656 11112 23662
rect 11060 23598 11112 23604
rect 10966 23488 11022 23497
rect 10966 23423 11022 23432
rect 10980 23118 11008 23423
rect 11072 23322 11100 23598
rect 11060 23316 11112 23322
rect 11060 23258 11112 23264
rect 10968 23112 11020 23118
rect 10968 23054 11020 23060
rect 11164 23050 11192 24647
rect 11256 23798 11284 27066
rect 11244 23792 11296 23798
rect 11244 23734 11296 23740
rect 11152 23044 11204 23050
rect 11152 22986 11204 22992
rect 11244 22636 11296 22642
rect 11244 22578 11296 22584
rect 10968 22432 11020 22438
rect 10968 22374 11020 22380
rect 10876 20052 10928 20058
rect 10876 19994 10928 20000
rect 10980 19786 11008 22374
rect 11060 21480 11112 21486
rect 11060 21422 11112 21428
rect 11072 20602 11100 21422
rect 11256 21350 11284 22578
rect 11348 22094 11376 30262
rect 11440 28490 11468 32778
rect 11610 32736 11666 32745
rect 11610 32671 11666 32680
rect 11518 32600 11574 32609
rect 11518 32535 11574 32544
rect 11532 32298 11560 32535
rect 11624 32502 11652 32671
rect 11612 32496 11664 32502
rect 11612 32438 11664 32444
rect 11520 32292 11572 32298
rect 11520 32234 11572 32240
rect 11716 31929 11744 36774
rect 11796 36576 11848 36582
rect 11796 36518 11848 36524
rect 11808 33930 11836 36518
rect 11888 36100 11940 36106
rect 11888 36042 11940 36048
rect 11900 35057 11928 36042
rect 12070 35456 12126 35465
rect 12070 35391 12126 35400
rect 11886 35048 11942 35057
rect 11886 34983 11942 34992
rect 11980 34400 12032 34406
rect 11980 34342 12032 34348
rect 11796 33924 11848 33930
rect 11796 33866 11848 33872
rect 11702 31920 11758 31929
rect 11702 31855 11758 31864
rect 11702 31512 11758 31521
rect 11702 31447 11758 31456
rect 11716 31414 11744 31447
rect 11704 31408 11756 31414
rect 11704 31350 11756 31356
rect 11704 31272 11756 31278
rect 11704 31214 11756 31220
rect 11612 31136 11664 31142
rect 11612 31078 11664 31084
rect 11520 30116 11572 30122
rect 11520 30058 11572 30064
rect 11532 29714 11560 30058
rect 11520 29708 11572 29714
rect 11520 29650 11572 29656
rect 11518 29608 11574 29617
rect 11518 29543 11520 29552
rect 11572 29543 11574 29552
rect 11520 29514 11572 29520
rect 11428 28484 11480 28490
rect 11428 28426 11480 28432
rect 11520 28484 11572 28490
rect 11520 28426 11572 28432
rect 11532 27674 11560 28426
rect 11520 27668 11572 27674
rect 11520 27610 11572 27616
rect 11520 26376 11572 26382
rect 11520 26318 11572 26324
rect 11428 25356 11480 25362
rect 11532 25344 11560 26318
rect 11480 25316 11560 25344
rect 11428 25298 11480 25304
rect 11428 25152 11480 25158
rect 11428 25094 11480 25100
rect 11440 24614 11468 25094
rect 11532 24750 11560 25316
rect 11520 24744 11572 24750
rect 11520 24686 11572 24692
rect 11428 24608 11480 24614
rect 11428 24550 11480 24556
rect 11624 23798 11652 31078
rect 11716 30190 11744 31214
rect 11704 30184 11756 30190
rect 11704 30126 11756 30132
rect 11704 28688 11756 28694
rect 11704 28630 11756 28636
rect 11716 28490 11744 28630
rect 11704 28484 11756 28490
rect 11704 28426 11756 28432
rect 11808 25906 11836 33866
rect 11992 33454 12020 34342
rect 12084 33833 12112 35391
rect 12268 35018 12296 39200
rect 13176 37664 13228 37670
rect 13176 37606 13228 37612
rect 13188 37330 13216 37606
rect 13176 37324 13228 37330
rect 13176 37266 13228 37272
rect 12530 37224 12586 37233
rect 12530 37159 12586 37168
rect 12716 37188 12768 37194
rect 12544 37126 12572 37159
rect 12716 37130 12768 37136
rect 12900 37188 12952 37194
rect 12900 37130 12952 37136
rect 12532 37120 12584 37126
rect 12532 37062 12584 37068
rect 12728 36310 12756 37130
rect 12912 36961 12940 37130
rect 12898 36952 12954 36961
rect 12898 36887 12954 36896
rect 13084 36644 13136 36650
rect 13084 36586 13136 36592
rect 12992 36576 13044 36582
rect 12992 36518 13044 36524
rect 12716 36304 12768 36310
rect 12716 36246 12768 36252
rect 12624 36236 12676 36242
rect 12624 36178 12676 36184
rect 12636 35630 12664 36178
rect 12624 35624 12676 35630
rect 12624 35566 12676 35572
rect 13004 35442 13032 36518
rect 13096 36242 13124 36586
rect 13084 36236 13136 36242
rect 13084 36178 13136 36184
rect 13452 36100 13504 36106
rect 13452 36042 13504 36048
rect 13176 36032 13228 36038
rect 13176 35974 13228 35980
rect 13268 36032 13320 36038
rect 13268 35974 13320 35980
rect 13084 35556 13136 35562
rect 13084 35498 13136 35504
rect 12820 35414 13032 35442
rect 12346 35320 12402 35329
rect 12346 35255 12402 35264
rect 12256 35012 12308 35018
rect 12256 34954 12308 34960
rect 12360 34950 12388 35255
rect 12348 34944 12400 34950
rect 12348 34886 12400 34892
rect 12532 34944 12584 34950
rect 12532 34886 12584 34892
rect 12164 34740 12216 34746
rect 12164 34682 12216 34688
rect 12176 34066 12204 34682
rect 12346 34232 12402 34241
rect 12346 34167 12348 34176
rect 12400 34167 12402 34176
rect 12348 34138 12400 34144
rect 12440 34128 12492 34134
rect 12438 34096 12440 34105
rect 12492 34096 12494 34105
rect 12164 34060 12216 34066
rect 12438 34031 12494 34040
rect 12164 34002 12216 34008
rect 12438 33960 12494 33969
rect 12438 33895 12440 33904
rect 12492 33895 12494 33904
rect 12440 33866 12492 33872
rect 12070 33824 12126 33833
rect 12544 33810 12572 34886
rect 12820 34241 12848 35414
rect 13096 35290 13124 35498
rect 13084 35284 13136 35290
rect 13084 35226 13136 35232
rect 13082 34640 13138 34649
rect 13082 34575 13138 34584
rect 13096 34542 13124 34575
rect 13084 34536 13136 34542
rect 13084 34478 13136 34484
rect 12806 34232 12862 34241
rect 12806 34167 12862 34176
rect 13188 33844 13216 35974
rect 13280 35086 13308 35974
rect 13268 35080 13320 35086
rect 13268 35022 13320 35028
rect 13268 34672 13320 34678
rect 13268 34614 13320 34620
rect 13280 33998 13308 34614
rect 13464 34377 13492 36042
rect 13556 34610 13584 39200
rect 15488 39114 15516 39200
rect 15580 39114 15608 39222
rect 15488 39086 15608 39114
rect 14280 37732 14332 37738
rect 14280 37674 14332 37680
rect 14004 37256 14056 37262
rect 14292 37210 14320 37674
rect 14556 37324 14608 37330
rect 14556 37266 14608 37272
rect 14004 37198 14056 37204
rect 14016 36718 14044 37198
rect 14200 37194 14320 37210
rect 14188 37188 14320 37194
rect 14240 37182 14320 37188
rect 14188 37130 14240 37136
rect 14004 36712 14056 36718
rect 14004 36654 14056 36660
rect 13726 36408 13782 36417
rect 13726 36343 13728 36352
rect 13780 36343 13782 36352
rect 13728 36314 13780 36320
rect 14016 36224 14044 36654
rect 14292 36582 14320 37182
rect 14568 36922 14596 37266
rect 14646 37224 14702 37233
rect 14646 37159 14648 37168
rect 14700 37159 14702 37168
rect 14648 37130 14700 37136
rect 15106 37088 15162 37097
rect 15106 37023 15162 37032
rect 14556 36916 14608 36922
rect 14556 36858 14608 36864
rect 14280 36576 14332 36582
rect 14280 36518 14332 36524
rect 14280 36236 14332 36242
rect 14016 36196 14280 36224
rect 14280 36178 14332 36184
rect 13912 36032 13964 36038
rect 13912 35974 13964 35980
rect 13818 35864 13874 35873
rect 13818 35799 13874 35808
rect 13832 35630 13860 35799
rect 13820 35624 13872 35630
rect 13820 35566 13872 35572
rect 13636 35488 13688 35494
rect 13636 35430 13688 35436
rect 13544 34604 13596 34610
rect 13544 34546 13596 34552
rect 13648 34542 13676 35430
rect 13924 35329 13952 35974
rect 14096 35692 14148 35698
rect 14096 35634 14148 35640
rect 13910 35320 13966 35329
rect 13910 35255 13966 35264
rect 13820 35080 13872 35086
rect 13820 35022 13872 35028
rect 13728 35012 13780 35018
rect 13728 34954 13780 34960
rect 13740 34921 13768 34954
rect 13726 34912 13782 34921
rect 13726 34847 13782 34856
rect 13636 34536 13688 34542
rect 13636 34478 13688 34484
rect 13450 34368 13506 34377
rect 13450 34303 13506 34312
rect 13268 33992 13320 33998
rect 13268 33934 13320 33940
rect 13544 33992 13596 33998
rect 13544 33934 13596 33940
rect 13188 33816 13308 33844
rect 12544 33782 12756 33810
rect 12070 33759 12126 33768
rect 12256 33584 12308 33590
rect 12308 33544 12480 33572
rect 12256 33526 12308 33532
rect 11980 33448 12032 33454
rect 11980 33390 12032 33396
rect 11992 33130 12020 33390
rect 11900 33102 12020 33130
rect 11900 28762 11928 33102
rect 12164 32972 12216 32978
rect 12164 32914 12216 32920
rect 11978 32600 12034 32609
rect 11978 32535 12034 32544
rect 11992 29238 12020 32535
rect 12072 32360 12124 32366
rect 12070 32328 12072 32337
rect 12124 32328 12126 32337
rect 12070 32263 12126 32272
rect 12072 32224 12124 32230
rect 12072 32166 12124 32172
rect 12084 32026 12112 32166
rect 12072 32020 12124 32026
rect 12072 31962 12124 31968
rect 12070 31920 12126 31929
rect 12070 31855 12126 31864
rect 12084 30569 12112 31855
rect 12070 30560 12126 30569
rect 12070 30495 12126 30504
rect 11980 29232 12032 29238
rect 11980 29174 12032 29180
rect 11992 28966 12020 29174
rect 11980 28960 12032 28966
rect 11980 28902 12032 28908
rect 11888 28756 11940 28762
rect 11888 28698 11940 28704
rect 11980 28688 12032 28694
rect 11980 28630 12032 28636
rect 11992 28218 12020 28630
rect 11980 28212 12032 28218
rect 11980 28154 12032 28160
rect 11888 27328 11940 27334
rect 11888 27270 11940 27276
rect 11900 27062 11928 27270
rect 11888 27056 11940 27062
rect 11888 26998 11940 27004
rect 11888 26580 11940 26586
rect 11888 26522 11940 26528
rect 11900 26382 11928 26522
rect 11888 26376 11940 26382
rect 11888 26318 11940 26324
rect 11796 25900 11848 25906
rect 11796 25842 11848 25848
rect 11704 25424 11756 25430
rect 11704 25366 11756 25372
rect 11716 25226 11744 25366
rect 11704 25220 11756 25226
rect 11704 25162 11756 25168
rect 11704 24064 11756 24070
rect 11704 24006 11756 24012
rect 11716 23866 11744 24006
rect 11704 23860 11756 23866
rect 11704 23802 11756 23808
rect 11612 23792 11664 23798
rect 11612 23734 11664 23740
rect 11716 23322 11744 23802
rect 11704 23316 11756 23322
rect 11704 23258 11756 23264
rect 11520 22976 11572 22982
rect 11520 22918 11572 22924
rect 11532 22778 11560 22918
rect 11520 22772 11572 22778
rect 11520 22714 11572 22720
rect 11716 22098 11744 23258
rect 11808 23186 11836 25842
rect 11888 25696 11940 25702
rect 11888 25638 11940 25644
rect 11900 24886 11928 25638
rect 12176 25344 12204 32914
rect 12256 32768 12308 32774
rect 12256 32710 12308 32716
rect 12268 31754 12296 32710
rect 12452 32026 12480 33544
rect 12728 33300 12756 33782
rect 13176 33448 13228 33454
rect 13176 33390 13228 33396
rect 12544 33272 12756 33300
rect 12440 32020 12492 32026
rect 12440 31962 12492 31968
rect 12544 31754 12572 33272
rect 12624 33040 12676 33046
rect 12624 32982 12676 32988
rect 12636 32910 12664 32982
rect 12624 32904 12676 32910
rect 12624 32846 12676 32852
rect 12900 32564 12952 32570
rect 12900 32506 12952 32512
rect 12808 32360 12860 32366
rect 12808 32302 12860 32308
rect 12820 32201 12848 32302
rect 12806 32192 12862 32201
rect 12806 32127 12862 32136
rect 12256 31748 12308 31754
rect 12544 31726 12664 31754
rect 12256 31690 12308 31696
rect 12268 31090 12296 31690
rect 12532 31680 12584 31686
rect 12532 31622 12584 31628
rect 12544 31521 12572 31622
rect 12530 31512 12586 31521
rect 12530 31447 12586 31456
rect 12268 31062 12480 31090
rect 12348 30932 12400 30938
rect 12348 30874 12400 30880
rect 12360 30841 12388 30874
rect 12346 30832 12402 30841
rect 12346 30767 12402 30776
rect 12256 30660 12308 30666
rect 12256 30602 12308 30608
rect 12268 30394 12296 30602
rect 12256 30388 12308 30394
rect 12256 30330 12308 30336
rect 12452 29510 12480 31062
rect 12636 30410 12664 31726
rect 12716 31408 12768 31414
rect 12716 31350 12768 31356
rect 12728 30938 12756 31350
rect 12808 31136 12860 31142
rect 12808 31078 12860 31084
rect 12716 30932 12768 30938
rect 12716 30874 12768 30880
rect 12820 30666 12848 31078
rect 12808 30660 12860 30666
rect 12808 30602 12860 30608
rect 12544 30382 12664 30410
rect 12714 30424 12770 30433
rect 12544 30190 12572 30382
rect 12714 30359 12770 30368
rect 12728 30326 12756 30359
rect 12716 30320 12768 30326
rect 12716 30262 12768 30268
rect 12532 30184 12584 30190
rect 12532 30126 12584 30132
rect 12530 29880 12586 29889
rect 12530 29815 12532 29824
rect 12584 29815 12586 29824
rect 12532 29786 12584 29792
rect 12912 29782 12940 32506
rect 12992 32496 13044 32502
rect 12992 32438 13044 32444
rect 13004 31890 13032 32438
rect 12992 31884 13044 31890
rect 12992 31826 13044 31832
rect 13004 31090 13032 31826
rect 13188 31498 13216 33390
rect 13280 32842 13308 33816
rect 13556 33590 13584 33934
rect 13452 33584 13504 33590
rect 13452 33526 13504 33532
rect 13544 33584 13596 33590
rect 13544 33526 13596 33532
rect 13464 32978 13492 33526
rect 13452 32972 13504 32978
rect 13452 32914 13504 32920
rect 13360 32904 13412 32910
rect 13360 32846 13412 32852
rect 13268 32836 13320 32842
rect 13268 32778 13320 32784
rect 13280 32745 13308 32778
rect 13266 32736 13322 32745
rect 13266 32671 13322 32680
rect 13372 31890 13400 32846
rect 13452 32020 13504 32026
rect 13452 31962 13504 31968
rect 13544 32020 13596 32026
rect 13544 31962 13596 31968
rect 13360 31884 13412 31890
rect 13360 31826 13412 31832
rect 13372 31657 13400 31826
rect 13358 31648 13414 31657
rect 13358 31583 13414 31592
rect 13188 31470 13308 31498
rect 13176 31408 13228 31414
rect 13176 31350 13228 31356
rect 13188 31278 13216 31350
rect 13280 31278 13308 31470
rect 13176 31272 13228 31278
rect 13176 31214 13228 31220
rect 13268 31272 13320 31278
rect 13268 31214 13320 31220
rect 13084 31136 13136 31142
rect 13004 31084 13084 31090
rect 13004 31078 13136 31084
rect 13004 31062 13124 31078
rect 13004 30734 13032 31062
rect 13280 30818 13308 31214
rect 13280 30790 13400 30818
rect 12992 30728 13044 30734
rect 12992 30670 13044 30676
rect 13176 30728 13228 30734
rect 13176 30670 13228 30676
rect 13004 30054 13032 30670
rect 13084 30592 13136 30598
rect 13084 30534 13136 30540
rect 12992 30048 13044 30054
rect 12992 29990 13044 29996
rect 12900 29776 12952 29782
rect 12900 29718 12952 29724
rect 12990 29744 13046 29753
rect 12990 29679 13046 29688
rect 12256 29504 12308 29510
rect 12256 29446 12308 29452
rect 12440 29504 12492 29510
rect 12440 29446 12492 29452
rect 12808 29504 12860 29510
rect 12808 29446 12860 29452
rect 12268 28082 12296 29446
rect 12624 28620 12676 28626
rect 12624 28562 12676 28568
rect 12636 28490 12664 28562
rect 12624 28484 12676 28490
rect 12624 28426 12676 28432
rect 12256 28076 12308 28082
rect 12256 28018 12308 28024
rect 12268 26926 12296 28018
rect 12440 27532 12492 27538
rect 12440 27474 12492 27480
rect 12256 26920 12308 26926
rect 12256 26862 12308 26868
rect 12452 26586 12480 27474
rect 12820 26790 12848 29446
rect 12900 28008 12952 28014
rect 12900 27950 12952 27956
rect 12912 27538 12940 27950
rect 13004 27554 13032 29679
rect 13096 29578 13124 30534
rect 13188 30190 13216 30670
rect 13268 30660 13320 30666
rect 13268 30602 13320 30608
rect 13176 30184 13228 30190
rect 13176 30126 13228 30132
rect 13084 29572 13136 29578
rect 13084 29514 13136 29520
rect 13188 29034 13216 30126
rect 13176 29028 13228 29034
rect 13176 28970 13228 28976
rect 12900 27532 12952 27538
rect 13004 27526 13216 27554
rect 12900 27474 12952 27480
rect 12808 26784 12860 26790
rect 12808 26726 12860 26732
rect 12440 26580 12492 26586
rect 12440 26522 12492 26528
rect 12912 26382 12940 27474
rect 13084 27396 13136 27402
rect 13084 27338 13136 27344
rect 12992 27328 13044 27334
rect 12992 27270 13044 27276
rect 12900 26376 12952 26382
rect 12900 26318 12952 26324
rect 12716 26240 12768 26246
rect 12716 26182 12768 26188
rect 12440 25764 12492 25770
rect 12440 25706 12492 25712
rect 12452 25362 12480 25706
rect 12532 25696 12584 25702
rect 12532 25638 12584 25644
rect 12084 25316 12204 25344
rect 12440 25356 12492 25362
rect 11888 24880 11940 24886
rect 11888 24822 11940 24828
rect 11796 23180 11848 23186
rect 11796 23122 11848 23128
rect 11348 22066 11652 22094
rect 11624 21842 11652 22066
rect 11704 22092 11756 22098
rect 11704 22034 11756 22040
rect 12084 21962 12112 25316
rect 12440 25298 12492 25304
rect 12544 24274 12572 25638
rect 12624 25492 12676 25498
rect 12624 25434 12676 25440
rect 12636 25401 12664 25434
rect 12622 25392 12678 25401
rect 12622 25327 12678 25336
rect 12728 24886 12756 26182
rect 12900 25764 12952 25770
rect 12900 25706 12952 25712
rect 12716 24880 12768 24886
rect 12716 24822 12768 24828
rect 12912 24818 12940 25706
rect 12900 24812 12952 24818
rect 12900 24754 12952 24760
rect 13004 24682 13032 27270
rect 13096 27062 13124 27338
rect 13084 27056 13136 27062
rect 13084 26998 13136 27004
rect 13084 26512 13136 26518
rect 13084 26454 13136 26460
rect 13096 25974 13124 26454
rect 13084 25968 13136 25974
rect 13084 25910 13136 25916
rect 13188 25702 13216 27526
rect 13176 25696 13228 25702
rect 13176 25638 13228 25644
rect 13084 25356 13136 25362
rect 13084 25298 13136 25304
rect 13096 24750 13124 25298
rect 13280 24750 13308 30602
rect 13372 29753 13400 30790
rect 13358 29744 13414 29753
rect 13358 29679 13414 29688
rect 13360 29572 13412 29578
rect 13360 29514 13412 29520
rect 13372 29306 13400 29514
rect 13360 29300 13412 29306
rect 13360 29242 13412 29248
rect 13360 28960 13412 28966
rect 13360 28902 13412 28908
rect 13372 28762 13400 28902
rect 13360 28756 13412 28762
rect 13360 28698 13412 28704
rect 13464 26994 13492 31962
rect 13556 28694 13584 31962
rect 13648 31958 13676 34478
rect 13728 33856 13780 33862
rect 13728 33798 13780 33804
rect 13636 31952 13688 31958
rect 13636 31894 13688 31900
rect 13636 31816 13688 31822
rect 13636 31758 13688 31764
rect 13648 29073 13676 31758
rect 13740 31736 13768 33798
rect 13832 32337 13860 35022
rect 13924 33425 13952 35255
rect 14108 34678 14136 35634
rect 14292 35494 14320 36178
rect 15120 36106 15148 37023
rect 15764 36922 15792 39222
rect 16762 39200 16818 39800
rect 18694 39200 18750 39800
rect 20626 39200 20682 39800
rect 21914 39200 21970 39800
rect 23846 39200 23902 39800
rect 25134 39200 25190 39800
rect 27066 39200 27122 39800
rect 28998 39200 29054 39800
rect 30286 39200 30342 39800
rect 32218 39200 32274 39800
rect 33506 39200 33562 39800
rect 35438 39200 35494 39800
rect 37370 39200 37426 39800
rect 38658 39200 38714 39800
rect 16120 37664 16172 37670
rect 16120 37606 16172 37612
rect 16488 37664 16540 37670
rect 16488 37606 16540 37612
rect 16028 37392 16080 37398
rect 16026 37360 16028 37369
rect 16080 37360 16082 37369
rect 16026 37295 16082 37304
rect 16040 37126 16068 37295
rect 16028 37120 16080 37126
rect 16028 37062 16080 37068
rect 15752 36916 15804 36922
rect 15752 36858 15804 36864
rect 16132 36582 16160 37606
rect 16396 37392 16448 37398
rect 16302 37360 16358 37369
rect 16396 37334 16448 37340
rect 16302 37295 16358 37304
rect 16316 36582 16344 37295
rect 16120 36576 16172 36582
rect 16120 36518 16172 36524
rect 16304 36576 16356 36582
rect 16304 36518 16356 36524
rect 15108 36100 15160 36106
rect 15108 36042 15160 36048
rect 15752 36100 15804 36106
rect 15752 36042 15804 36048
rect 15014 36000 15070 36009
rect 15120 35986 15148 36042
rect 15764 36009 15792 36042
rect 15070 35958 15148 35986
rect 15750 36000 15806 36009
rect 15014 35935 15070 35944
rect 15750 35935 15806 35944
rect 15750 35864 15806 35873
rect 15750 35799 15806 35808
rect 14924 35760 14976 35766
rect 14924 35702 14976 35708
rect 15108 35760 15160 35766
rect 15108 35702 15160 35708
rect 15476 35760 15528 35766
rect 15476 35702 15528 35708
rect 14936 35601 14964 35702
rect 14922 35592 14978 35601
rect 14372 35556 14424 35562
rect 14922 35527 14978 35536
rect 14372 35498 14424 35504
rect 14280 35488 14332 35494
rect 14280 35430 14332 35436
rect 14188 35284 14240 35290
rect 14188 35226 14240 35232
rect 14200 34785 14228 35226
rect 14292 34950 14320 35430
rect 14384 35222 14412 35498
rect 15014 35320 15070 35329
rect 15014 35255 15070 35264
rect 14372 35216 14424 35222
rect 14372 35158 14424 35164
rect 15028 35086 15056 35255
rect 15016 35080 15068 35086
rect 15016 35022 15068 35028
rect 14280 34944 14332 34950
rect 14280 34886 14332 34892
rect 15016 34944 15068 34950
rect 15016 34886 15068 34892
rect 14186 34776 14242 34785
rect 14292 34746 14320 34886
rect 14646 34776 14702 34785
rect 14186 34711 14242 34720
rect 14280 34740 14332 34746
rect 14280 34682 14332 34688
rect 14372 34740 14424 34746
rect 14646 34711 14702 34720
rect 14372 34682 14424 34688
rect 14096 34672 14148 34678
rect 14384 34626 14412 34682
rect 14096 34614 14148 34620
rect 14200 34598 14412 34626
rect 14660 34610 14688 34711
rect 14830 34640 14886 34649
rect 14648 34604 14700 34610
rect 13910 33416 13966 33425
rect 13910 33351 13966 33360
rect 13818 32328 13874 32337
rect 13818 32263 13874 32272
rect 14200 32065 14228 34598
rect 14830 34575 14832 34584
rect 14648 34546 14700 34552
rect 14884 34575 14886 34584
rect 14832 34546 14884 34552
rect 14556 34536 14608 34542
rect 14556 34478 14608 34484
rect 14280 34196 14332 34202
rect 14280 34138 14332 34144
rect 14372 34196 14424 34202
rect 14372 34138 14424 34144
rect 14292 33862 14320 34138
rect 14280 33856 14332 33862
rect 14280 33798 14332 33804
rect 14384 33658 14412 34138
rect 14372 33652 14424 33658
rect 14372 33594 14424 33600
rect 14464 33652 14516 33658
rect 14464 33594 14516 33600
rect 14372 33516 14424 33522
rect 14372 33458 14424 33464
rect 14280 32972 14332 32978
rect 14280 32914 14332 32920
rect 14186 32056 14242 32065
rect 14186 31991 14242 32000
rect 14004 31884 14056 31890
rect 14004 31826 14056 31832
rect 13912 31748 13964 31754
rect 13740 31708 13860 31736
rect 13832 31657 13860 31708
rect 13912 31690 13964 31696
rect 13818 31648 13874 31657
rect 13818 31583 13874 31592
rect 13924 31210 13952 31690
rect 13912 31204 13964 31210
rect 13912 31146 13964 31152
rect 13910 30832 13966 30841
rect 13910 30767 13966 30776
rect 13818 30016 13874 30025
rect 13818 29951 13874 29960
rect 13832 29238 13860 29951
rect 13820 29232 13872 29238
rect 13820 29174 13872 29180
rect 13634 29064 13690 29073
rect 13634 28999 13690 29008
rect 13544 28688 13596 28694
rect 13544 28630 13596 28636
rect 13636 28484 13688 28490
rect 13636 28426 13688 28432
rect 13648 28150 13676 28426
rect 13636 28144 13688 28150
rect 13636 28086 13688 28092
rect 13452 26988 13504 26994
rect 13452 26930 13504 26936
rect 13084 24744 13136 24750
rect 13084 24686 13136 24692
rect 13268 24744 13320 24750
rect 13268 24686 13320 24692
rect 12992 24676 13044 24682
rect 12992 24618 13044 24624
rect 13176 24676 13228 24682
rect 13176 24618 13228 24624
rect 13188 24342 13216 24618
rect 13360 24608 13412 24614
rect 13360 24550 13412 24556
rect 13176 24336 13228 24342
rect 13176 24278 13228 24284
rect 13372 24274 13400 24550
rect 12532 24268 12584 24274
rect 12532 24210 12584 24216
rect 13360 24268 13412 24274
rect 13360 24210 13412 24216
rect 12256 24200 12308 24206
rect 12256 24142 12308 24148
rect 12268 23730 12296 24142
rect 13360 23860 13412 23866
rect 13360 23802 13412 23808
rect 12256 23724 12308 23730
rect 12256 23666 12308 23672
rect 13372 23526 13400 23802
rect 13360 23520 13412 23526
rect 13360 23462 13412 23468
rect 12532 23112 12584 23118
rect 12532 23054 12584 23060
rect 12348 23044 12400 23050
rect 12348 22986 12400 22992
rect 12164 22432 12216 22438
rect 12164 22374 12216 22380
rect 12072 21956 12124 21962
rect 12072 21898 12124 21904
rect 11532 21814 11652 21842
rect 11244 21344 11296 21350
rect 11244 21286 11296 21292
rect 11256 20942 11284 21286
rect 11532 20942 11560 21814
rect 11612 21480 11664 21486
rect 11612 21422 11664 21428
rect 11624 21146 11652 21422
rect 11612 21140 11664 21146
rect 11612 21082 11664 21088
rect 11244 20936 11296 20942
rect 11244 20878 11296 20884
rect 11520 20936 11572 20942
rect 11520 20878 11572 20884
rect 11060 20596 11112 20602
rect 11060 20538 11112 20544
rect 10968 19780 11020 19786
rect 10968 19722 11020 19728
rect 11256 19718 11284 20878
rect 11532 20602 11560 20878
rect 12084 20806 12112 21898
rect 12176 21690 12204 22374
rect 12360 22166 12388 22986
rect 12348 22160 12400 22166
rect 12348 22102 12400 22108
rect 12164 21684 12216 21690
rect 12164 21626 12216 21632
rect 12072 20800 12124 20806
rect 12072 20742 12124 20748
rect 11520 20596 11572 20602
rect 11520 20538 11572 20544
rect 12176 20398 12204 21626
rect 12348 20596 12400 20602
rect 12348 20538 12400 20544
rect 12164 20392 12216 20398
rect 12164 20334 12216 20340
rect 12360 19990 12388 20538
rect 12440 20324 12492 20330
rect 12440 20266 12492 20272
rect 12348 19984 12400 19990
rect 12348 19926 12400 19932
rect 12452 19854 12480 20266
rect 12544 20058 12572 23054
rect 13360 22976 13412 22982
rect 13360 22918 13412 22924
rect 12624 22636 12676 22642
rect 12624 22578 12676 22584
rect 12636 22030 12664 22578
rect 13372 22098 13400 22918
rect 13360 22092 13412 22098
rect 13360 22034 13412 22040
rect 12624 22024 12676 22030
rect 12624 21966 12676 21972
rect 12532 20052 12584 20058
rect 12532 19994 12584 20000
rect 12440 19848 12492 19854
rect 12440 19790 12492 19796
rect 10600 19712 10652 19718
rect 10600 19654 10652 19660
rect 11244 19712 11296 19718
rect 11244 19654 11296 19660
rect 10612 19514 10640 19654
rect 10600 19508 10652 19514
rect 10600 19450 10652 19456
rect 11256 19446 11284 19654
rect 12452 19514 12480 19790
rect 12440 19508 12492 19514
rect 12440 19450 12492 19456
rect 11244 19440 11296 19446
rect 11244 19382 11296 19388
rect 12452 18970 12480 19450
rect 12440 18964 12492 18970
rect 12440 18906 12492 18912
rect 10876 11076 10928 11082
rect 10876 11018 10928 11024
rect 10508 7336 10560 7342
rect 10508 7278 10560 7284
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 8576 2848 8628 2854
rect 8576 2790 8628 2796
rect 8588 2446 8616 2790
rect 8680 2650 8708 2994
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 10888 2446 10916 11018
rect 12636 10810 12664 21966
rect 13268 21548 13320 21554
rect 13268 21490 13320 21496
rect 12808 21480 12860 21486
rect 12808 21422 12860 21428
rect 12820 21010 12848 21422
rect 12808 21004 12860 21010
rect 12808 20946 12860 20952
rect 13084 20936 13136 20942
rect 13084 20878 13136 20884
rect 12716 20800 12768 20806
rect 12716 20742 12768 20748
rect 12728 19786 12756 20742
rect 13096 20058 13124 20878
rect 13084 20052 13136 20058
rect 13084 19994 13136 20000
rect 12716 19780 12768 19786
rect 12716 19722 12768 19728
rect 12728 19514 12756 19722
rect 12716 19508 12768 19514
rect 12716 19450 12768 19456
rect 13280 19310 13308 21490
rect 13464 21434 13492 26930
rect 13636 26784 13688 26790
rect 13636 26726 13688 26732
rect 13648 25906 13676 26726
rect 13728 26580 13780 26586
rect 13728 26522 13780 26528
rect 13740 26042 13768 26522
rect 13924 26246 13952 30767
rect 13912 26240 13964 26246
rect 13912 26182 13964 26188
rect 13728 26036 13780 26042
rect 13728 25978 13780 25984
rect 13912 26036 13964 26042
rect 13912 25978 13964 25984
rect 13636 25900 13688 25906
rect 13636 25842 13688 25848
rect 13544 25832 13596 25838
rect 13544 25774 13596 25780
rect 13556 25430 13584 25774
rect 13648 25430 13676 25842
rect 13924 25838 13952 25978
rect 13912 25832 13964 25838
rect 13912 25774 13964 25780
rect 14016 25786 14044 31826
rect 14200 31686 14228 31991
rect 14292 31929 14320 32914
rect 14278 31920 14334 31929
rect 14278 31855 14334 31864
rect 14188 31680 14240 31686
rect 14188 31622 14240 31628
rect 14280 31340 14332 31346
rect 14280 31282 14332 31288
rect 14292 30734 14320 31282
rect 14280 30728 14332 30734
rect 14280 30670 14332 30676
rect 14188 30592 14240 30598
rect 14188 30534 14240 30540
rect 14280 30592 14332 30598
rect 14280 30534 14332 30540
rect 14096 30184 14148 30190
rect 14096 30126 14148 30132
rect 14108 29345 14136 30126
rect 14094 29336 14150 29345
rect 14094 29271 14150 29280
rect 14200 29238 14228 30534
rect 14188 29232 14240 29238
rect 14188 29174 14240 29180
rect 14108 29102 14136 29133
rect 14096 29096 14148 29102
rect 14094 29064 14096 29073
rect 14148 29064 14150 29073
rect 14094 28999 14150 29008
rect 14108 26926 14136 28999
rect 14292 28150 14320 30534
rect 14280 28144 14332 28150
rect 14280 28086 14332 28092
rect 14384 27962 14412 33458
rect 14476 33318 14504 33594
rect 14464 33312 14516 33318
rect 14464 33254 14516 33260
rect 14464 29776 14516 29782
rect 14464 29718 14516 29724
rect 14476 28150 14504 29718
rect 14568 29578 14596 34478
rect 14646 34096 14702 34105
rect 14646 34031 14702 34040
rect 14660 32910 14688 34031
rect 15028 33930 15056 34886
rect 15120 34746 15148 35702
rect 15384 35080 15436 35086
rect 15384 35022 15436 35028
rect 15198 34912 15254 34921
rect 15198 34847 15254 34856
rect 15108 34740 15160 34746
rect 15108 34682 15160 34688
rect 15212 34406 15240 34847
rect 15292 34604 15344 34610
rect 15292 34546 15344 34552
rect 15200 34400 15252 34406
rect 15200 34342 15252 34348
rect 15200 33992 15252 33998
rect 15200 33934 15252 33940
rect 14924 33924 14976 33930
rect 14924 33866 14976 33872
rect 15016 33924 15068 33930
rect 15016 33866 15068 33872
rect 14740 33312 14792 33318
rect 14740 33254 14792 33260
rect 14648 32904 14700 32910
rect 14648 32846 14700 32852
rect 14752 32842 14780 33254
rect 14740 32836 14792 32842
rect 14792 32796 14872 32824
rect 14740 32778 14792 32784
rect 14648 31884 14700 31890
rect 14648 31826 14700 31832
rect 14556 29572 14608 29578
rect 14556 29514 14608 29520
rect 14660 29034 14688 31826
rect 14844 30122 14872 32796
rect 14936 30326 14964 33866
rect 15028 31278 15056 33866
rect 15108 32496 15160 32502
rect 15108 32438 15160 32444
rect 15120 32201 15148 32438
rect 15212 32366 15240 33934
rect 15200 32360 15252 32366
rect 15200 32302 15252 32308
rect 15106 32192 15162 32201
rect 15106 32127 15162 32136
rect 15304 31521 15332 34546
rect 15396 34406 15424 35022
rect 15384 34400 15436 34406
rect 15384 34342 15436 34348
rect 15396 33289 15424 34342
rect 15382 33280 15438 33289
rect 15382 33215 15438 33224
rect 15384 32564 15436 32570
rect 15384 32506 15436 32512
rect 15396 32026 15424 32506
rect 15384 32020 15436 32026
rect 15384 31962 15436 31968
rect 15396 31890 15424 31962
rect 15384 31884 15436 31890
rect 15384 31826 15436 31832
rect 15290 31512 15346 31521
rect 15120 31470 15290 31498
rect 15016 31272 15068 31278
rect 15016 31214 15068 31220
rect 15028 30802 15056 31214
rect 15016 30796 15068 30802
rect 15016 30738 15068 30744
rect 15120 30716 15148 31470
rect 15290 31447 15346 31456
rect 15304 31387 15332 31447
rect 15200 31272 15252 31278
rect 15200 31214 15252 31220
rect 15212 30841 15240 31214
rect 15292 31136 15344 31142
rect 15292 31078 15344 31084
rect 15384 31136 15436 31142
rect 15384 31078 15436 31084
rect 15198 30832 15254 30841
rect 15198 30767 15254 30776
rect 15120 30688 15240 30716
rect 15016 30592 15068 30598
rect 15016 30534 15068 30540
rect 14924 30320 14976 30326
rect 14924 30262 14976 30268
rect 14832 30116 14884 30122
rect 14832 30058 14884 30064
rect 14740 30048 14792 30054
rect 14740 29990 14792 29996
rect 14752 29578 14780 29990
rect 14740 29572 14792 29578
rect 14740 29514 14792 29520
rect 14648 29028 14700 29034
rect 14648 28970 14700 28976
rect 14464 28144 14516 28150
rect 14464 28086 14516 28092
rect 14660 28014 14688 28970
rect 14844 28626 14872 30058
rect 14924 29572 14976 29578
rect 14924 29514 14976 29520
rect 14832 28620 14884 28626
rect 14832 28562 14884 28568
rect 14648 28008 14700 28014
rect 14384 27934 14504 27962
rect 14648 27950 14700 27956
rect 14372 27872 14424 27878
rect 14372 27814 14424 27820
rect 14384 27062 14412 27814
rect 14476 27690 14504 27934
rect 14554 27704 14610 27713
rect 14476 27662 14554 27690
rect 14554 27639 14610 27648
rect 14568 27470 14596 27639
rect 14660 27606 14688 27950
rect 14648 27600 14700 27606
rect 14648 27542 14700 27548
rect 14556 27464 14608 27470
rect 14556 27406 14608 27412
rect 14936 27062 14964 29514
rect 15028 28014 15056 30534
rect 15212 29481 15240 30688
rect 15304 30326 15332 31078
rect 15292 30320 15344 30326
rect 15292 30262 15344 30268
rect 15198 29472 15254 29481
rect 15198 29407 15254 29416
rect 15396 29238 15424 31078
rect 15488 29510 15516 35702
rect 15660 35148 15712 35154
rect 15660 35090 15712 35096
rect 15566 35048 15622 35057
rect 15566 34983 15622 34992
rect 15580 33386 15608 34983
rect 15672 34746 15700 35090
rect 15764 35057 15792 35799
rect 16132 35680 16160 36518
rect 16408 35698 16436 37334
rect 16500 37262 16528 37606
rect 16672 37324 16724 37330
rect 16672 37266 16724 37272
rect 16488 37256 16540 37262
rect 16488 37198 16540 37204
rect 16578 37224 16634 37233
rect 16578 37159 16634 37168
rect 16592 37126 16620 37159
rect 16580 37120 16632 37126
rect 16580 37062 16632 37068
rect 16684 36938 16712 37266
rect 16776 37126 16804 39200
rect 18050 37496 18106 37505
rect 18050 37431 18106 37440
rect 16856 37256 16908 37262
rect 16856 37198 16908 37204
rect 17132 37256 17184 37262
rect 17132 37198 17184 37204
rect 16764 37120 16816 37126
rect 16764 37062 16816 37068
rect 16592 36910 16712 36938
rect 16592 36038 16620 36910
rect 16672 36576 16724 36582
rect 16672 36518 16724 36524
rect 16580 36032 16632 36038
rect 16580 35974 16632 35980
rect 16684 35698 16712 36518
rect 16762 36272 16818 36281
rect 16762 36207 16818 36216
rect 16776 36174 16804 36207
rect 16764 36168 16816 36174
rect 16764 36110 16816 36116
rect 16396 35692 16448 35698
rect 16132 35652 16344 35680
rect 15750 35048 15806 35057
rect 16210 35048 16266 35057
rect 15750 34983 15806 34992
rect 15844 35012 15896 35018
rect 16210 34983 16266 34992
rect 15844 34954 15896 34960
rect 15660 34740 15712 34746
rect 15660 34682 15712 34688
rect 15660 34536 15712 34542
rect 15660 34478 15712 34484
rect 15752 34536 15804 34542
rect 15752 34478 15804 34484
rect 15568 33380 15620 33386
rect 15568 33322 15620 33328
rect 15566 32192 15622 32201
rect 15566 32127 15622 32136
rect 15580 32026 15608 32127
rect 15568 32020 15620 32026
rect 15568 31962 15620 31968
rect 15672 31754 15700 34478
rect 15764 31890 15792 34478
rect 15856 33930 15884 34954
rect 16028 34944 16080 34950
rect 16028 34886 16080 34892
rect 15844 33924 15896 33930
rect 15844 33866 15896 33872
rect 16040 33590 16068 34886
rect 16120 33924 16172 33930
rect 16120 33866 16172 33872
rect 15844 33584 15896 33590
rect 16028 33584 16080 33590
rect 15896 33544 15976 33572
rect 15844 33526 15896 33532
rect 15948 33454 15976 33544
rect 16028 33526 16080 33532
rect 15844 33448 15896 33454
rect 15844 33390 15896 33396
rect 15936 33448 15988 33454
rect 15936 33390 15988 33396
rect 15752 31884 15804 31890
rect 15752 31826 15804 31832
rect 15660 31748 15712 31754
rect 15660 31690 15712 31696
rect 15856 31278 15884 33390
rect 16132 32978 16160 33866
rect 16120 32972 16172 32978
rect 16120 32914 16172 32920
rect 16026 32192 16082 32201
rect 16026 32127 16082 32136
rect 16040 31958 16068 32127
rect 16028 31952 16080 31958
rect 16028 31894 16080 31900
rect 16028 31340 16080 31346
rect 16028 31282 16080 31288
rect 15844 31272 15896 31278
rect 15844 31214 15896 31220
rect 15844 30660 15896 30666
rect 15844 30602 15896 30608
rect 15566 29744 15622 29753
rect 15566 29679 15568 29688
rect 15620 29679 15622 29688
rect 15568 29650 15620 29656
rect 15476 29504 15528 29510
rect 15476 29446 15528 29452
rect 15384 29232 15436 29238
rect 15384 29174 15436 29180
rect 15292 29096 15344 29102
rect 15292 29038 15344 29044
rect 15016 28008 15068 28014
rect 15016 27950 15068 27956
rect 15200 27872 15252 27878
rect 15200 27814 15252 27820
rect 15212 27418 15240 27814
rect 15120 27402 15240 27418
rect 15108 27396 15240 27402
rect 15160 27390 15240 27396
rect 15108 27338 15160 27344
rect 14372 27056 14424 27062
rect 14372 26998 14424 27004
rect 14924 27056 14976 27062
rect 14924 26998 14976 27004
rect 15108 27056 15160 27062
rect 15108 26998 15160 27004
rect 14096 26920 14148 26926
rect 14096 26862 14148 26868
rect 14108 25974 14136 26862
rect 14936 26450 14964 26998
rect 15120 26586 15148 26998
rect 15108 26580 15160 26586
rect 15108 26522 15160 26528
rect 14924 26444 14976 26450
rect 14924 26386 14976 26392
rect 14556 26308 14608 26314
rect 14556 26250 14608 26256
rect 14096 25968 14148 25974
rect 14096 25910 14148 25916
rect 14188 25832 14240 25838
rect 14016 25758 14136 25786
rect 14188 25774 14240 25780
rect 13728 25696 13780 25702
rect 13728 25638 13780 25644
rect 13820 25696 13872 25702
rect 13820 25638 13872 25644
rect 13544 25424 13596 25430
rect 13544 25366 13596 25372
rect 13636 25424 13688 25430
rect 13636 25366 13688 25372
rect 13648 25294 13676 25366
rect 13636 25288 13688 25294
rect 13636 25230 13688 25236
rect 13740 24614 13768 25638
rect 13832 25362 13860 25638
rect 13820 25356 13872 25362
rect 13820 25298 13872 25304
rect 13820 25152 13872 25158
rect 13820 25094 13872 25100
rect 13544 24608 13596 24614
rect 13544 24550 13596 24556
rect 13728 24608 13780 24614
rect 13728 24550 13780 24556
rect 13556 23798 13584 24550
rect 13832 24410 13860 25094
rect 14004 24608 14056 24614
rect 14004 24550 14056 24556
rect 14016 24410 14044 24550
rect 13820 24404 13872 24410
rect 13820 24346 13872 24352
rect 14004 24404 14056 24410
rect 14004 24346 14056 24352
rect 13636 24200 13688 24206
rect 13636 24142 13688 24148
rect 13544 23792 13596 23798
rect 13544 23734 13596 23740
rect 13648 23526 13676 24142
rect 13832 23662 13860 24346
rect 14004 23724 14056 23730
rect 14004 23666 14056 23672
rect 13820 23656 13872 23662
rect 13820 23598 13872 23604
rect 13636 23520 13688 23526
rect 13636 23462 13688 23468
rect 13544 22568 13596 22574
rect 13544 22510 13596 22516
rect 13556 21894 13584 22510
rect 13544 21888 13596 21894
rect 13544 21830 13596 21836
rect 13372 21406 13492 21434
rect 13268 19304 13320 19310
rect 13268 19246 13320 19252
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12728 3194 12756 10406
rect 13372 8974 13400 21406
rect 13556 20806 13584 21830
rect 13544 20800 13596 20806
rect 13544 20742 13596 20748
rect 13556 20398 13584 20742
rect 13544 20392 13596 20398
rect 13544 20334 13596 20340
rect 13360 8968 13412 8974
rect 13360 8910 13412 8916
rect 13648 8838 13676 23462
rect 13832 22098 13860 23598
rect 14016 23118 14044 23666
rect 14004 23112 14056 23118
rect 14004 23054 14056 23060
rect 14108 23050 14136 25758
rect 14200 24954 14228 25774
rect 14464 25764 14516 25770
rect 14464 25706 14516 25712
rect 14476 25226 14504 25706
rect 14372 25220 14424 25226
rect 14372 25162 14424 25168
rect 14464 25220 14516 25226
rect 14464 25162 14516 25168
rect 14188 24948 14240 24954
rect 14188 24890 14240 24896
rect 14384 24682 14412 25162
rect 14568 24818 14596 26250
rect 14648 26240 14700 26246
rect 14648 26182 14700 26188
rect 14556 24812 14608 24818
rect 14556 24754 14608 24760
rect 14372 24676 14424 24682
rect 14372 24618 14424 24624
rect 14660 24206 14688 26182
rect 14832 25900 14884 25906
rect 14832 25842 14884 25848
rect 14844 24954 14872 25842
rect 14936 25430 14964 26386
rect 14924 25424 14976 25430
rect 14924 25366 14976 25372
rect 14832 24948 14884 24954
rect 14832 24890 14884 24896
rect 14740 24812 14792 24818
rect 14740 24754 14792 24760
rect 14648 24200 14700 24206
rect 14648 24142 14700 24148
rect 14752 24070 14780 24754
rect 14740 24064 14792 24070
rect 14740 24006 14792 24012
rect 14372 23588 14424 23594
rect 14372 23530 14424 23536
rect 14384 23254 14412 23530
rect 14372 23248 14424 23254
rect 14372 23190 14424 23196
rect 14096 23044 14148 23050
rect 14096 22986 14148 22992
rect 14096 22568 14148 22574
rect 14096 22510 14148 22516
rect 13820 22092 13872 22098
rect 13820 22034 13872 22040
rect 14108 21622 14136 22510
rect 14384 22506 14412 23190
rect 14752 22642 14780 24006
rect 14740 22636 14792 22642
rect 14740 22578 14792 22584
rect 14372 22500 14424 22506
rect 14372 22442 14424 22448
rect 13912 21616 13964 21622
rect 13912 21558 13964 21564
rect 14096 21616 14148 21622
rect 14096 21558 14148 21564
rect 13924 21010 13952 21558
rect 13912 21004 13964 21010
rect 13912 20946 13964 20952
rect 13924 20330 13952 20946
rect 13912 20324 13964 20330
rect 13912 20266 13964 20272
rect 14280 19712 14332 19718
rect 14280 19654 14332 19660
rect 14292 18290 14320 19654
rect 14280 18284 14332 18290
rect 14280 18226 14332 18232
rect 14384 10674 14412 22442
rect 14844 22094 14872 24890
rect 15120 24682 15148 26522
rect 15108 24676 15160 24682
rect 15108 24618 15160 24624
rect 14924 24132 14976 24138
rect 14924 24074 14976 24080
rect 14752 22066 14872 22094
rect 14752 19854 14780 22066
rect 14832 20868 14884 20874
rect 14832 20810 14884 20816
rect 14844 20602 14872 20810
rect 14832 20596 14884 20602
rect 14832 20538 14884 20544
rect 14832 20324 14884 20330
rect 14832 20266 14884 20272
rect 14844 19922 14872 20266
rect 14832 19916 14884 19922
rect 14832 19858 14884 19864
rect 14740 19848 14792 19854
rect 14740 19790 14792 19796
rect 14752 19378 14780 19790
rect 14740 19372 14792 19378
rect 14740 19314 14792 19320
rect 14372 10668 14424 10674
rect 14372 10610 14424 10616
rect 13636 8832 13688 8838
rect 13636 8774 13688 8780
rect 12716 3188 12768 3194
rect 12716 3130 12768 3136
rect 14936 3126 14964 24074
rect 15200 23588 15252 23594
rect 15200 23530 15252 23536
rect 15212 22506 15240 23530
rect 15200 22500 15252 22506
rect 15200 22442 15252 22448
rect 15304 22030 15332 29038
rect 15580 28694 15608 29650
rect 15856 29345 15884 30602
rect 15934 30560 15990 30569
rect 15934 30495 15990 30504
rect 15948 29782 15976 30495
rect 15936 29776 15988 29782
rect 15936 29718 15988 29724
rect 15842 29336 15898 29345
rect 15842 29271 15898 29280
rect 15568 28688 15620 28694
rect 15568 28630 15620 28636
rect 15568 27940 15620 27946
rect 15568 27882 15620 27888
rect 15384 26784 15436 26790
rect 15384 26726 15436 26732
rect 15396 26450 15424 26726
rect 15384 26444 15436 26450
rect 15384 26386 15436 26392
rect 15476 26240 15528 26246
rect 15476 26182 15528 26188
rect 15488 24886 15516 26182
rect 15580 25702 15608 27882
rect 15856 27538 15884 29271
rect 16040 28762 16068 31282
rect 16224 31226 16252 34983
rect 16132 31198 16252 31226
rect 16132 30598 16160 31198
rect 16212 31136 16264 31142
rect 16212 31078 16264 31084
rect 16224 30870 16252 31078
rect 16212 30864 16264 30870
rect 16212 30806 16264 30812
rect 16120 30592 16172 30598
rect 16120 30534 16172 30540
rect 16224 30274 16252 30806
rect 16316 30802 16344 35652
rect 16396 35634 16448 35640
rect 16672 35692 16724 35698
rect 16672 35634 16724 35640
rect 16580 35624 16632 35630
rect 16580 35566 16632 35572
rect 16486 35456 16542 35465
rect 16486 35391 16542 35400
rect 16396 35080 16448 35086
rect 16396 35022 16448 35028
rect 16408 34950 16436 35022
rect 16500 35018 16528 35391
rect 16488 35012 16540 35018
rect 16488 34954 16540 34960
rect 16396 34944 16448 34950
rect 16396 34886 16448 34892
rect 16408 33114 16436 34886
rect 16592 34649 16620 35566
rect 16776 35562 16804 36110
rect 16764 35556 16816 35562
rect 16764 35498 16816 35504
rect 16868 35086 16896 37198
rect 17040 36780 17092 36786
rect 17040 36722 17092 36728
rect 17052 36310 17080 36722
rect 17040 36304 17092 36310
rect 17040 36246 17092 36252
rect 16948 35692 17000 35698
rect 16948 35634 17000 35640
rect 16960 35465 16988 35634
rect 17040 35488 17092 35494
rect 16946 35456 17002 35465
rect 17040 35430 17092 35436
rect 16946 35391 17002 35400
rect 16856 35080 16908 35086
rect 16856 35022 16908 35028
rect 16578 34640 16634 34649
rect 16578 34575 16634 34584
rect 16856 34604 16908 34610
rect 16856 34546 16908 34552
rect 16488 34060 16540 34066
rect 16488 34002 16540 34008
rect 16500 33930 16528 34002
rect 16488 33924 16540 33930
rect 16488 33866 16540 33872
rect 16500 33318 16528 33866
rect 16672 33516 16724 33522
rect 16672 33458 16724 33464
rect 16488 33312 16540 33318
rect 16488 33254 16540 33260
rect 16396 33108 16448 33114
rect 16396 33050 16448 33056
rect 16580 33108 16632 33114
rect 16580 33050 16632 33056
rect 16592 32978 16620 33050
rect 16580 32972 16632 32978
rect 16580 32914 16632 32920
rect 16396 32836 16448 32842
rect 16396 32778 16448 32784
rect 16408 32586 16436 32778
rect 16580 32768 16632 32774
rect 16684 32756 16712 33458
rect 16764 32836 16816 32842
rect 16764 32778 16816 32784
rect 16632 32728 16712 32756
rect 16580 32710 16632 32716
rect 16776 32586 16804 32778
rect 16408 32558 16804 32586
rect 16868 32570 16896 34546
rect 16948 32972 17000 32978
rect 16948 32914 17000 32920
rect 16856 32564 16908 32570
rect 16856 32506 16908 32512
rect 16960 32337 16988 32914
rect 17052 32774 17080 35430
rect 17040 32768 17092 32774
rect 17040 32710 17092 32716
rect 16946 32328 17002 32337
rect 16946 32263 17002 32272
rect 16396 31952 16448 31958
rect 16396 31894 16448 31900
rect 16948 31952 17000 31958
rect 16948 31894 17000 31900
rect 16304 30796 16356 30802
rect 16304 30738 16356 30744
rect 16132 30246 16252 30274
rect 16132 30190 16160 30246
rect 16120 30184 16172 30190
rect 16120 30126 16172 30132
rect 16132 29238 16160 30126
rect 16120 29232 16172 29238
rect 16212 29232 16264 29238
rect 16120 29174 16172 29180
rect 16210 29200 16212 29209
rect 16264 29200 16266 29209
rect 16210 29135 16266 29144
rect 16408 29050 16436 31894
rect 16580 31884 16632 31890
rect 16580 31826 16632 31832
rect 16592 31754 16620 31826
rect 16960 31804 16988 31894
rect 16868 31776 16988 31804
rect 16592 31726 16712 31754
rect 16580 31680 16632 31686
rect 16580 31622 16632 31628
rect 16592 30190 16620 31622
rect 16580 30184 16632 30190
rect 16580 30126 16632 30132
rect 16488 30116 16540 30122
rect 16488 30058 16540 30064
rect 16500 29850 16528 30058
rect 16592 29850 16620 30126
rect 16488 29844 16540 29850
rect 16488 29786 16540 29792
rect 16580 29844 16632 29850
rect 16580 29786 16632 29792
rect 16132 29022 16436 29050
rect 16028 28756 16080 28762
rect 16028 28698 16080 28704
rect 15936 28688 15988 28694
rect 15936 28630 15988 28636
rect 15844 27532 15896 27538
rect 15844 27474 15896 27480
rect 15660 25900 15712 25906
rect 15660 25842 15712 25848
rect 15672 25702 15700 25842
rect 15568 25696 15620 25702
rect 15568 25638 15620 25644
rect 15660 25696 15712 25702
rect 15660 25638 15712 25644
rect 15476 24880 15528 24886
rect 15476 24822 15528 24828
rect 15580 24342 15608 25638
rect 15672 24834 15700 25638
rect 15844 25152 15896 25158
rect 15844 25094 15896 25100
rect 15856 24886 15884 25094
rect 15844 24880 15896 24886
rect 15672 24806 15792 24834
rect 15844 24822 15896 24828
rect 15660 24744 15712 24750
rect 15660 24686 15712 24692
rect 15568 24336 15620 24342
rect 15568 24278 15620 24284
rect 15672 24274 15700 24686
rect 15764 24290 15792 24806
rect 15660 24268 15712 24274
rect 15764 24262 15884 24290
rect 15660 24210 15712 24216
rect 15752 24132 15804 24138
rect 15752 24074 15804 24080
rect 15764 23866 15792 24074
rect 15568 23860 15620 23866
rect 15568 23802 15620 23808
rect 15752 23860 15804 23866
rect 15752 23802 15804 23808
rect 15580 23746 15608 23802
rect 15856 23746 15884 24262
rect 15580 23718 15884 23746
rect 15384 23520 15436 23526
rect 15384 23462 15436 23468
rect 15396 22642 15424 23462
rect 15568 23044 15620 23050
rect 15568 22986 15620 22992
rect 15384 22636 15436 22642
rect 15384 22578 15436 22584
rect 15580 22506 15608 22986
rect 15568 22500 15620 22506
rect 15568 22442 15620 22448
rect 15292 22024 15344 22030
rect 15292 21966 15344 21972
rect 15292 21548 15344 21554
rect 15292 21490 15344 21496
rect 15108 21344 15160 21350
rect 15108 21286 15160 21292
rect 15016 20392 15068 20398
rect 15016 20334 15068 20340
rect 15028 19514 15056 20334
rect 15120 19718 15148 21286
rect 15108 19712 15160 19718
rect 15108 19654 15160 19660
rect 15016 19508 15068 19514
rect 15016 19450 15068 19456
rect 15200 19304 15252 19310
rect 15200 19246 15252 19252
rect 15212 6914 15240 19246
rect 15304 19242 15332 21490
rect 15384 21480 15436 21486
rect 15384 21422 15436 21428
rect 15396 20874 15424 21422
rect 15580 21418 15608 22442
rect 15856 22094 15884 23718
rect 15764 22066 15884 22094
rect 15660 21888 15712 21894
rect 15660 21830 15712 21836
rect 15672 21554 15700 21830
rect 15660 21548 15712 21554
rect 15660 21490 15712 21496
rect 15568 21412 15620 21418
rect 15568 21354 15620 21360
rect 15476 21004 15528 21010
rect 15476 20946 15528 20952
rect 15384 20868 15436 20874
rect 15384 20810 15436 20816
rect 15292 19236 15344 19242
rect 15292 19178 15344 19184
rect 15396 12442 15424 20810
rect 15488 20466 15516 20946
rect 15568 20800 15620 20806
rect 15568 20742 15620 20748
rect 15476 20460 15528 20466
rect 15476 20402 15528 20408
rect 15384 12436 15436 12442
rect 15384 12378 15436 12384
rect 15212 6886 15424 6914
rect 14924 3120 14976 3126
rect 14924 3062 14976 3068
rect 11978 2680 12034 2689
rect 11978 2615 12034 2624
rect 11992 2582 12020 2615
rect 11980 2576 12032 2582
rect 11980 2518 12032 2524
rect 15396 2514 15424 6886
rect 15580 2990 15608 20742
rect 15764 6914 15792 22066
rect 15672 6886 15792 6914
rect 15568 2984 15620 2990
rect 15568 2926 15620 2932
rect 15672 2582 15700 6886
rect 15948 3194 15976 28630
rect 16040 28082 16068 28698
rect 16132 28626 16160 29022
rect 16212 28960 16264 28966
rect 16212 28902 16264 28908
rect 16120 28620 16172 28626
rect 16120 28562 16172 28568
rect 16028 28076 16080 28082
rect 16028 28018 16080 28024
rect 16132 27130 16160 28562
rect 16224 28490 16252 28902
rect 16684 28778 16712 31726
rect 16764 31748 16816 31754
rect 16868 31736 16896 31776
rect 16816 31708 16896 31736
rect 16764 31690 16816 31696
rect 17038 31648 17094 31657
rect 17038 31583 17094 31592
rect 16764 30660 16816 30666
rect 16816 30620 16896 30648
rect 16764 30602 16816 30608
rect 16684 28750 16804 28778
rect 16868 28762 16896 30620
rect 17052 30326 17080 31583
rect 17040 30320 17092 30326
rect 17040 30262 17092 30268
rect 16948 30184 17000 30190
rect 16948 30126 17000 30132
rect 16960 29306 16988 30126
rect 16948 29300 17000 29306
rect 16948 29242 17000 29248
rect 16672 28688 16724 28694
rect 16672 28630 16724 28636
rect 16212 28484 16264 28490
rect 16212 28426 16264 28432
rect 16396 28416 16448 28422
rect 16396 28358 16448 28364
rect 16408 28218 16436 28358
rect 16396 28212 16448 28218
rect 16396 28154 16448 28160
rect 16580 28144 16632 28150
rect 16580 28086 16632 28092
rect 16488 28076 16540 28082
rect 16488 28018 16540 28024
rect 16500 27538 16528 28018
rect 16488 27532 16540 27538
rect 16488 27474 16540 27480
rect 16592 27130 16620 28086
rect 16684 27402 16712 28630
rect 16672 27396 16724 27402
rect 16672 27338 16724 27344
rect 16120 27124 16172 27130
rect 16120 27066 16172 27072
rect 16580 27124 16632 27130
rect 16580 27066 16632 27072
rect 16120 26988 16172 26994
rect 16120 26930 16172 26936
rect 16132 26790 16160 26930
rect 16120 26784 16172 26790
rect 16120 26726 16172 26732
rect 16132 23769 16160 26726
rect 16396 26512 16448 26518
rect 16396 26454 16448 26460
rect 16304 26240 16356 26246
rect 16304 26182 16356 26188
rect 16316 25906 16344 26182
rect 16304 25900 16356 25906
rect 16304 25842 16356 25848
rect 16408 25294 16436 26454
rect 16396 25288 16448 25294
rect 16396 25230 16448 25236
rect 16776 24274 16804 28750
rect 16856 28756 16908 28762
rect 16856 28698 16908 28704
rect 17040 28756 17092 28762
rect 17040 28698 17092 28704
rect 16948 28620 17000 28626
rect 16948 28562 17000 28568
rect 16960 28014 16988 28562
rect 16948 28008 17000 28014
rect 16948 27950 17000 27956
rect 16856 27940 16908 27946
rect 16856 27882 16908 27888
rect 16868 27674 16896 27882
rect 16856 27668 16908 27674
rect 16856 27610 16908 27616
rect 16856 27396 16908 27402
rect 16856 27338 16908 27344
rect 16868 25922 16896 27338
rect 16948 27328 17000 27334
rect 16948 27270 17000 27276
rect 16960 26382 16988 27270
rect 17052 26466 17080 28698
rect 17144 26586 17172 37198
rect 17684 37120 17736 37126
rect 17314 37088 17370 37097
rect 17684 37062 17736 37068
rect 17314 37023 17370 37032
rect 17224 36916 17276 36922
rect 17224 36858 17276 36864
rect 17236 36718 17264 36858
rect 17224 36712 17276 36718
rect 17224 36654 17276 36660
rect 17328 36553 17356 37023
rect 17500 36780 17552 36786
rect 17500 36722 17552 36728
rect 17314 36544 17370 36553
rect 17314 36479 17370 36488
rect 17222 36272 17278 36281
rect 17222 36207 17278 36216
rect 17236 36174 17264 36207
rect 17224 36168 17276 36174
rect 17224 36110 17276 36116
rect 17236 34105 17264 36110
rect 17408 36032 17460 36038
rect 17408 35974 17460 35980
rect 17314 35728 17370 35737
rect 17314 35663 17370 35672
rect 17328 35465 17356 35663
rect 17314 35456 17370 35465
rect 17314 35391 17370 35400
rect 17316 35080 17368 35086
rect 17316 35022 17368 35028
rect 17222 34096 17278 34105
rect 17222 34031 17278 34040
rect 17224 33992 17276 33998
rect 17224 33934 17276 33940
rect 17236 33862 17264 33934
rect 17224 33856 17276 33862
rect 17224 33798 17276 33804
rect 17224 32972 17276 32978
rect 17224 32914 17276 32920
rect 17236 32473 17264 32914
rect 17222 32464 17278 32473
rect 17222 32399 17278 32408
rect 17328 31414 17356 35022
rect 17420 34678 17448 35974
rect 17408 34672 17460 34678
rect 17408 34614 17460 34620
rect 17512 34218 17540 36722
rect 17696 34678 17724 37062
rect 17868 36780 17920 36786
rect 17868 36722 17920 36728
rect 17880 36174 17908 36722
rect 17868 36168 17920 36174
rect 17868 36110 17920 36116
rect 17880 34921 17908 36110
rect 18064 36038 18092 37431
rect 18708 37126 18736 39200
rect 18880 37664 18932 37670
rect 18880 37606 18932 37612
rect 18696 37120 18748 37126
rect 18696 37062 18748 37068
rect 18604 36576 18656 36582
rect 18604 36518 18656 36524
rect 18616 36417 18644 36518
rect 18602 36408 18658 36417
rect 18602 36343 18658 36352
rect 18788 36100 18840 36106
rect 18788 36042 18840 36048
rect 17960 36032 18012 36038
rect 17960 35974 18012 35980
rect 18052 36032 18104 36038
rect 18052 35974 18104 35980
rect 17866 34912 17922 34921
rect 17866 34847 17922 34856
rect 17866 34776 17922 34785
rect 17866 34711 17922 34720
rect 17880 34678 17908 34711
rect 17684 34672 17736 34678
rect 17684 34614 17736 34620
rect 17868 34672 17920 34678
rect 17868 34614 17920 34620
rect 17512 34190 17816 34218
rect 17500 33924 17552 33930
rect 17500 33866 17552 33872
rect 17512 33590 17540 33866
rect 17684 33856 17736 33862
rect 17684 33798 17736 33804
rect 17500 33584 17552 33590
rect 17500 33526 17552 33532
rect 17408 33108 17460 33114
rect 17408 33050 17460 33056
rect 17316 31408 17368 31414
rect 17316 31350 17368 31356
rect 17224 31272 17276 31278
rect 17224 31214 17276 31220
rect 17236 26926 17264 31214
rect 17420 30190 17448 33050
rect 17512 32366 17540 33526
rect 17500 32360 17552 32366
rect 17500 32302 17552 32308
rect 17592 31884 17644 31890
rect 17592 31826 17644 31832
rect 17604 31754 17632 31826
rect 17696 31754 17724 33798
rect 17592 31748 17644 31754
rect 17592 31690 17644 31696
rect 17684 31748 17736 31754
rect 17684 31690 17736 31696
rect 17500 31680 17552 31686
rect 17500 31622 17552 31628
rect 17408 30184 17460 30190
rect 17408 30126 17460 30132
rect 17316 29640 17368 29646
rect 17512 29617 17540 31622
rect 17592 30660 17644 30666
rect 17592 30602 17644 30608
rect 17316 29582 17368 29588
rect 17498 29608 17554 29617
rect 17328 29102 17356 29582
rect 17498 29543 17554 29552
rect 17500 29504 17552 29510
rect 17500 29446 17552 29452
rect 17512 29238 17540 29446
rect 17604 29238 17632 30602
rect 17500 29232 17552 29238
rect 17500 29174 17552 29180
rect 17592 29232 17644 29238
rect 17592 29174 17644 29180
rect 17316 29096 17368 29102
rect 17316 29038 17368 29044
rect 17316 28756 17368 28762
rect 17316 28698 17368 28704
rect 17328 27713 17356 28698
rect 17314 27704 17370 27713
rect 17314 27639 17370 27648
rect 17224 26920 17276 26926
rect 17224 26862 17276 26868
rect 17132 26580 17184 26586
rect 17132 26522 17184 26528
rect 17224 26580 17276 26586
rect 17224 26522 17276 26528
rect 17236 26466 17264 26522
rect 17052 26438 17264 26466
rect 17498 26480 17554 26489
rect 17498 26415 17554 26424
rect 17512 26382 17540 26415
rect 16948 26376 17000 26382
rect 16948 26318 17000 26324
rect 17500 26376 17552 26382
rect 17500 26318 17552 26324
rect 16868 25894 16988 25922
rect 17512 25906 17540 26318
rect 16856 24744 16908 24750
rect 16856 24686 16908 24692
rect 16764 24268 16816 24274
rect 16764 24210 16816 24216
rect 16580 24064 16632 24070
rect 16580 24006 16632 24012
rect 16118 23760 16174 23769
rect 16118 23695 16174 23704
rect 16028 23044 16080 23050
rect 16028 22986 16080 22992
rect 16488 23044 16540 23050
rect 16592 23032 16620 24006
rect 16776 23186 16804 24210
rect 16868 23662 16896 24686
rect 16856 23656 16908 23662
rect 16856 23598 16908 23604
rect 16764 23180 16816 23186
rect 16764 23122 16816 23128
rect 16540 23004 16620 23032
rect 16488 22986 16540 22992
rect 16040 21486 16068 22986
rect 16776 22506 16804 23122
rect 16764 22500 16816 22506
rect 16764 22442 16816 22448
rect 16960 22094 16988 25894
rect 17500 25900 17552 25906
rect 17420 25860 17500 25888
rect 17040 25764 17092 25770
rect 17040 25706 17092 25712
rect 17052 25294 17080 25706
rect 17040 25288 17092 25294
rect 17040 25230 17092 25236
rect 17420 24818 17448 25860
rect 17500 25842 17552 25848
rect 17500 25356 17552 25362
rect 17500 25298 17552 25304
rect 17408 24812 17460 24818
rect 17408 24754 17460 24760
rect 17512 24410 17540 25298
rect 17040 24404 17092 24410
rect 17040 24346 17092 24352
rect 17500 24404 17552 24410
rect 17500 24346 17552 24352
rect 17052 23866 17080 24346
rect 17040 23860 17092 23866
rect 17040 23802 17092 23808
rect 17052 23730 17080 23802
rect 17040 23724 17092 23730
rect 17040 23666 17092 23672
rect 17604 23526 17632 29174
rect 17684 27396 17736 27402
rect 17684 27338 17736 27344
rect 17696 26994 17724 27338
rect 17684 26988 17736 26994
rect 17684 26930 17736 26936
rect 17788 25498 17816 34190
rect 17868 33992 17920 33998
rect 17868 33934 17920 33940
rect 17880 33590 17908 33934
rect 17972 33930 18000 35974
rect 18236 35488 18288 35494
rect 18236 35430 18288 35436
rect 18052 35012 18104 35018
rect 18052 34954 18104 34960
rect 17960 33924 18012 33930
rect 17960 33866 18012 33872
rect 17958 33824 18014 33833
rect 17958 33759 18014 33768
rect 17868 33584 17920 33590
rect 17868 33526 17920 33532
rect 17972 33522 18000 33759
rect 17960 33516 18012 33522
rect 17960 33458 18012 33464
rect 17868 33312 17920 33318
rect 17868 33254 17920 33260
rect 17880 30666 17908 33254
rect 18064 32745 18092 34954
rect 18248 33930 18276 35430
rect 18696 35080 18748 35086
rect 18696 35022 18748 35028
rect 18326 34232 18382 34241
rect 18326 34167 18382 34176
rect 18144 33924 18196 33930
rect 18144 33866 18196 33872
rect 18236 33924 18288 33930
rect 18236 33866 18288 33872
rect 18050 32736 18106 32745
rect 18050 32671 18106 32680
rect 17958 32600 18014 32609
rect 17958 32535 18014 32544
rect 17972 32366 18000 32535
rect 17960 32360 18012 32366
rect 17960 32302 18012 32308
rect 17958 31920 18014 31929
rect 17958 31855 17960 31864
rect 18012 31855 18014 31864
rect 17960 31826 18012 31832
rect 17960 30864 18012 30870
rect 17960 30806 18012 30812
rect 17868 30660 17920 30666
rect 17868 30602 17920 30608
rect 17868 30184 17920 30190
rect 17868 30126 17920 30132
rect 17880 30025 17908 30126
rect 17866 30016 17922 30025
rect 17866 29951 17922 29960
rect 17868 29096 17920 29102
rect 17868 29038 17920 29044
rect 17880 26858 17908 29038
rect 17972 27062 18000 30806
rect 17960 27056 18012 27062
rect 17960 26998 18012 27004
rect 17868 26852 17920 26858
rect 17868 26794 17920 26800
rect 17776 25492 17828 25498
rect 17776 25434 17828 25440
rect 17684 25288 17736 25294
rect 17684 25230 17736 25236
rect 17696 24614 17724 25230
rect 17880 25158 17908 26794
rect 17960 26308 18012 26314
rect 17960 26250 18012 26256
rect 17972 25906 18000 26250
rect 17960 25900 18012 25906
rect 17960 25842 18012 25848
rect 17868 25152 17920 25158
rect 17868 25094 17920 25100
rect 17868 24744 17920 24750
rect 17868 24686 17920 24692
rect 17684 24608 17736 24614
rect 17684 24550 17736 24556
rect 17592 23520 17644 23526
rect 17592 23462 17644 23468
rect 17696 23322 17724 24550
rect 17880 24274 17908 24686
rect 18064 24410 18092 32671
rect 18156 31142 18184 33866
rect 18340 32910 18368 34167
rect 18604 33312 18656 33318
rect 18604 33254 18656 33260
rect 18328 32904 18380 32910
rect 18328 32846 18380 32852
rect 18512 32768 18564 32774
rect 18512 32710 18564 32716
rect 18328 32496 18380 32502
rect 18328 32438 18380 32444
rect 18340 32201 18368 32438
rect 18420 32292 18472 32298
rect 18420 32234 18472 32240
rect 18326 32192 18382 32201
rect 18326 32127 18382 32136
rect 18432 31754 18460 32234
rect 18236 31748 18288 31754
rect 18236 31690 18288 31696
rect 18340 31726 18460 31754
rect 18248 31414 18276 31690
rect 18236 31408 18288 31414
rect 18236 31350 18288 31356
rect 18144 31136 18196 31142
rect 18144 31078 18196 31084
rect 18340 30546 18368 31726
rect 18524 31414 18552 32710
rect 18512 31408 18564 31414
rect 18512 31350 18564 31356
rect 18418 31240 18474 31249
rect 18418 31175 18474 31184
rect 18432 30734 18460 31175
rect 18420 30728 18472 30734
rect 18420 30670 18472 30676
rect 18340 30518 18460 30546
rect 18236 30048 18288 30054
rect 18236 29990 18288 29996
rect 18248 29578 18276 29990
rect 18432 29578 18460 30518
rect 18144 29572 18196 29578
rect 18144 29514 18196 29520
rect 18236 29572 18288 29578
rect 18236 29514 18288 29520
rect 18420 29572 18472 29578
rect 18420 29514 18472 29520
rect 18156 28218 18184 29514
rect 18236 29096 18288 29102
rect 18236 29038 18288 29044
rect 18512 29096 18564 29102
rect 18512 29038 18564 29044
rect 18248 28422 18276 29038
rect 18524 28490 18552 29038
rect 18512 28484 18564 28490
rect 18512 28426 18564 28432
rect 18236 28416 18288 28422
rect 18236 28358 18288 28364
rect 18420 28416 18472 28422
rect 18420 28358 18472 28364
rect 18144 28212 18196 28218
rect 18144 28154 18196 28160
rect 18156 26450 18184 28154
rect 18432 27826 18460 28358
rect 18524 27946 18552 28426
rect 18616 28150 18644 33254
rect 18708 32502 18736 35022
rect 18800 33930 18828 36042
rect 18892 35630 18920 37606
rect 19248 37324 19300 37330
rect 19248 37266 19300 37272
rect 18972 36780 19024 36786
rect 18972 36722 19024 36728
rect 18984 36174 19012 36722
rect 19156 36576 19208 36582
rect 19156 36518 19208 36524
rect 19062 36272 19118 36281
rect 19062 36207 19064 36216
rect 19116 36207 19118 36216
rect 19064 36178 19116 36184
rect 18972 36168 19024 36174
rect 18972 36110 19024 36116
rect 18880 35624 18932 35630
rect 18880 35566 18932 35572
rect 18984 34610 19012 36110
rect 19064 35216 19116 35222
rect 19064 35158 19116 35164
rect 19076 35018 19104 35158
rect 19064 35012 19116 35018
rect 19064 34954 19116 34960
rect 18972 34604 19024 34610
rect 18972 34546 19024 34552
rect 18788 33924 18840 33930
rect 18788 33866 18840 33872
rect 18800 32502 18828 33866
rect 18984 33522 19012 34546
rect 18972 33516 19024 33522
rect 18972 33458 19024 33464
rect 18696 32496 18748 32502
rect 18696 32438 18748 32444
rect 18788 32496 18840 32502
rect 18788 32438 18840 32444
rect 18788 31816 18840 31822
rect 18788 31758 18840 31764
rect 18800 30433 18828 31758
rect 19168 31482 19196 36518
rect 19260 34746 19288 37266
rect 19432 37256 19484 37262
rect 19432 37198 19484 37204
rect 19984 37256 20036 37262
rect 20640 37244 20668 39200
rect 21548 37732 21600 37738
rect 21548 37674 21600 37680
rect 21560 37398 21588 37674
rect 21548 37392 21600 37398
rect 21548 37334 21600 37340
rect 20720 37256 20772 37262
rect 20640 37216 20720 37244
rect 19984 37198 20036 37204
rect 20720 37198 20772 37204
rect 19444 36378 19472 37198
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19432 36372 19484 36378
rect 19432 36314 19484 36320
rect 19430 36136 19486 36145
rect 19430 36071 19486 36080
rect 19444 35766 19472 36071
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19996 35834 20024 37198
rect 20444 37188 20496 37194
rect 20444 37130 20496 37136
rect 20456 36786 20484 37130
rect 20720 36848 20772 36854
rect 20718 36816 20720 36825
rect 20772 36816 20774 36825
rect 20444 36780 20496 36786
rect 20718 36751 20774 36760
rect 20444 36722 20496 36728
rect 20168 36712 20220 36718
rect 20168 36654 20220 36660
rect 19984 35828 20036 35834
rect 19984 35770 20036 35776
rect 19432 35760 19484 35766
rect 19432 35702 19484 35708
rect 19800 35760 19852 35766
rect 19800 35702 19852 35708
rect 20076 35760 20128 35766
rect 20076 35702 20128 35708
rect 19812 35290 19840 35702
rect 19984 35692 20036 35698
rect 19984 35634 20036 35640
rect 19800 35284 19852 35290
rect 19800 35226 19852 35232
rect 19432 35148 19484 35154
rect 19432 35090 19484 35096
rect 19248 34740 19300 34746
rect 19248 34682 19300 34688
rect 19444 34649 19472 35090
rect 19996 35018 20024 35634
rect 20088 35154 20116 35702
rect 20180 35698 20208 36654
rect 20456 36174 20484 36722
rect 20628 36712 20680 36718
rect 20628 36654 20680 36660
rect 20640 36174 20668 36654
rect 20720 36304 20772 36310
rect 20720 36246 20772 36252
rect 20444 36168 20496 36174
rect 20444 36110 20496 36116
rect 20628 36168 20680 36174
rect 20628 36110 20680 36116
rect 20168 35692 20220 35698
rect 20168 35634 20220 35640
rect 20260 35488 20312 35494
rect 20260 35430 20312 35436
rect 20076 35148 20128 35154
rect 20076 35090 20128 35096
rect 19984 35012 20036 35018
rect 19984 34954 20036 34960
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19430 34640 19486 34649
rect 19996 34610 20024 34954
rect 19430 34575 19486 34584
rect 19984 34604 20036 34610
rect 19984 34546 20036 34552
rect 19432 34468 19484 34474
rect 19432 34410 19484 34416
rect 19444 33658 19472 34410
rect 19522 34096 19578 34105
rect 19522 34031 19524 34040
rect 19576 34031 19578 34040
rect 19524 34002 19576 34008
rect 19996 33998 20024 34546
rect 20272 34377 20300 35430
rect 20258 34368 20314 34377
rect 20258 34303 20314 34312
rect 20536 34128 20588 34134
rect 20536 34070 20588 34076
rect 19984 33992 20036 33998
rect 19984 33934 20036 33940
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19248 33652 19300 33658
rect 19248 33594 19300 33600
rect 19432 33652 19484 33658
rect 19432 33594 19484 33600
rect 19260 33114 19288 33594
rect 19340 33516 19392 33522
rect 19340 33458 19392 33464
rect 19248 33108 19300 33114
rect 19248 33050 19300 33056
rect 19352 32910 19380 33458
rect 19340 32904 19392 32910
rect 19340 32846 19392 32852
rect 19352 31754 19380 32846
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19996 32434 20024 33934
rect 20548 33930 20576 34070
rect 20536 33924 20588 33930
rect 20536 33866 20588 33872
rect 20640 33522 20668 36110
rect 20732 36106 20760 36246
rect 20720 36100 20772 36106
rect 20720 36042 20772 36048
rect 21270 35728 21326 35737
rect 20812 35692 20864 35698
rect 21270 35663 21326 35672
rect 21454 35728 21510 35737
rect 21454 35663 21510 35672
rect 20812 35634 20864 35640
rect 20824 34406 20852 35634
rect 21284 35329 21312 35663
rect 21086 35320 21142 35329
rect 21086 35255 21142 35264
rect 21270 35320 21326 35329
rect 21270 35255 21326 35264
rect 21100 35086 21128 35255
rect 21364 35216 21416 35222
rect 21364 35158 21416 35164
rect 21088 35080 21140 35086
rect 21088 35022 21140 35028
rect 20996 35012 21048 35018
rect 20996 34954 21048 34960
rect 21008 34649 21036 34954
rect 21376 34746 21404 35158
rect 21468 35057 21496 35663
rect 21454 35048 21510 35057
rect 21454 34983 21510 34992
rect 21364 34740 21416 34746
rect 21364 34682 21416 34688
rect 20994 34640 21050 34649
rect 20994 34575 21050 34584
rect 20720 34400 20772 34406
rect 20720 34342 20772 34348
rect 20812 34400 20864 34406
rect 20812 34342 20864 34348
rect 20732 34134 20760 34342
rect 20720 34128 20772 34134
rect 20720 34070 20772 34076
rect 20824 33998 20852 34342
rect 20812 33992 20864 33998
rect 20812 33934 20864 33940
rect 20824 33590 20852 33934
rect 20904 33856 20956 33862
rect 20904 33798 20956 33804
rect 20812 33584 20864 33590
rect 20812 33526 20864 33532
rect 20628 33516 20680 33522
rect 20628 33458 20680 33464
rect 20640 32910 20668 33458
rect 20720 33448 20772 33454
rect 20720 33390 20772 33396
rect 20732 32978 20760 33390
rect 20916 33114 20944 33798
rect 20904 33108 20956 33114
rect 20904 33050 20956 33056
rect 20720 32972 20772 32978
rect 20720 32914 20772 32920
rect 20628 32904 20680 32910
rect 20628 32846 20680 32852
rect 20076 32836 20128 32842
rect 20076 32778 20128 32784
rect 19432 32428 19484 32434
rect 19432 32370 19484 32376
rect 19984 32428 20036 32434
rect 19984 32370 20036 32376
rect 19444 31822 19472 32370
rect 20088 31822 20116 32778
rect 20352 32768 20404 32774
rect 20352 32710 20404 32716
rect 20260 32428 20312 32434
rect 20260 32370 20312 32376
rect 20168 31952 20220 31958
rect 20168 31894 20220 31900
rect 19432 31816 19484 31822
rect 19432 31758 19484 31764
rect 20076 31816 20128 31822
rect 20076 31758 20128 31764
rect 19340 31748 19392 31754
rect 19340 31690 19392 31696
rect 19338 31512 19394 31521
rect 19156 31476 19208 31482
rect 19156 31418 19208 31424
rect 19248 31476 19300 31482
rect 19338 31447 19394 31456
rect 19248 31418 19300 31424
rect 19260 31249 19288 31418
rect 19352 31414 19380 31447
rect 19340 31408 19392 31414
rect 19340 31350 19392 31356
rect 19444 31346 19472 31758
rect 19984 31748 20036 31754
rect 19984 31690 20036 31696
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19996 31346 20024 31690
rect 19432 31340 19484 31346
rect 19432 31282 19484 31288
rect 19984 31340 20036 31346
rect 19984 31282 20036 31288
rect 19246 31240 19302 31249
rect 19246 31175 19302 31184
rect 19432 31136 19484 31142
rect 19432 31078 19484 31084
rect 18786 30424 18842 30433
rect 18786 30359 18842 30368
rect 18880 30252 18932 30258
rect 18880 30194 18932 30200
rect 18696 30048 18748 30054
rect 18696 29990 18748 29996
rect 18708 28490 18736 29990
rect 18892 29578 18920 30194
rect 19444 30190 19472 31078
rect 20180 30938 20208 31894
rect 20272 31414 20300 32370
rect 20364 31482 20392 32710
rect 20732 32366 20760 32914
rect 20916 32434 20944 33050
rect 20904 32428 20956 32434
rect 20904 32370 20956 32376
rect 20720 32360 20772 32366
rect 20720 32302 20772 32308
rect 20732 31822 20760 32302
rect 20810 32056 20866 32065
rect 20810 31991 20812 32000
rect 20864 31991 20866 32000
rect 20812 31962 20864 31968
rect 20720 31816 20772 31822
rect 20720 31758 20772 31764
rect 20904 31680 20956 31686
rect 20904 31622 20956 31628
rect 20916 31482 20944 31622
rect 20352 31476 20404 31482
rect 20352 31418 20404 31424
rect 20904 31476 20956 31482
rect 20904 31418 20956 31424
rect 20260 31408 20312 31414
rect 20260 31350 20312 31356
rect 20168 30932 20220 30938
rect 20168 30874 20220 30880
rect 20272 30734 20300 31350
rect 20364 30802 20392 31418
rect 20718 31376 20774 31385
rect 20718 31311 20774 31320
rect 20444 31272 20496 31278
rect 20444 31214 20496 31220
rect 20352 30796 20404 30802
rect 20352 30738 20404 30744
rect 20260 30728 20312 30734
rect 20260 30670 20312 30676
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19614 30288 19670 30297
rect 19614 30223 19616 30232
rect 19668 30223 19670 30232
rect 19616 30194 19668 30200
rect 19432 30184 19484 30190
rect 19432 30126 19484 30132
rect 20272 30054 20300 30670
rect 20352 30320 20404 30326
rect 20352 30262 20404 30268
rect 20364 30122 20392 30262
rect 20352 30116 20404 30122
rect 20352 30058 20404 30064
rect 18972 30048 19024 30054
rect 18972 29990 19024 29996
rect 20260 30048 20312 30054
rect 20260 29990 20312 29996
rect 18788 29572 18840 29578
rect 18788 29514 18840 29520
rect 18880 29572 18932 29578
rect 18880 29514 18932 29520
rect 18696 28484 18748 28490
rect 18696 28426 18748 28432
rect 18800 28370 18828 29514
rect 18892 29306 18920 29514
rect 18880 29300 18932 29306
rect 18880 29242 18932 29248
rect 18984 29238 19012 29990
rect 19352 29838 19564 29866
rect 19352 29646 19380 29838
rect 19536 29832 19564 29838
rect 19616 29844 19668 29850
rect 19536 29804 19616 29832
rect 19616 29786 19668 29792
rect 19432 29776 19484 29782
rect 19432 29718 19484 29724
rect 19444 29646 19472 29718
rect 19340 29640 19392 29646
rect 19340 29582 19392 29588
rect 19432 29640 19484 29646
rect 19432 29582 19484 29588
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 18972 29232 19024 29238
rect 18972 29174 19024 29180
rect 19432 29164 19484 29170
rect 19432 29106 19484 29112
rect 20260 29164 20312 29170
rect 20364 29152 20392 30058
rect 20312 29124 20392 29152
rect 20260 29106 20312 29112
rect 18972 29028 19024 29034
rect 18972 28970 19024 28976
rect 18984 28626 19012 28970
rect 18972 28620 19024 28626
rect 18972 28562 19024 28568
rect 19156 28552 19208 28558
rect 19156 28494 19208 28500
rect 18708 28342 18828 28370
rect 18604 28144 18656 28150
rect 18604 28086 18656 28092
rect 18708 28014 18736 28342
rect 18696 28008 18748 28014
rect 18696 27950 18748 27956
rect 18880 28008 18932 28014
rect 18880 27950 18932 27956
rect 18512 27940 18564 27946
rect 18512 27882 18564 27888
rect 18432 27798 18552 27826
rect 18236 27464 18288 27470
rect 18236 27406 18288 27412
rect 18248 27130 18276 27406
rect 18236 27124 18288 27130
rect 18236 27066 18288 27072
rect 18144 26444 18196 26450
rect 18144 26386 18196 26392
rect 18328 26444 18380 26450
rect 18328 26386 18380 26392
rect 18340 26042 18368 26386
rect 18420 26376 18472 26382
rect 18420 26318 18472 26324
rect 18432 26042 18460 26318
rect 18328 26036 18380 26042
rect 18328 25978 18380 25984
rect 18420 26036 18472 26042
rect 18420 25978 18472 25984
rect 18236 25832 18288 25838
rect 18236 25774 18288 25780
rect 18248 25362 18276 25774
rect 18236 25356 18288 25362
rect 18236 25298 18288 25304
rect 18328 25220 18380 25226
rect 18328 25162 18380 25168
rect 18144 24608 18196 24614
rect 18144 24550 18196 24556
rect 18052 24404 18104 24410
rect 18052 24346 18104 24352
rect 17868 24268 17920 24274
rect 17868 24210 17920 24216
rect 17776 23656 17828 23662
rect 17776 23598 17828 23604
rect 17684 23316 17736 23322
rect 17684 23258 17736 23264
rect 17132 22976 17184 22982
rect 17132 22918 17184 22924
rect 17144 22710 17172 22918
rect 17132 22704 17184 22710
rect 17132 22646 17184 22652
rect 17132 22568 17184 22574
rect 17132 22510 17184 22516
rect 16868 22066 16988 22094
rect 16028 21480 16080 21486
rect 16028 21422 16080 21428
rect 16672 21480 16724 21486
rect 16672 21422 16724 21428
rect 16684 21146 16712 21422
rect 16672 21140 16724 21146
rect 16672 21082 16724 21088
rect 16672 20868 16724 20874
rect 16672 20810 16724 20816
rect 16684 20058 16712 20810
rect 16672 20052 16724 20058
rect 16672 19994 16724 20000
rect 16580 19916 16632 19922
rect 16580 19858 16632 19864
rect 16028 19236 16080 19242
rect 16028 19178 16080 19184
rect 16040 8974 16068 19178
rect 16592 19174 16620 19858
rect 16580 19168 16632 19174
rect 16580 19110 16632 19116
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 16028 8968 16080 8974
rect 16028 8910 16080 8916
rect 15936 3188 15988 3194
rect 15936 3130 15988 3136
rect 16132 3058 16160 12038
rect 16868 10266 16896 22066
rect 17144 21894 17172 22510
rect 17788 21894 17816 23598
rect 17880 23118 17908 24210
rect 18064 24206 18092 24346
rect 18052 24200 18104 24206
rect 18052 24142 18104 24148
rect 17868 23112 17920 23118
rect 17868 23054 17920 23060
rect 17868 22568 17920 22574
rect 17868 22510 17920 22516
rect 17132 21888 17184 21894
rect 17132 21830 17184 21836
rect 17776 21888 17828 21894
rect 17776 21830 17828 21836
rect 16948 20936 17000 20942
rect 16948 20878 17000 20884
rect 16960 20602 16988 20878
rect 16948 20596 17000 20602
rect 16948 20538 17000 20544
rect 17788 19174 17816 21830
rect 17880 21486 17908 22510
rect 17868 21480 17920 21486
rect 17868 21422 17920 21428
rect 17880 20534 17908 21422
rect 18064 21146 18092 24142
rect 18156 23798 18184 24550
rect 18340 24410 18368 25162
rect 18524 24682 18552 27798
rect 18892 27674 18920 27950
rect 19168 27878 19196 28494
rect 19248 28484 19300 28490
rect 19248 28426 19300 28432
rect 19260 27878 19288 28426
rect 19340 28008 19392 28014
rect 19340 27950 19392 27956
rect 19156 27872 19208 27878
rect 19156 27814 19208 27820
rect 19248 27872 19300 27878
rect 19248 27814 19300 27820
rect 18880 27668 18932 27674
rect 18880 27610 18932 27616
rect 18604 26988 18656 26994
rect 18604 26930 18656 26936
rect 18616 26858 18644 26930
rect 18604 26852 18656 26858
rect 18604 26794 18656 26800
rect 18892 26586 18920 27610
rect 18696 26580 18748 26586
rect 18696 26522 18748 26528
rect 18880 26580 18932 26586
rect 18880 26522 18932 26528
rect 18708 26314 18736 26522
rect 18696 26308 18748 26314
rect 18696 26250 18748 26256
rect 18604 26240 18656 26246
rect 18604 26182 18656 26188
rect 18512 24676 18564 24682
rect 18512 24618 18564 24624
rect 18328 24404 18380 24410
rect 18328 24346 18380 24352
rect 18328 24132 18380 24138
rect 18328 24074 18380 24080
rect 18340 23866 18368 24074
rect 18328 23860 18380 23866
rect 18328 23802 18380 23808
rect 18144 23792 18196 23798
rect 18144 23734 18196 23740
rect 18340 22642 18368 23802
rect 18616 23254 18644 26182
rect 19260 25770 19288 27814
rect 19352 27062 19380 27950
rect 19340 27056 19392 27062
rect 19340 26998 19392 27004
rect 19340 26920 19392 26926
rect 19340 26862 19392 26868
rect 19248 25764 19300 25770
rect 19248 25706 19300 25712
rect 19352 24682 19380 26862
rect 19444 25974 19472 29106
rect 19984 28416 20036 28422
rect 19984 28358 20036 28364
rect 20076 28416 20128 28422
rect 20076 28358 20128 28364
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19996 28082 20024 28358
rect 19984 28076 20036 28082
rect 19984 28018 20036 28024
rect 20088 27538 20116 28358
rect 20456 27538 20484 31214
rect 20732 30938 20760 31311
rect 20720 30932 20772 30938
rect 20720 30874 20772 30880
rect 20732 30258 20760 30874
rect 20812 30660 20864 30666
rect 20812 30602 20864 30608
rect 20720 30252 20772 30258
rect 20720 30194 20772 30200
rect 20824 29850 20852 30602
rect 21560 29850 21588 37334
rect 21928 37126 21956 39200
rect 22836 37460 22888 37466
rect 22836 37402 22888 37408
rect 22744 37256 22796 37262
rect 22744 37198 22796 37204
rect 21916 37120 21968 37126
rect 21916 37062 21968 37068
rect 22652 37120 22704 37126
rect 22652 37062 22704 37068
rect 22560 36848 22612 36854
rect 22560 36790 22612 36796
rect 22572 36582 22600 36790
rect 22560 36576 22612 36582
rect 22560 36518 22612 36524
rect 21640 36304 21692 36310
rect 21640 36246 21692 36252
rect 20812 29844 20864 29850
rect 20812 29786 20864 29792
rect 21548 29844 21600 29850
rect 21548 29786 21600 29792
rect 21560 29714 21588 29786
rect 21548 29708 21600 29714
rect 21548 29650 21600 29656
rect 20720 29640 20772 29646
rect 20720 29582 20772 29588
rect 20732 29102 20760 29582
rect 20904 29164 20956 29170
rect 20904 29106 20956 29112
rect 20720 29096 20772 29102
rect 20720 29038 20772 29044
rect 20076 27532 20128 27538
rect 20076 27474 20128 27480
rect 20444 27532 20496 27538
rect 20444 27474 20496 27480
rect 20352 27396 20404 27402
rect 20352 27338 20404 27344
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 20364 27130 20392 27338
rect 20352 27124 20404 27130
rect 20352 27066 20404 27072
rect 19524 27056 19576 27062
rect 19524 26998 19576 27004
rect 19536 26602 19564 26998
rect 19536 26586 19656 26602
rect 19536 26580 19668 26586
rect 19536 26574 19616 26580
rect 19616 26522 19668 26528
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19432 25968 19484 25974
rect 19432 25910 19484 25916
rect 19892 25832 19944 25838
rect 19892 25774 19944 25780
rect 19904 25226 19932 25774
rect 20456 25430 20484 27474
rect 20720 26988 20772 26994
rect 20720 26930 20772 26936
rect 20732 26586 20760 26930
rect 20536 26580 20588 26586
rect 20536 26522 20588 26528
rect 20720 26580 20772 26586
rect 20720 26522 20772 26528
rect 20548 26042 20576 26522
rect 20628 26376 20680 26382
rect 20628 26318 20680 26324
rect 20536 26036 20588 26042
rect 20536 25978 20588 25984
rect 20444 25424 20496 25430
rect 20444 25366 20496 25372
rect 19432 25220 19484 25226
rect 19432 25162 19484 25168
rect 19892 25220 19944 25226
rect 19892 25162 19944 25168
rect 19984 25220 20036 25226
rect 19984 25162 20036 25168
rect 18696 24676 18748 24682
rect 18696 24618 18748 24624
rect 19340 24676 19392 24682
rect 19340 24618 19392 24624
rect 18708 23798 18736 24618
rect 18696 23792 18748 23798
rect 18696 23734 18748 23740
rect 18604 23248 18656 23254
rect 18604 23190 18656 23196
rect 18328 22636 18380 22642
rect 18328 22578 18380 22584
rect 19352 22574 19380 24618
rect 19340 22568 19392 22574
rect 19340 22510 19392 22516
rect 18052 21140 18104 21146
rect 18052 21082 18104 21088
rect 18064 20942 18092 21082
rect 18052 20936 18104 20942
rect 18052 20878 18104 20884
rect 17868 20528 17920 20534
rect 17868 20470 17920 20476
rect 17776 19168 17828 19174
rect 17776 19110 17828 19116
rect 17788 18086 17816 19110
rect 17776 18080 17828 18086
rect 17776 18022 17828 18028
rect 17880 17338 17908 20470
rect 19444 18970 19472 25162
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19892 24744 19944 24750
rect 19892 24686 19944 24692
rect 19904 24290 19932 24686
rect 19996 24410 20024 25162
rect 20076 24948 20128 24954
rect 20076 24890 20128 24896
rect 20088 24410 20116 24890
rect 20640 24750 20668 26318
rect 20732 25974 20760 26522
rect 20720 25968 20772 25974
rect 20720 25910 20772 25916
rect 20628 24744 20680 24750
rect 20628 24686 20680 24692
rect 19984 24404 20036 24410
rect 19984 24346 20036 24352
rect 20076 24404 20128 24410
rect 20076 24346 20128 24352
rect 20732 24342 20760 25910
rect 20720 24336 20772 24342
rect 19904 24262 20024 24290
rect 20720 24278 20772 24284
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19432 18964 19484 18970
rect 19432 18906 19484 18912
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 17868 17332 17920 17338
rect 17868 17274 17920 17280
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19996 10810 20024 24262
rect 20916 22094 20944 29106
rect 21180 27328 21232 27334
rect 21180 27270 21232 27276
rect 21192 27062 21220 27270
rect 21180 27056 21232 27062
rect 21180 26998 21232 27004
rect 21652 26994 21680 36246
rect 22664 36106 22692 37062
rect 22756 36922 22784 37198
rect 22744 36916 22796 36922
rect 22744 36858 22796 36864
rect 22744 36712 22796 36718
rect 22744 36654 22796 36660
rect 22756 36242 22784 36654
rect 22848 36582 22876 37402
rect 22928 37120 22980 37126
rect 22928 37062 22980 37068
rect 22836 36576 22888 36582
rect 22836 36518 22888 36524
rect 22744 36236 22796 36242
rect 22744 36178 22796 36184
rect 22652 36100 22704 36106
rect 22652 36042 22704 36048
rect 22744 35692 22796 35698
rect 22744 35634 22796 35640
rect 22836 35692 22888 35698
rect 22836 35634 22888 35640
rect 22376 35556 22428 35562
rect 22376 35498 22428 35504
rect 22100 35488 22152 35494
rect 22098 35456 22100 35465
rect 22152 35456 22154 35465
rect 22098 35391 22154 35400
rect 22388 34950 22416 35498
rect 22756 35494 22784 35634
rect 22744 35488 22796 35494
rect 22744 35430 22796 35436
rect 22376 34944 22428 34950
rect 22376 34886 22428 34892
rect 21824 34672 21876 34678
rect 21824 34614 21876 34620
rect 21732 34196 21784 34202
rect 21732 34138 21784 34144
rect 21744 33114 21772 34138
rect 21732 33108 21784 33114
rect 21732 33050 21784 33056
rect 21836 32026 21864 34614
rect 22100 33856 22152 33862
rect 22100 33798 22152 33804
rect 22112 33318 22140 33798
rect 22100 33312 22152 33318
rect 22100 33254 22152 33260
rect 22112 32774 22140 33254
rect 22192 33040 22244 33046
rect 22192 32982 22244 32988
rect 22100 32768 22152 32774
rect 22100 32710 22152 32716
rect 22112 32366 22140 32710
rect 22204 32570 22232 32982
rect 22284 32904 22336 32910
rect 22284 32846 22336 32852
rect 22192 32564 22244 32570
rect 22192 32506 22244 32512
rect 22296 32450 22324 32846
rect 22204 32434 22324 32450
rect 22192 32428 22324 32434
rect 22244 32422 22324 32428
rect 22192 32370 22244 32376
rect 22100 32360 22152 32366
rect 22100 32302 22152 32308
rect 22112 32026 22140 32302
rect 21824 32020 21876 32026
rect 21824 31962 21876 31968
rect 22100 32020 22152 32026
rect 22100 31962 22152 31968
rect 22112 31482 22140 31962
rect 22204 31890 22232 32370
rect 22388 32314 22416 34886
rect 22756 34746 22784 35430
rect 22848 35222 22876 35634
rect 22836 35216 22888 35222
rect 22836 35158 22888 35164
rect 22744 34740 22796 34746
rect 22744 34682 22796 34688
rect 22836 34196 22888 34202
rect 22836 34138 22888 34144
rect 22744 33924 22796 33930
rect 22744 33866 22796 33872
rect 22296 32286 22416 32314
rect 22296 32230 22324 32286
rect 22284 32224 22336 32230
rect 22284 32166 22336 32172
rect 22192 31884 22244 31890
rect 22192 31826 22244 31832
rect 22100 31476 22152 31482
rect 22100 31418 22152 31424
rect 22204 30734 22232 31826
rect 22192 30728 22244 30734
rect 22192 30670 22244 30676
rect 21824 30592 21876 30598
rect 21824 30534 21876 30540
rect 21836 30394 21864 30534
rect 21824 30388 21876 30394
rect 21824 30330 21876 30336
rect 22296 27062 22324 32166
rect 22756 31754 22784 33866
rect 22848 33522 22876 34138
rect 22836 33516 22888 33522
rect 22836 33458 22888 33464
rect 22848 31958 22876 33458
rect 22836 31952 22888 31958
rect 22836 31894 22888 31900
rect 22664 31726 22784 31754
rect 22560 31476 22612 31482
rect 22560 31418 22612 31424
rect 22572 29850 22600 31418
rect 22560 29844 22612 29850
rect 22560 29786 22612 29792
rect 22664 28150 22692 31726
rect 22940 29306 22968 37062
rect 23860 36922 23888 39200
rect 23938 37360 23994 37369
rect 23938 37295 23940 37304
rect 23992 37295 23994 37304
rect 23940 37266 23992 37272
rect 25148 37126 25176 39200
rect 25320 37256 25372 37262
rect 25320 37198 25372 37204
rect 26516 37256 26568 37262
rect 26516 37198 26568 37204
rect 24768 37120 24820 37126
rect 24768 37062 24820 37068
rect 25136 37120 25188 37126
rect 25136 37062 25188 37068
rect 24780 36922 24808 37062
rect 23848 36916 23900 36922
rect 23848 36858 23900 36864
rect 24768 36916 24820 36922
rect 24768 36858 24820 36864
rect 23020 36780 23072 36786
rect 23020 36722 23072 36728
rect 23032 36378 23060 36722
rect 24032 36712 24084 36718
rect 24030 36680 24032 36689
rect 24084 36680 24086 36689
rect 24030 36615 24086 36624
rect 24676 36576 24728 36582
rect 23846 36544 23902 36553
rect 24676 36518 24728 36524
rect 23846 36479 23902 36488
rect 23860 36378 23888 36479
rect 23020 36372 23072 36378
rect 23020 36314 23072 36320
rect 23848 36372 23900 36378
rect 23848 36314 23900 36320
rect 24688 36038 24716 36518
rect 24676 36032 24728 36038
rect 24676 35974 24728 35980
rect 23204 35624 23256 35630
rect 23202 35592 23204 35601
rect 23256 35592 23258 35601
rect 23202 35527 23258 35536
rect 24688 35494 24716 35974
rect 23756 35488 23808 35494
rect 23756 35430 23808 35436
rect 24032 35488 24084 35494
rect 24032 35430 24084 35436
rect 24676 35488 24728 35494
rect 24676 35430 24728 35436
rect 23768 35329 23796 35430
rect 23754 35320 23810 35329
rect 23754 35255 23810 35264
rect 23204 35012 23256 35018
rect 23204 34954 23256 34960
rect 23216 34678 23244 34954
rect 24044 34950 24072 35430
rect 25134 35184 25190 35193
rect 25134 35119 25136 35128
rect 25188 35119 25190 35128
rect 25136 35090 25188 35096
rect 24032 34944 24084 34950
rect 24032 34886 24084 34892
rect 23204 34672 23256 34678
rect 23204 34614 23256 34620
rect 23216 34202 23244 34614
rect 24044 34474 24072 34886
rect 24308 34536 24360 34542
rect 24306 34504 24308 34513
rect 24360 34504 24362 34513
rect 24032 34468 24084 34474
rect 24306 34439 24362 34448
rect 24032 34410 24084 34416
rect 23664 34400 23716 34406
rect 23664 34342 23716 34348
rect 23204 34196 23256 34202
rect 23204 34138 23256 34144
rect 23216 33658 23244 34138
rect 23676 33862 23704 34342
rect 23664 33856 23716 33862
rect 23664 33798 23716 33804
rect 23204 33652 23256 33658
rect 23204 33594 23256 33600
rect 23216 33114 23244 33594
rect 23676 33114 23704 33798
rect 24044 33318 24072 34410
rect 25228 33992 25280 33998
rect 25228 33934 25280 33940
rect 25240 33658 25268 33934
rect 25228 33652 25280 33658
rect 25228 33594 25280 33600
rect 24032 33312 24084 33318
rect 24032 33254 24084 33260
rect 23204 33108 23256 33114
rect 23204 33050 23256 33056
rect 23664 33108 23716 33114
rect 23664 33050 23716 33056
rect 23676 31482 23704 33050
rect 24044 32774 24072 33254
rect 25240 33114 25268 33594
rect 25228 33108 25280 33114
rect 25228 33050 25280 33056
rect 24032 32768 24084 32774
rect 24032 32710 24084 32716
rect 24044 32366 24072 32710
rect 24032 32360 24084 32366
rect 24032 32302 24084 32308
rect 23664 31476 23716 31482
rect 23664 31418 23716 31424
rect 22928 29300 22980 29306
rect 22928 29242 22980 29248
rect 22836 28756 22888 28762
rect 22836 28698 22888 28704
rect 22652 28144 22704 28150
rect 22652 28086 22704 28092
rect 22664 27674 22692 28086
rect 22848 27674 22876 28698
rect 23572 28212 23624 28218
rect 23572 28154 23624 28160
rect 22652 27668 22704 27674
rect 22652 27610 22704 27616
rect 22836 27668 22888 27674
rect 22836 27610 22888 27616
rect 22664 27130 22692 27610
rect 22652 27124 22704 27130
rect 22652 27066 22704 27072
rect 22284 27056 22336 27062
rect 22284 26998 22336 27004
rect 21640 26988 21692 26994
rect 21640 26930 21692 26936
rect 22296 26790 22324 26998
rect 23584 26994 23612 28154
rect 25332 27130 25360 37198
rect 26528 37126 26556 37198
rect 27080 37126 27108 39200
rect 29012 37126 29040 39200
rect 30300 37346 30328 39200
rect 29184 37324 29236 37330
rect 30300 37318 30420 37346
rect 29184 37266 29236 37272
rect 26516 37120 26568 37126
rect 26516 37062 26568 37068
rect 27068 37120 27120 37126
rect 27068 37062 27120 37068
rect 28448 37120 28500 37126
rect 28448 37062 28500 37068
rect 29000 37120 29052 37126
rect 29000 37062 29052 37068
rect 25688 36712 25740 36718
rect 25688 36654 25740 36660
rect 25780 36712 25832 36718
rect 25780 36654 25832 36660
rect 25700 35290 25728 36654
rect 25688 35284 25740 35290
rect 25688 35226 25740 35232
rect 25792 35222 25820 36654
rect 26240 35488 26292 35494
rect 26240 35430 26292 35436
rect 26252 35290 26280 35430
rect 26240 35284 26292 35290
rect 26240 35226 26292 35232
rect 25780 35216 25832 35222
rect 25780 35158 25832 35164
rect 25688 34468 25740 34474
rect 25688 34410 25740 34416
rect 25700 34202 25728 34410
rect 25688 34196 25740 34202
rect 25688 34138 25740 34144
rect 26332 34196 26384 34202
rect 26332 34138 26384 34144
rect 25412 34128 25464 34134
rect 26344 34105 26372 34138
rect 25412 34070 25464 34076
rect 26330 34096 26386 34105
rect 25424 33998 25452 34070
rect 26330 34031 26386 34040
rect 25412 33992 25464 33998
rect 25412 33934 25464 33940
rect 26422 33552 26478 33561
rect 26422 33487 26424 33496
rect 26476 33487 26478 33496
rect 26424 33458 26476 33464
rect 25870 33416 25926 33425
rect 25870 33351 25872 33360
rect 25924 33351 25926 33360
rect 25872 33322 25924 33328
rect 25688 32904 25740 32910
rect 25686 32872 25688 32881
rect 25740 32872 25742 32881
rect 25686 32807 25742 32816
rect 26240 27940 26292 27946
rect 26240 27882 26292 27888
rect 25320 27124 25372 27130
rect 25320 27066 25372 27072
rect 23572 26988 23624 26994
rect 23572 26930 23624 26936
rect 22284 26784 22336 26790
rect 22284 26726 22336 26732
rect 20996 25900 21048 25906
rect 20996 25842 21048 25848
rect 21008 25702 21036 25842
rect 21088 25832 21140 25838
rect 21088 25774 21140 25780
rect 20996 25696 21048 25702
rect 20996 25638 21048 25644
rect 21008 25294 21036 25638
rect 21100 25498 21128 25774
rect 21088 25492 21140 25498
rect 21088 25434 21140 25440
rect 26252 25362 26280 27882
rect 26240 25356 26292 25362
rect 26240 25298 26292 25304
rect 20996 25288 21048 25294
rect 20996 25230 21048 25236
rect 20824 22066 20944 22094
rect 20824 20874 20852 22066
rect 26528 21078 26556 37062
rect 27068 36848 27120 36854
rect 27068 36790 27120 36796
rect 27080 36650 27108 36790
rect 27068 36644 27120 36650
rect 27068 36586 27120 36592
rect 28460 36582 28488 37062
rect 28448 36576 28500 36582
rect 28448 36518 28500 36524
rect 28460 36038 28488 36518
rect 27344 36032 27396 36038
rect 27344 35974 27396 35980
rect 27896 36032 27948 36038
rect 27896 35974 27948 35980
rect 28448 36032 28500 36038
rect 28448 35974 28500 35980
rect 29000 36032 29052 36038
rect 29000 35974 29052 35980
rect 27160 35760 27212 35766
rect 27158 35728 27160 35737
rect 27212 35728 27214 35737
rect 27158 35663 27214 35672
rect 27356 29714 27384 35974
rect 27908 31793 27936 35974
rect 28460 35562 28488 35974
rect 28448 35556 28500 35562
rect 28448 35498 28500 35504
rect 27988 35488 28040 35494
rect 27988 35430 28040 35436
rect 27894 31784 27950 31793
rect 27894 31719 27950 31728
rect 27344 29708 27396 29714
rect 27344 29650 27396 29656
rect 27252 23860 27304 23866
rect 27252 23802 27304 23808
rect 27264 23322 27292 23802
rect 28000 23322 28028 35430
rect 29012 34746 29040 35974
rect 29000 34740 29052 34746
rect 29000 34682 29052 34688
rect 29196 30190 29224 37266
rect 30392 37262 30420 37318
rect 29736 37256 29788 37262
rect 29642 37224 29698 37233
rect 29736 37198 29788 37204
rect 30380 37256 30432 37262
rect 30380 37198 30432 37204
rect 29642 37159 29698 37168
rect 29656 36718 29684 37159
rect 29748 36922 29776 37198
rect 30564 37188 30616 37194
rect 30564 37130 30616 37136
rect 29736 36916 29788 36922
rect 29736 36858 29788 36864
rect 29644 36712 29696 36718
rect 29644 36654 29696 36660
rect 30576 35698 30604 37130
rect 32232 37126 32260 39200
rect 32312 37256 32364 37262
rect 32312 37198 32364 37204
rect 32220 37120 32272 37126
rect 32220 37062 32272 37068
rect 32324 36786 32352 37198
rect 33520 37126 33548 39200
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 35452 37330 35480 39200
rect 37186 38856 37242 38865
rect 37186 38791 37242 38800
rect 35440 37324 35492 37330
rect 35440 37266 35492 37272
rect 33968 37256 34020 37262
rect 33968 37198 34020 37204
rect 33508 37120 33560 37126
rect 33508 37062 33560 37068
rect 32312 36780 32364 36786
rect 32312 36722 32364 36728
rect 30564 35692 30616 35698
rect 30564 35634 30616 35640
rect 29184 30184 29236 30190
rect 29184 30126 29236 30132
rect 29460 30048 29512 30054
rect 29460 29990 29512 29996
rect 29472 29782 29500 29990
rect 29460 29776 29512 29782
rect 29460 29718 29512 29724
rect 33980 28762 34008 37198
rect 36820 37120 36872 37126
rect 36820 37062 36872 37068
rect 36832 36854 36860 37062
rect 36820 36848 36872 36854
rect 36820 36790 36872 36796
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 37200 36378 37228 38791
rect 37384 37126 37412 39200
rect 38290 37496 38346 37505
rect 38200 37460 38252 37466
rect 38672 37466 38700 39200
rect 38290 37431 38346 37440
rect 38660 37460 38712 37466
rect 38200 37402 38252 37408
rect 37372 37120 37424 37126
rect 37372 37062 37424 37068
rect 38212 36854 38240 37402
rect 38200 36848 38252 36854
rect 38200 36790 38252 36796
rect 38016 36644 38068 36650
rect 38016 36586 38068 36592
rect 37464 36576 37516 36582
rect 37464 36518 37516 36524
rect 37924 36576 37976 36582
rect 37924 36518 37976 36524
rect 37188 36372 37240 36378
rect 37188 36314 37240 36320
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 37476 34202 37504 36518
rect 37936 36174 37964 36518
rect 37832 36168 37884 36174
rect 37832 36110 37884 36116
rect 37924 36168 37976 36174
rect 37924 36110 37976 36116
rect 37740 34672 37792 34678
rect 37740 34614 37792 34620
rect 37464 34196 37516 34202
rect 37464 34138 37516 34144
rect 37372 33380 37424 33386
rect 37372 33322 37424 33328
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 37280 30864 37332 30870
rect 37280 30806 37332 30812
rect 37292 30258 37320 30806
rect 37280 30252 37332 30258
rect 37280 30194 37332 30200
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 37384 29238 37412 33322
rect 37648 30184 37700 30190
rect 37648 30126 37700 30132
rect 37660 29510 37688 30126
rect 37648 29504 37700 29510
rect 37648 29446 37700 29452
rect 37372 29232 37424 29238
rect 37372 29174 37424 29180
rect 34520 29164 34572 29170
rect 34520 29106 34572 29112
rect 33968 28756 34020 28762
rect 33968 28698 34020 28704
rect 34532 28694 34560 29106
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34520 28688 34572 28694
rect 34520 28630 34572 28636
rect 30748 28552 30800 28558
rect 30748 28494 30800 28500
rect 34152 28552 34204 28558
rect 34152 28494 34204 28500
rect 30760 28121 30788 28494
rect 30746 28112 30802 28121
rect 30746 28047 30802 28056
rect 34164 27402 34192 28494
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34152 27396 34204 27402
rect 34152 27338 34204 27344
rect 34796 27396 34848 27402
rect 34796 27338 34848 27344
rect 27252 23316 27304 23322
rect 27252 23258 27304 23264
rect 27988 23316 28040 23322
rect 27988 23258 28040 23264
rect 27264 23118 27292 23258
rect 33692 23180 33744 23186
rect 33692 23122 33744 23128
rect 27252 23112 27304 23118
rect 27252 23054 27304 23060
rect 26516 21072 26568 21078
rect 26516 21014 26568 21020
rect 20812 20868 20864 20874
rect 20812 20810 20864 20816
rect 28540 19508 28592 19514
rect 28540 19450 28592 19456
rect 22376 18624 22428 18630
rect 22376 18566 22428 18572
rect 19984 10804 20036 10810
rect 19984 10746 20036 10752
rect 22008 10532 22060 10538
rect 22008 10474 22060 10480
rect 16856 10260 16908 10266
rect 16856 10202 16908 10208
rect 16868 10062 16896 10202
rect 16856 10056 16908 10062
rect 16856 9998 16908 10004
rect 18604 9988 18656 9994
rect 18604 9930 18656 9936
rect 18144 9104 18196 9110
rect 18144 9046 18196 9052
rect 16856 8900 16908 8906
rect 16856 8842 16908 8848
rect 15752 3052 15804 3058
rect 15752 2994 15804 3000
rect 16120 3052 16172 3058
rect 16120 2994 16172 3000
rect 15764 2650 15792 2994
rect 15752 2644 15804 2650
rect 15752 2586 15804 2592
rect 15660 2576 15712 2582
rect 15660 2518 15712 2524
rect 15384 2508 15436 2514
rect 15384 2450 15436 2456
rect 16868 2446 16896 8842
rect 18156 2446 18184 9046
rect 18616 2446 18644 9930
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 20628 3120 20680 3126
rect 20812 3120 20864 3126
rect 20680 3068 20812 3074
rect 20628 3062 20864 3068
rect 20640 3046 20852 3062
rect 22020 2446 22048 10474
rect 22388 7410 22416 18566
rect 24400 16992 24452 16998
rect 24400 16934 24452 16940
rect 22376 7404 22428 7410
rect 22376 7346 22428 7352
rect 22560 7200 22612 7206
rect 22560 7142 22612 7148
rect 22572 2446 22600 7142
rect 24412 6322 24440 16934
rect 24400 6316 24452 6322
rect 24400 6258 24452 6264
rect 24952 6112 25004 6118
rect 24952 6054 25004 6060
rect 23388 2848 23440 2854
rect 23388 2790 23440 2796
rect 6828 2440 6880 2446
rect 6828 2382 6880 2388
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 10876 2440 10928 2446
rect 10876 2382 10928 2388
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 18144 2440 18196 2446
rect 18144 2382 18196 2388
rect 18604 2440 18656 2446
rect 18604 2382 18656 2388
rect 22008 2440 22060 2446
rect 22008 2382 22060 2388
rect 22560 2440 22612 2446
rect 22560 2382 22612 2388
rect 4528 2372 4580 2378
rect 4528 2314 4580 2320
rect 3240 2304 3292 2310
rect 3240 2246 3292 2252
rect 1674 1456 1730 1465
rect 1674 1391 1730 1400
rect 3252 800 3280 2246
rect 4540 800 4568 2314
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 6472 800 6500 2246
rect 8404 800 8432 2246
rect 9692 800 9720 2382
rect 23400 2378 23428 2790
rect 24964 2446 24992 6054
rect 28552 2650 28580 19450
rect 29000 10668 29052 10674
rect 29000 10610 29052 10616
rect 29012 3058 29040 10610
rect 29000 3052 29052 3058
rect 29000 2994 29052 3000
rect 30288 2984 30340 2990
rect 30288 2926 30340 2932
rect 29184 2848 29236 2854
rect 29184 2790 29236 2796
rect 28540 2644 28592 2650
rect 28540 2586 28592 2592
rect 29196 2446 29224 2790
rect 30300 2582 30328 2926
rect 33704 2650 33732 23122
rect 34704 3188 34756 3194
rect 34704 3130 34756 3136
rect 33692 2644 33744 2650
rect 33692 2586 33744 2592
rect 30288 2576 30340 2582
rect 30288 2518 30340 2524
rect 34716 2446 34744 3130
rect 34808 2582 34836 27338
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 37280 25220 37332 25226
rect 37280 25162 37332 25168
rect 36820 25152 36872 25158
rect 36820 25094 36872 25100
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 36832 21554 36860 25094
rect 37292 23730 37320 25162
rect 37280 23724 37332 23730
rect 37280 23666 37332 23672
rect 36820 21548 36872 21554
rect 36820 21490 36872 21496
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 37660 16114 37688 29446
rect 37752 27062 37780 34614
rect 37740 27056 37792 27062
rect 37740 26998 37792 27004
rect 37740 26308 37792 26314
rect 37740 26250 37792 26256
rect 37752 25294 37780 26250
rect 37844 26042 37872 36110
rect 38028 34134 38056 36586
rect 38304 36378 38332 37431
rect 38660 37402 38712 37408
rect 38292 36372 38344 36378
rect 38292 36314 38344 36320
rect 38200 35488 38252 35494
rect 38198 35456 38200 35465
rect 38252 35456 38254 35465
rect 38198 35391 38254 35400
rect 38016 34128 38068 34134
rect 38016 34070 38068 34076
rect 38200 33516 38252 33522
rect 38200 33458 38252 33464
rect 38212 33425 38240 33458
rect 38198 33416 38254 33425
rect 38198 33351 38254 33360
rect 38016 32428 38068 32434
rect 38016 32370 38068 32376
rect 38028 29850 38056 32370
rect 38200 32224 38252 32230
rect 38200 32166 38252 32172
rect 38212 32065 38240 32166
rect 38198 32056 38254 32065
rect 38198 31991 38254 32000
rect 38200 30048 38252 30054
rect 38198 30016 38200 30025
rect 38252 30016 38254 30025
rect 38198 29951 38254 29960
rect 38016 29844 38068 29850
rect 38016 29786 38068 29792
rect 38200 29028 38252 29034
rect 38200 28970 38252 28976
rect 38212 28665 38240 28970
rect 38198 28656 38254 28665
rect 38198 28591 38254 28600
rect 37924 27328 37976 27334
rect 37924 27270 37976 27276
rect 37832 26036 37884 26042
rect 37832 25978 37884 25984
rect 37740 25288 37792 25294
rect 37740 25230 37792 25236
rect 37936 21434 37964 27270
rect 38200 26988 38252 26994
rect 38200 26930 38252 26936
rect 38212 26625 38240 26930
rect 38292 26852 38344 26858
rect 38292 26794 38344 26800
rect 38198 26616 38254 26625
rect 38198 26551 38254 26560
rect 38108 25288 38160 25294
rect 38108 25230 38160 25236
rect 38016 25152 38068 25158
rect 38016 25094 38068 25100
rect 38028 24818 38056 25094
rect 38016 24812 38068 24818
rect 38016 24754 38068 24760
rect 37752 21406 37964 21434
rect 37648 16108 37700 16114
rect 37648 16050 37700 16056
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 37280 12708 37332 12714
rect 37280 12650 37332 12656
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 37292 7546 37320 12650
rect 37280 7540 37332 7546
rect 37280 7482 37332 7488
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 37372 3392 37424 3398
rect 37372 3334 37424 3340
rect 37280 3120 37332 3126
rect 37280 3062 37332 3068
rect 36728 2984 36780 2990
rect 36728 2926 36780 2932
rect 36360 2848 36412 2854
rect 36360 2790 36412 2796
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34796 2576 34848 2582
rect 34796 2518 34848 2524
rect 36372 2446 36400 2790
rect 24952 2440 25004 2446
rect 24952 2382 25004 2388
rect 29184 2440 29236 2446
rect 29184 2382 29236 2388
rect 34704 2440 34756 2446
rect 34704 2382 34756 2388
rect 36360 2440 36412 2446
rect 36360 2382 36412 2388
rect 36740 2378 36768 2926
rect 37292 2514 37320 3062
rect 37384 2922 37412 3334
rect 37752 3126 37780 21406
rect 38120 19922 38148 25230
rect 38200 24608 38252 24614
rect 38198 24576 38200 24585
rect 38252 24576 38254 24585
rect 38198 24511 38254 24520
rect 38200 23520 38252 23526
rect 38200 23462 38252 23468
rect 38212 23225 38240 23462
rect 38198 23216 38254 23225
rect 38198 23151 38254 23160
rect 38200 21344 38252 21350
rect 38200 21286 38252 21292
rect 38212 21185 38240 21286
rect 38198 21176 38254 21185
rect 38198 21111 38254 21120
rect 38304 19938 38332 26794
rect 38384 26240 38436 26246
rect 38384 26182 38436 26188
rect 38396 25906 38424 26182
rect 38384 25900 38436 25906
rect 38384 25842 38436 25848
rect 38108 19916 38160 19922
rect 38108 19858 38160 19864
rect 38212 19910 38332 19938
rect 38212 19802 38240 19910
rect 38292 19848 38344 19854
rect 37936 19774 38240 19802
rect 38290 19816 38292 19825
rect 38344 19816 38346 19825
rect 37832 11144 37884 11150
rect 37832 11086 37884 11092
rect 37844 6118 37872 11086
rect 37936 7478 37964 19774
rect 38290 19751 38346 19760
rect 38304 19514 38332 19751
rect 38292 19508 38344 19514
rect 38292 19450 38344 19456
rect 38016 18284 38068 18290
rect 38016 18226 38068 18232
rect 38028 14482 38056 18226
rect 38292 16040 38344 16046
rect 38292 15982 38344 15988
rect 38304 15745 38332 15982
rect 38290 15736 38346 15745
rect 38290 15671 38292 15680
rect 38344 15671 38346 15680
rect 38292 15642 38344 15648
rect 38016 14476 38068 14482
rect 38016 14418 38068 14424
rect 38028 12238 38056 14418
rect 38292 14408 38344 14414
rect 38290 14376 38292 14385
rect 38344 14376 38346 14385
rect 38290 14311 38346 14320
rect 38304 14074 38332 14311
rect 38292 14068 38344 14074
rect 38292 14010 38344 14016
rect 38200 12844 38252 12850
rect 38200 12786 38252 12792
rect 38212 12345 38240 12786
rect 38198 12336 38254 12345
rect 38198 12271 38254 12280
rect 38016 12232 38068 12238
rect 38016 12174 38068 12180
rect 38016 12096 38068 12102
rect 38016 12038 38068 12044
rect 38028 8974 38056 12038
rect 38200 11076 38252 11082
rect 38200 11018 38252 11024
rect 38212 10985 38240 11018
rect 38198 10976 38254 10985
rect 38198 10911 38254 10920
rect 38016 8968 38068 8974
rect 38016 8910 38068 8916
rect 38198 8936 38254 8945
rect 38198 8871 38254 8880
rect 38212 8838 38240 8871
rect 38200 8832 38252 8838
rect 38200 8774 38252 8780
rect 37924 7472 37976 7478
rect 37924 7414 37976 7420
rect 38200 7404 38252 7410
rect 38200 7346 38252 7352
rect 38212 6905 38240 7346
rect 38198 6896 38254 6905
rect 38198 6831 38254 6840
rect 37832 6112 37884 6118
rect 37832 6054 37884 6060
rect 38396 5914 38424 25842
rect 38384 5908 38436 5914
rect 38384 5850 38436 5856
rect 38200 5636 38252 5642
rect 38200 5578 38252 5584
rect 38212 5545 38240 5578
rect 38198 5536 38254 5545
rect 38198 5471 38254 5480
rect 38108 3936 38160 3942
rect 38108 3878 38160 3884
rect 37740 3120 37792 3126
rect 37740 3062 37792 3068
rect 37372 2916 37424 2922
rect 37372 2858 37424 2864
rect 37280 2508 37332 2514
rect 37280 2450 37332 2456
rect 38120 2446 38148 3878
rect 38198 3496 38254 3505
rect 38198 3431 38254 3440
rect 38212 3398 38240 3431
rect 38200 3392 38252 3398
rect 38200 3334 38252 3340
rect 38200 3052 38252 3058
rect 38200 2994 38252 3000
rect 37188 2440 37240 2446
rect 38108 2440 38160 2446
rect 37188 2382 37240 2388
rect 38028 2388 38108 2394
rect 38028 2382 38160 2388
rect 11612 2372 11664 2378
rect 11612 2314 11664 2320
rect 14832 2372 14884 2378
rect 14832 2314 14884 2320
rect 23388 2372 23440 2378
rect 23388 2314 23440 2320
rect 28356 2372 28408 2378
rect 28356 2314 28408 2320
rect 33508 2372 33560 2378
rect 33508 2314 33560 2320
rect 36728 2372 36780 2378
rect 36728 2314 36780 2320
rect 11624 800 11652 2314
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 12912 800 12940 2246
rect 14844 800 14872 2314
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 18052 2304 18104 2310
rect 18052 2246 18104 2252
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 21272 2304 21324 2310
rect 21272 2246 21324 2252
rect 23204 2304 23256 2310
rect 23204 2246 23256 2252
rect 25136 2304 25188 2310
rect 25136 2246 25188 2252
rect 26424 2304 26476 2310
rect 26424 2246 26476 2252
rect 16776 800 16804 2246
rect 18064 800 18092 2246
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19996 800 20024 2246
rect 21284 800 21312 2246
rect 23216 800 23244 2246
rect 25148 800 25176 2246
rect 26436 800 26464 2246
rect 28368 800 28396 2314
rect 29644 2304 29696 2310
rect 29644 2246 29696 2252
rect 31760 2304 31812 2310
rect 31760 2246 31812 2252
rect 29656 800 29684 2246
rect 31772 1714 31800 2246
rect 31588 1686 31800 1714
rect 31588 800 31616 1686
rect 33520 800 33548 2314
rect 34796 2304 34848 2310
rect 34796 2246 34848 2252
rect 34808 800 34836 2246
rect 36740 800 36768 2314
rect 18 200 74 800
rect 1306 200 1362 800
rect 3238 200 3294 800
rect 4526 200 4582 800
rect 6458 200 6514 800
rect 8390 200 8446 800
rect 9678 200 9734 800
rect 11610 200 11666 800
rect 12898 200 12954 800
rect 14830 200 14886 800
rect 16762 200 16818 800
rect 18050 200 18106 800
rect 19982 200 20038 800
rect 21270 200 21326 800
rect 23202 200 23258 800
rect 25134 200 25190 800
rect 26422 200 26478 800
rect 28354 200 28410 800
rect 29642 200 29698 800
rect 31574 200 31630 800
rect 33506 200 33562 800
rect 34794 200 34850 800
rect 36726 200 36782 800
rect 37200 105 37228 2382
rect 38028 2366 38148 2382
rect 38028 800 38056 2366
rect 38212 2145 38240 2994
rect 38198 2136 38254 2145
rect 38198 2071 38254 2080
rect 38014 200 38070 800
rect 37186 96 37242 105
rect 37186 31 37242 40
<< via2 >>
rect 1674 32272 1730 32328
rect 1674 31340 1730 31376
rect 1674 31320 1676 31340
rect 1676 31320 1728 31340
rect 1728 31320 1730 31340
rect 3054 38800 3110 38856
rect 1858 31204 1914 31240
rect 1858 31184 1860 31204
rect 1860 31184 1912 31204
rect 1912 31184 1914 31204
rect 1674 30116 1730 30152
rect 1674 30096 1676 30116
rect 1676 30096 1728 30116
rect 1728 30096 1730 30116
rect 1674 29960 1730 30016
rect 1766 29008 1822 29064
rect 1674 27940 1730 27976
rect 1674 27920 1676 27940
rect 1676 27920 1728 27940
rect 1728 27920 1730 27940
rect 1674 26560 1730 26616
rect 1674 24556 1676 24576
rect 1676 24556 1728 24576
rect 1728 24556 1730 24576
rect 1674 24520 1730 24556
rect 1950 24656 2006 24712
rect 2502 33224 2558 33280
rect 2594 31728 2650 31784
rect 1674 22500 1730 22536
rect 1674 22480 1676 22500
rect 1676 22480 1728 22500
rect 1728 22480 1730 22500
rect 1582 21140 1638 21176
rect 1582 21120 1584 21140
rect 1584 21120 1636 21140
rect 1636 21120 1638 21140
rect 1582 20596 1638 20632
rect 1582 20576 1584 20596
rect 1584 20576 1636 20596
rect 1636 20576 1638 20596
rect 1582 19080 1638 19136
rect 1674 17720 1730 17776
rect 1674 15680 1730 15736
rect 1582 13640 1638 13696
rect 1674 12280 1730 12336
rect 1674 10240 1730 10296
rect 1674 8900 1730 8936
rect 1674 8880 1676 8900
rect 1676 8880 1728 8900
rect 1728 8880 1730 8900
rect 1582 6840 1638 6896
rect 2778 36760 2834 36816
rect 2962 35944 3018 36000
rect 2870 33516 2926 33552
rect 2870 33496 2872 33516
rect 2872 33496 2924 33516
rect 2924 33496 2926 33516
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 3054 32272 3110 32328
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 3330 32952 3386 33008
rect 3698 32816 3754 32872
rect 3698 32544 3754 32600
rect 2870 27376 2926 27432
rect 3882 31864 3938 31920
rect 4618 34620 4620 34640
rect 4620 34620 4672 34640
rect 4672 34620 4674 34640
rect 4618 34584 4674 34620
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 3698 24928 3754 24984
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 5722 35808 5778 35864
rect 5262 35708 5264 35728
rect 5264 35708 5316 35728
rect 5316 35708 5318 35728
rect 5262 35672 5318 35708
rect 5170 33088 5226 33144
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4526 28076 4582 28112
rect 4526 28056 4528 28076
rect 4528 28056 4580 28076
rect 4580 28056 4582 28076
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4066 26288 4122 26344
rect 4526 25880 4582 25936
rect 5078 28484 5134 28520
rect 5078 28464 5080 28484
rect 5080 28464 5132 28484
rect 5132 28464 5134 28484
rect 5078 28328 5134 28384
rect 4894 27004 4896 27024
rect 4896 27004 4948 27024
rect 4948 27004 4950 27024
rect 4894 26968 4950 27004
rect 4802 26152 4858 26208
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4618 25472 4674 25528
rect 5078 26424 5134 26480
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 3330 20052 3386 20088
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 3330 20032 3332 20052
rect 3332 20032 3384 20052
rect 3384 20032 3386 20052
rect 2226 18964 2282 19000
rect 2226 18944 2228 18964
rect 2228 18944 2280 18964
rect 2280 18944 2282 18964
rect 1582 4820 1638 4856
rect 1582 4800 1584 4820
rect 1584 4800 1636 4820
rect 1636 4800 1638 4820
rect 1674 3476 1676 3496
rect 1676 3476 1728 3496
rect 1728 3476 1730 3496
rect 1674 3440 1730 3476
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 5538 30912 5594 30968
rect 6366 32680 6422 32736
rect 6274 32000 6330 32056
rect 5446 28328 5502 28384
rect 5354 26424 5410 26480
rect 5446 26016 5502 26072
rect 5354 24556 5356 24576
rect 5356 24556 5408 24576
rect 5408 24556 5410 24576
rect 5354 24520 5410 24556
rect 5814 27376 5870 27432
rect 6182 27956 6184 27976
rect 6184 27956 6236 27976
rect 6236 27956 6238 27976
rect 6182 27920 6238 27956
rect 5814 25064 5870 25120
rect 5722 23316 5778 23352
rect 5722 23296 5724 23316
rect 5724 23296 5776 23316
rect 5776 23296 5778 23316
rect 7102 36488 7158 36544
rect 7654 35284 7710 35320
rect 7654 35264 7656 35284
rect 7656 35264 7708 35284
rect 7708 35264 7710 35284
rect 7378 35128 7434 35184
rect 6550 32408 6606 32464
rect 6734 31728 6790 31784
rect 6458 27104 6514 27160
rect 6642 26324 6644 26344
rect 6644 26324 6696 26344
rect 6696 26324 6698 26344
rect 6642 26288 6698 26324
rect 6826 28464 6882 28520
rect 7286 33108 7342 33144
rect 7286 33088 7288 33108
rect 7288 33088 7340 33108
rect 7340 33088 7342 33108
rect 7286 32544 7342 32600
rect 7286 31864 7342 31920
rect 7562 27512 7618 27568
rect 7562 27276 7564 27296
rect 7564 27276 7616 27296
rect 7616 27276 7618 27296
rect 7562 27240 7618 27276
rect 7378 26152 7434 26208
rect 7286 25880 7342 25936
rect 7378 25336 7434 25392
rect 7194 23588 7250 23624
rect 7194 23568 7196 23588
rect 7196 23568 7248 23588
rect 7248 23568 7250 23588
rect 8206 36116 8208 36136
rect 8208 36116 8260 36136
rect 8260 36116 8262 36136
rect 8206 36080 8262 36116
rect 9034 36216 9090 36272
rect 8298 35400 8354 35456
rect 8206 34740 8262 34776
rect 8206 34720 8208 34740
rect 8208 34720 8260 34740
rect 8260 34720 8262 34740
rect 8206 32000 8262 32056
rect 7838 27376 7894 27432
rect 7838 27004 7840 27024
rect 7840 27004 7892 27024
rect 7892 27004 7894 27024
rect 7838 26968 7894 27004
rect 8298 29280 8354 29336
rect 8298 27276 8300 27296
rect 8300 27276 8352 27296
rect 8352 27276 8354 27296
rect 8298 27240 8354 27276
rect 8114 26152 8170 26208
rect 7746 24148 7748 24168
rect 7748 24148 7800 24168
rect 7800 24148 7802 24168
rect 7746 24112 7802 24148
rect 7746 23724 7802 23760
rect 7746 23704 7748 23724
rect 7748 23704 7800 23724
rect 7800 23704 7802 23724
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 8942 35264 8998 35320
rect 8942 34584 8998 34640
rect 8942 34484 8944 34504
rect 8944 34484 8996 34504
rect 8996 34484 8998 34504
rect 8942 34448 8998 34484
rect 9126 35128 9182 35184
rect 10690 37440 10746 37496
rect 10966 37304 11022 37360
rect 10782 37168 10838 37224
rect 10598 35536 10654 35592
rect 10966 36796 10968 36816
rect 10968 36796 11020 36816
rect 11020 36796 11022 36816
rect 10966 36760 11022 36796
rect 10506 34604 10562 34640
rect 10506 34584 10508 34604
rect 10508 34584 10560 34604
rect 10560 34584 10562 34604
rect 8574 28056 8630 28112
rect 8482 24520 8538 24576
rect 10782 34176 10838 34232
rect 10598 34040 10654 34096
rect 10506 33224 10562 33280
rect 10598 32544 10654 32600
rect 9954 31728 10010 31784
rect 9586 29844 9642 29880
rect 9586 29824 9588 29844
rect 9588 29824 9640 29844
rect 9640 29824 9642 29844
rect 9678 29416 9734 29472
rect 9402 29280 9458 29336
rect 9586 28464 9642 28520
rect 9494 27648 9550 27704
rect 9310 27512 9366 27568
rect 9218 27104 9274 27160
rect 9126 25880 9182 25936
rect 10598 31728 10654 31784
rect 10782 32136 10838 32192
rect 9678 26308 9734 26344
rect 9678 26288 9680 26308
rect 9680 26288 9732 26308
rect 9732 26288 9734 26308
rect 8850 24656 8906 24712
rect 9770 25916 9772 25936
rect 9772 25916 9824 25936
rect 9824 25916 9826 25936
rect 9770 25880 9826 25916
rect 9218 23568 9274 23624
rect 10230 25100 10232 25120
rect 10232 25100 10284 25120
rect 10284 25100 10286 25120
rect 10230 25064 10286 25100
rect 10414 24112 10470 24168
rect 10414 23432 10470 23488
rect 10598 30640 10654 30696
rect 11150 34856 11206 34912
rect 11886 36916 11942 36952
rect 11886 36896 11888 36916
rect 11888 36896 11940 36916
rect 11940 36896 11942 36916
rect 11334 33904 11390 33960
rect 10782 29144 10838 29200
rect 11150 29280 11206 29336
rect 10874 26424 10930 26480
rect 10966 25900 11022 25936
rect 10966 25880 10968 25900
rect 10968 25880 11020 25900
rect 11020 25880 11022 25900
rect 11150 24656 11206 24712
rect 10966 23432 11022 23488
rect 11610 32680 11666 32736
rect 11518 32544 11574 32600
rect 12070 35400 12126 35456
rect 11886 34992 11942 35048
rect 11702 31864 11758 31920
rect 11702 31456 11758 31512
rect 11518 29572 11574 29608
rect 11518 29552 11520 29572
rect 11520 29552 11572 29572
rect 11572 29552 11574 29572
rect 12530 37168 12586 37224
rect 12898 36896 12954 36952
rect 12346 35264 12402 35320
rect 12346 34196 12402 34232
rect 12346 34176 12348 34196
rect 12348 34176 12400 34196
rect 12400 34176 12402 34196
rect 12438 34076 12440 34096
rect 12440 34076 12492 34096
rect 12492 34076 12494 34096
rect 12438 34040 12494 34076
rect 12438 33924 12494 33960
rect 12438 33904 12440 33924
rect 12440 33904 12492 33924
rect 12492 33904 12494 33924
rect 12070 33768 12126 33824
rect 13082 34584 13138 34640
rect 12806 34176 12862 34232
rect 13726 36372 13782 36408
rect 13726 36352 13728 36372
rect 13728 36352 13780 36372
rect 13780 36352 13782 36372
rect 14646 37188 14702 37224
rect 14646 37168 14648 37188
rect 14648 37168 14700 37188
rect 14700 37168 14702 37188
rect 15106 37032 15162 37088
rect 13818 35808 13874 35864
rect 13910 35264 13966 35320
rect 13726 34856 13782 34912
rect 13450 34312 13506 34368
rect 11978 32544 12034 32600
rect 12070 32308 12072 32328
rect 12072 32308 12124 32328
rect 12124 32308 12126 32328
rect 12070 32272 12126 32308
rect 12070 31864 12126 31920
rect 12070 30504 12126 30560
rect 12806 32136 12862 32192
rect 12530 31456 12586 31512
rect 12346 30776 12402 30832
rect 12714 30368 12770 30424
rect 12530 29844 12586 29880
rect 12530 29824 12532 29844
rect 12532 29824 12584 29844
rect 12584 29824 12586 29844
rect 13266 32680 13322 32736
rect 13358 31592 13414 31648
rect 12990 29688 13046 29744
rect 12622 25336 12678 25392
rect 13358 29688 13414 29744
rect 16026 37340 16028 37360
rect 16028 37340 16080 37360
rect 16080 37340 16082 37360
rect 16026 37304 16082 37340
rect 16302 37304 16358 37360
rect 15014 35944 15070 36000
rect 15750 35944 15806 36000
rect 15750 35808 15806 35864
rect 14922 35536 14978 35592
rect 15014 35264 15070 35320
rect 14186 34720 14242 34776
rect 14646 34720 14702 34776
rect 13910 33360 13966 33416
rect 13818 32272 13874 32328
rect 14830 34604 14886 34640
rect 14830 34584 14832 34604
rect 14832 34584 14884 34604
rect 14884 34584 14886 34604
rect 14186 32000 14242 32056
rect 13818 31592 13874 31648
rect 13910 30776 13966 30832
rect 13818 29960 13874 30016
rect 13634 29008 13690 29064
rect 14278 31864 14334 31920
rect 14094 29280 14150 29336
rect 14094 29044 14096 29064
rect 14096 29044 14148 29064
rect 14148 29044 14150 29064
rect 14094 29008 14150 29044
rect 14646 34040 14702 34096
rect 15198 34856 15254 34912
rect 15106 32136 15162 32192
rect 15382 33224 15438 33280
rect 15290 31456 15346 31512
rect 15198 30776 15254 30832
rect 14554 27648 14610 27704
rect 15198 29416 15254 29472
rect 15566 34992 15622 35048
rect 16578 37168 16634 37224
rect 18050 37440 18106 37496
rect 16762 36216 16818 36272
rect 15750 34992 15806 35048
rect 16210 34992 16266 35048
rect 15566 32136 15622 32192
rect 16026 32136 16082 32192
rect 15566 29708 15622 29744
rect 15566 29688 15568 29708
rect 15568 29688 15620 29708
rect 15620 29688 15622 29708
rect 15934 30504 15990 30560
rect 15842 29280 15898 29336
rect 16486 35400 16542 35456
rect 16946 35400 17002 35456
rect 16578 34584 16634 34640
rect 16946 32272 17002 32328
rect 16210 29180 16212 29200
rect 16212 29180 16264 29200
rect 16264 29180 16266 29200
rect 16210 29144 16266 29180
rect 11978 2624 12034 2680
rect 17038 31592 17094 31648
rect 17314 37032 17370 37088
rect 17314 36488 17370 36544
rect 17222 36216 17278 36272
rect 17314 35672 17370 35728
rect 17314 35400 17370 35456
rect 17222 34040 17278 34096
rect 17222 32408 17278 32464
rect 18602 36352 18658 36408
rect 17866 34856 17922 34912
rect 17866 34720 17922 34776
rect 17498 29552 17554 29608
rect 17314 27648 17370 27704
rect 17498 26424 17554 26480
rect 16118 23704 16174 23760
rect 17958 33768 18014 33824
rect 18326 34176 18382 34232
rect 18050 32680 18106 32736
rect 17958 32544 18014 32600
rect 17958 31884 18014 31920
rect 17958 31864 17960 31884
rect 17960 31864 18012 31884
rect 18012 31864 18014 31884
rect 17866 29960 17922 30016
rect 18326 32136 18382 32192
rect 18418 31184 18474 31240
rect 19062 36236 19118 36272
rect 19062 36216 19064 36236
rect 19064 36216 19116 36236
rect 19116 36216 19118 36236
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19430 36080 19486 36136
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 20718 36796 20720 36816
rect 20720 36796 20772 36816
rect 20772 36796 20774 36816
rect 20718 36760 20774 36796
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19430 34584 19486 34640
rect 19522 34060 19578 34096
rect 19522 34040 19524 34060
rect 19524 34040 19576 34060
rect 19576 34040 19578 34060
rect 20258 34312 20314 34368
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 21270 35672 21326 35728
rect 21454 35672 21510 35728
rect 21086 35264 21142 35320
rect 21270 35264 21326 35320
rect 21454 34992 21510 35048
rect 20994 34584 21050 34640
rect 19338 31456 19394 31512
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19246 31184 19302 31240
rect 18786 30368 18842 30424
rect 20810 32020 20866 32056
rect 20810 32000 20812 32020
rect 20812 32000 20864 32020
rect 20864 32000 20866 32020
rect 20718 31320 20774 31376
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19614 30252 19670 30288
rect 19614 30232 19616 30252
rect 19616 30232 19668 30252
rect 19668 30232 19670 30252
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 22098 35436 22100 35456
rect 22100 35436 22152 35456
rect 22152 35436 22154 35456
rect 22098 35400 22154 35436
rect 23938 37324 23994 37360
rect 23938 37304 23940 37324
rect 23940 37304 23992 37324
rect 23992 37304 23994 37324
rect 24030 36660 24032 36680
rect 24032 36660 24084 36680
rect 24084 36660 24086 36680
rect 24030 36624 24086 36660
rect 23846 36488 23902 36544
rect 23202 35572 23204 35592
rect 23204 35572 23256 35592
rect 23256 35572 23258 35592
rect 23202 35536 23258 35572
rect 23754 35264 23810 35320
rect 25134 35148 25190 35184
rect 25134 35128 25136 35148
rect 25136 35128 25188 35148
rect 25188 35128 25190 35148
rect 24306 34484 24308 34504
rect 24308 34484 24360 34504
rect 24360 34484 24362 34504
rect 24306 34448 24362 34484
rect 26330 34040 26386 34096
rect 26422 33516 26478 33552
rect 26422 33496 26424 33516
rect 26424 33496 26476 33516
rect 26476 33496 26478 33516
rect 25870 33380 25926 33416
rect 25870 33360 25872 33380
rect 25872 33360 25924 33380
rect 25924 33360 25926 33380
rect 25686 32852 25688 32872
rect 25688 32852 25740 32872
rect 25740 32852 25742 32872
rect 25686 32816 25742 32852
rect 27158 35708 27160 35728
rect 27160 35708 27212 35728
rect 27212 35708 27214 35728
rect 27158 35672 27214 35708
rect 27894 31728 27950 31784
rect 29642 37168 29698 37224
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 37186 38800 37242 38856
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 38290 37440 38346 37496
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 30746 28056 30802 28112
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 1674 1400 1730 1456
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 38198 35436 38200 35456
rect 38200 35436 38252 35456
rect 38252 35436 38254 35456
rect 38198 35400 38254 35436
rect 38198 33360 38254 33416
rect 38198 32000 38254 32056
rect 38198 29996 38200 30016
rect 38200 29996 38252 30016
rect 38252 29996 38254 30016
rect 38198 29960 38254 29996
rect 38198 28600 38254 28656
rect 38198 26560 38254 26616
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 38198 24556 38200 24576
rect 38200 24556 38252 24576
rect 38252 24556 38254 24576
rect 38198 24520 38254 24556
rect 38198 23160 38254 23216
rect 38198 21120 38254 21176
rect 38290 19796 38292 19816
rect 38292 19796 38344 19816
rect 38344 19796 38346 19816
rect 38290 19760 38346 19796
rect 38290 15700 38346 15736
rect 38290 15680 38292 15700
rect 38292 15680 38344 15700
rect 38344 15680 38346 15700
rect 38290 14356 38292 14376
rect 38292 14356 38344 14376
rect 38344 14356 38346 14376
rect 38290 14320 38346 14356
rect 38198 12280 38254 12336
rect 38198 10920 38254 10976
rect 38198 8880 38254 8936
rect 38198 6840 38254 6896
rect 38198 5480 38254 5536
rect 38198 3440 38254 3496
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 38198 2080 38254 2136
rect 37186 40 37242 96
<< metal3 >>
rect 200 38858 800 38888
rect 3049 38858 3115 38861
rect 200 38856 3115 38858
rect 200 38800 3054 38856
rect 3110 38800 3115 38856
rect 200 38798 3115 38800
rect 200 38768 800 38798
rect 3049 38795 3115 38798
rect 37181 38858 37247 38861
rect 39200 38858 39800 38888
rect 37181 38856 39800 38858
rect 37181 38800 37186 38856
rect 37242 38800 39800 38856
rect 37181 38798 39800 38800
rect 37181 38795 37247 38798
rect 39200 38768 39800 38798
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 10685 37498 10751 37501
rect 18045 37498 18111 37501
rect 10685 37496 18111 37498
rect 10685 37440 10690 37496
rect 10746 37440 18050 37496
rect 18106 37440 18111 37496
rect 10685 37438 18111 37440
rect 10685 37435 10751 37438
rect 18045 37435 18111 37438
rect 38285 37498 38351 37501
rect 39200 37498 39800 37528
rect 38285 37496 39800 37498
rect 38285 37440 38290 37496
rect 38346 37440 39800 37496
rect 38285 37438 39800 37440
rect 38285 37435 38351 37438
rect 39200 37408 39800 37438
rect 10961 37362 11027 37365
rect 16021 37362 16087 37365
rect 16297 37362 16363 37365
rect 23933 37362 23999 37365
rect 10961 37360 16087 37362
rect 10961 37304 10966 37360
rect 11022 37304 16026 37360
rect 16082 37304 16087 37360
rect 10961 37302 16087 37304
rect 10961 37299 11027 37302
rect 16021 37299 16087 37302
rect 16254 37360 23999 37362
rect 16254 37304 16302 37360
rect 16358 37304 23938 37360
rect 23994 37304 23999 37360
rect 16254 37302 23999 37304
rect 16254 37299 16363 37302
rect 23933 37299 23999 37302
rect 10777 37226 10843 37229
rect 12525 37226 12591 37229
rect 10777 37224 12591 37226
rect 10777 37168 10782 37224
rect 10838 37168 12530 37224
rect 12586 37168 12591 37224
rect 10777 37166 12591 37168
rect 10777 37163 10843 37166
rect 12525 37163 12591 37166
rect 14641 37226 14707 37229
rect 16254 37226 16314 37299
rect 14641 37224 16314 37226
rect 14641 37168 14646 37224
rect 14702 37168 16314 37224
rect 14641 37166 16314 37168
rect 16573 37226 16639 37229
rect 19374 37226 19380 37228
rect 16573 37224 19380 37226
rect 16573 37168 16578 37224
rect 16634 37168 19380 37224
rect 16573 37166 19380 37168
rect 14641 37163 14707 37166
rect 16573 37163 16639 37166
rect 19374 37164 19380 37166
rect 19444 37226 19450 37228
rect 29637 37226 29703 37229
rect 19444 37224 29703 37226
rect 19444 37168 29642 37224
rect 29698 37168 29703 37224
rect 19444 37166 29703 37168
rect 19444 37164 19450 37166
rect 29637 37163 29703 37166
rect 15101 37090 15167 37093
rect 17309 37090 17375 37093
rect 15101 37088 17375 37090
rect 15101 37032 15106 37088
rect 15162 37032 17314 37088
rect 17370 37032 17375 37088
rect 15101 37030 17375 37032
rect 15101 37027 15167 37030
rect 17309 37027 17375 37030
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 11881 36954 11947 36957
rect 12893 36954 12959 36957
rect 11881 36952 12959 36954
rect 11881 36896 11886 36952
rect 11942 36896 12898 36952
rect 12954 36896 12959 36952
rect 11881 36894 12959 36896
rect 11881 36891 11947 36894
rect 12893 36891 12959 36894
rect 200 36818 800 36848
rect 2773 36818 2839 36821
rect 200 36816 2839 36818
rect 200 36760 2778 36816
rect 2834 36760 2839 36816
rect 200 36758 2839 36760
rect 200 36728 800 36758
rect 2773 36755 2839 36758
rect 10961 36818 11027 36821
rect 20713 36818 20779 36821
rect 10961 36816 20779 36818
rect 10961 36760 10966 36816
rect 11022 36760 20718 36816
rect 20774 36760 20779 36816
rect 10961 36758 20779 36760
rect 10961 36755 11027 36758
rect 20713 36755 20779 36758
rect 24025 36682 24091 36685
rect 17174 36680 24091 36682
rect 17174 36624 24030 36680
rect 24086 36624 24091 36680
rect 17174 36622 24091 36624
rect 7097 36546 7163 36549
rect 17174 36546 17234 36622
rect 24025 36619 24091 36622
rect 7097 36544 17234 36546
rect 7097 36488 7102 36544
rect 7158 36488 17234 36544
rect 7097 36486 17234 36488
rect 17309 36546 17375 36549
rect 23841 36546 23907 36549
rect 17309 36544 23907 36546
rect 17309 36488 17314 36544
rect 17370 36488 23846 36544
rect 23902 36488 23907 36544
rect 17309 36486 23907 36488
rect 7097 36483 7163 36486
rect 17309 36483 17375 36486
rect 23841 36483 23907 36486
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 13721 36410 13787 36413
rect 18597 36410 18663 36413
rect 13721 36408 18663 36410
rect 13721 36352 13726 36408
rect 13782 36352 18602 36408
rect 18658 36352 18663 36408
rect 13721 36350 18663 36352
rect 13721 36347 13787 36350
rect 18597 36347 18663 36350
rect 9029 36274 9095 36277
rect 16757 36274 16823 36277
rect 9029 36272 16823 36274
rect 9029 36216 9034 36272
rect 9090 36216 16762 36272
rect 16818 36216 16823 36272
rect 9029 36214 16823 36216
rect 9029 36211 9095 36214
rect 16757 36211 16823 36214
rect 17217 36274 17283 36277
rect 19057 36274 19123 36277
rect 17217 36272 19123 36274
rect 17217 36216 17222 36272
rect 17278 36216 19062 36272
rect 19118 36216 19123 36272
rect 17217 36214 19123 36216
rect 17217 36211 17283 36214
rect 19057 36211 19123 36214
rect 8201 36138 8267 36141
rect 19425 36138 19491 36141
rect 8201 36136 19491 36138
rect 8201 36080 8206 36136
rect 8262 36080 19430 36136
rect 19486 36080 19491 36136
rect 8201 36078 19491 36080
rect 8201 36075 8267 36078
rect 19425 36075 19491 36078
rect 2814 35940 2820 36004
rect 2884 36002 2890 36004
rect 2957 36002 3023 36005
rect 2884 36000 3023 36002
rect 2884 35944 2962 36000
rect 3018 35944 3023 36000
rect 2884 35942 3023 35944
rect 2884 35940 2890 35942
rect 2957 35939 3023 35942
rect 14590 35940 14596 36004
rect 14660 36002 14666 36004
rect 15009 36002 15075 36005
rect 14660 36000 15075 36002
rect 14660 35944 15014 36000
rect 15070 35944 15075 36000
rect 14660 35942 15075 35944
rect 14660 35940 14666 35942
rect 15009 35939 15075 35942
rect 15142 35940 15148 36004
rect 15212 36002 15218 36004
rect 15745 36002 15811 36005
rect 15212 36000 16498 36002
rect 15212 35944 15750 36000
rect 15806 35944 16498 36000
rect 15212 35942 16498 35944
rect 15212 35940 15218 35942
rect 15745 35939 15811 35942
rect 5717 35866 5783 35869
rect 13813 35866 13879 35869
rect 15745 35866 15811 35869
rect 5717 35864 15811 35866
rect 5717 35808 5722 35864
rect 5778 35808 13818 35864
rect 13874 35808 15750 35864
rect 15806 35808 15811 35864
rect 5717 35806 15811 35808
rect 16438 35866 16498 35942
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 16438 35806 19442 35866
rect 5717 35803 5783 35806
rect 13813 35803 13879 35806
rect 15745 35803 15811 35806
rect 5257 35730 5323 35733
rect 17309 35730 17375 35733
rect 5257 35728 17375 35730
rect 5257 35672 5262 35728
rect 5318 35672 17314 35728
rect 17370 35672 17375 35728
rect 5257 35670 17375 35672
rect 19382 35730 19442 35806
rect 21265 35730 21331 35733
rect 19382 35728 21331 35730
rect 19382 35672 21270 35728
rect 21326 35672 21331 35728
rect 19382 35670 21331 35672
rect 5257 35667 5323 35670
rect 17309 35667 17375 35670
rect 21265 35667 21331 35670
rect 21449 35730 21515 35733
rect 27153 35730 27219 35733
rect 21449 35728 27219 35730
rect 21449 35672 21454 35728
rect 21510 35672 27158 35728
rect 27214 35672 27219 35728
rect 21449 35670 27219 35672
rect 21449 35667 21515 35670
rect 27153 35667 27219 35670
rect 10593 35594 10659 35597
rect 10593 35592 12772 35594
rect 10593 35536 10598 35592
rect 10654 35536 12772 35592
rect 10593 35534 12772 35536
rect 10593 35531 10659 35534
rect 200 35368 800 35488
rect 8293 35458 8359 35461
rect 12065 35458 12131 35461
rect 8293 35456 12131 35458
rect 8293 35400 8298 35456
rect 8354 35400 12070 35456
rect 12126 35400 12131 35456
rect 8293 35398 12131 35400
rect 12712 35458 12772 35534
rect 14406 35532 14412 35596
rect 14476 35594 14482 35596
rect 14917 35594 14983 35597
rect 23197 35594 23263 35597
rect 14476 35592 23263 35594
rect 14476 35536 14922 35592
rect 14978 35536 23202 35592
rect 23258 35536 23263 35592
rect 14476 35534 23263 35536
rect 14476 35532 14482 35534
rect 14917 35531 14983 35534
rect 23197 35531 23263 35534
rect 16481 35458 16547 35461
rect 12712 35456 16547 35458
rect 12712 35400 16486 35456
rect 16542 35400 16547 35456
rect 12712 35398 16547 35400
rect 8293 35395 8359 35398
rect 12065 35395 12131 35398
rect 16481 35395 16547 35398
rect 16798 35396 16804 35460
rect 16868 35458 16874 35460
rect 16941 35458 17007 35461
rect 16868 35456 17007 35458
rect 16868 35400 16946 35456
rect 17002 35400 17007 35456
rect 16868 35398 17007 35400
rect 16868 35396 16874 35398
rect 16941 35395 17007 35398
rect 17309 35458 17375 35461
rect 22093 35458 22159 35461
rect 17309 35456 22159 35458
rect 17309 35400 17314 35456
rect 17370 35400 22098 35456
rect 22154 35400 22159 35456
rect 17309 35398 22159 35400
rect 17309 35395 17375 35398
rect 22093 35395 22159 35398
rect 38193 35458 38259 35461
rect 39200 35458 39800 35488
rect 38193 35456 39800 35458
rect 38193 35400 38198 35456
rect 38254 35400 39800 35456
rect 38193 35398 39800 35400
rect 38193 35395 38259 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 39200 35368 39800 35398
rect 34930 35327 35246 35328
rect 7649 35322 7715 35325
rect 8937 35322 9003 35325
rect 7649 35320 9003 35322
rect 7649 35264 7654 35320
rect 7710 35264 8942 35320
rect 8998 35264 9003 35320
rect 7649 35262 9003 35264
rect 7649 35259 7715 35262
rect 8937 35259 9003 35262
rect 12341 35322 12407 35325
rect 13905 35322 13971 35325
rect 12341 35320 13971 35322
rect 12341 35264 12346 35320
rect 12402 35264 13910 35320
rect 13966 35264 13971 35320
rect 12341 35262 13971 35264
rect 12341 35259 12407 35262
rect 13905 35259 13971 35262
rect 15009 35322 15075 35325
rect 21081 35322 21147 35325
rect 15009 35320 21147 35322
rect 15009 35264 15014 35320
rect 15070 35264 21086 35320
rect 21142 35264 21147 35320
rect 15009 35262 21147 35264
rect 15009 35259 15075 35262
rect 21081 35259 21147 35262
rect 21265 35322 21331 35325
rect 23749 35322 23815 35325
rect 21265 35320 23815 35322
rect 21265 35264 21270 35320
rect 21326 35264 23754 35320
rect 23810 35264 23815 35320
rect 21265 35262 23815 35264
rect 21265 35259 21331 35262
rect 23749 35259 23815 35262
rect 7373 35186 7439 35189
rect 9121 35186 9187 35189
rect 25129 35186 25195 35189
rect 7373 35184 25195 35186
rect 7373 35128 7378 35184
rect 7434 35128 9126 35184
rect 9182 35128 25134 35184
rect 25190 35128 25195 35184
rect 7373 35126 25195 35128
rect 7373 35123 7439 35126
rect 9121 35123 9187 35126
rect 25129 35123 25195 35126
rect 11881 35050 11947 35053
rect 15561 35050 15627 35053
rect 11881 35048 15627 35050
rect 11881 34992 11886 35048
rect 11942 34992 15566 35048
rect 15622 34992 15627 35048
rect 11881 34990 15627 34992
rect 11881 34987 11947 34990
rect 15561 34987 15627 34990
rect 15745 35050 15811 35053
rect 16205 35050 16271 35053
rect 21449 35050 21515 35053
rect 15745 35048 21515 35050
rect 15745 34992 15750 35048
rect 15806 34992 16210 35048
rect 16266 34992 21454 35048
rect 21510 34992 21515 35048
rect 15745 34990 21515 34992
rect 15745 34987 15811 34990
rect 16205 34987 16271 34990
rect 21449 34987 21515 34990
rect 11145 34914 11211 34917
rect 13721 34914 13787 34917
rect 11145 34912 13787 34914
rect 11145 34856 11150 34912
rect 11206 34856 13726 34912
rect 13782 34856 13787 34912
rect 11145 34854 13787 34856
rect 11145 34851 11211 34854
rect 13721 34851 13787 34854
rect 15193 34914 15259 34917
rect 17861 34914 17927 34917
rect 15193 34912 17927 34914
rect 15193 34856 15198 34912
rect 15254 34856 17866 34912
rect 17922 34856 17927 34912
rect 15193 34854 17927 34856
rect 15193 34851 15259 34854
rect 17861 34851 17927 34854
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 8201 34778 8267 34781
rect 14181 34778 14247 34781
rect 8201 34776 14247 34778
rect 8201 34720 8206 34776
rect 8262 34720 14186 34776
rect 14242 34720 14247 34776
rect 8201 34718 14247 34720
rect 8201 34715 8267 34718
rect 14181 34715 14247 34718
rect 14641 34778 14707 34781
rect 17861 34778 17927 34781
rect 14641 34776 17927 34778
rect 14641 34720 14646 34776
rect 14702 34720 17866 34776
rect 17922 34720 17927 34776
rect 14641 34718 17927 34720
rect 14641 34715 14707 34718
rect 17861 34715 17927 34718
rect 4613 34644 4679 34645
rect 4613 34640 4660 34644
rect 4724 34642 4730 34644
rect 8937 34642 9003 34645
rect 10501 34642 10567 34645
rect 4613 34584 4618 34640
rect 4613 34580 4660 34584
rect 4724 34582 4770 34642
rect 8937 34640 10567 34642
rect 8937 34584 8942 34640
rect 8998 34584 10506 34640
rect 10562 34584 10567 34640
rect 8937 34582 10567 34584
rect 4724 34580 4730 34582
rect 4613 34579 4679 34580
rect 8937 34579 9003 34582
rect 10501 34579 10567 34582
rect 13077 34642 13143 34645
rect 14825 34642 14891 34645
rect 16573 34642 16639 34645
rect 13077 34640 16639 34642
rect 13077 34584 13082 34640
rect 13138 34584 14830 34640
rect 14886 34584 16578 34640
rect 16634 34584 16639 34640
rect 13077 34582 16639 34584
rect 13077 34579 13143 34582
rect 14825 34579 14891 34582
rect 16573 34579 16639 34582
rect 19425 34642 19491 34645
rect 20989 34642 21055 34645
rect 19425 34640 21055 34642
rect 19425 34584 19430 34640
rect 19486 34584 20994 34640
rect 21050 34584 21055 34640
rect 19425 34582 21055 34584
rect 19425 34579 19491 34582
rect 20989 34579 21055 34582
rect 8937 34506 9003 34509
rect 24301 34506 24367 34509
rect 8937 34504 24367 34506
rect 8937 34448 8942 34504
rect 8998 34448 24306 34504
rect 24362 34448 24367 34504
rect 8937 34446 24367 34448
rect 8937 34443 9003 34446
rect 24301 34443 24367 34446
rect 13445 34370 13511 34373
rect 20253 34370 20319 34373
rect 13445 34368 20319 34370
rect 13445 34312 13450 34368
rect 13506 34312 20258 34368
rect 20314 34312 20319 34368
rect 13445 34310 20319 34312
rect 13445 34307 13511 34310
rect 20253 34307 20319 34310
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 10777 34234 10843 34237
rect 12341 34234 12407 34237
rect 10777 34232 12407 34234
rect 10777 34176 10782 34232
rect 10838 34176 12346 34232
rect 12402 34176 12407 34232
rect 10777 34174 12407 34176
rect 10777 34171 10843 34174
rect 12341 34171 12407 34174
rect 12801 34234 12867 34237
rect 18321 34234 18387 34237
rect 12801 34232 19350 34234
rect 12801 34176 12806 34232
rect 12862 34176 18326 34232
rect 18382 34176 19350 34232
rect 12801 34174 19350 34176
rect 12801 34171 12867 34174
rect 18321 34171 18387 34174
rect 10593 34098 10659 34101
rect 12433 34098 12499 34101
rect 10593 34096 12499 34098
rect 10593 34040 10598 34096
rect 10654 34040 12438 34096
rect 12494 34040 12499 34096
rect 10593 34038 12499 34040
rect 10593 34035 10659 34038
rect 12433 34035 12499 34038
rect 14641 34098 14707 34101
rect 17217 34098 17283 34101
rect 14641 34096 17283 34098
rect 14641 34040 14646 34096
rect 14702 34040 17222 34096
rect 17278 34040 17283 34096
rect 14641 34038 17283 34040
rect 19290 34098 19350 34174
rect 19517 34098 19583 34101
rect 26325 34098 26391 34101
rect 19290 34096 26391 34098
rect 19290 34040 19522 34096
rect 19578 34040 26330 34096
rect 26386 34040 26391 34096
rect 19290 34038 26391 34040
rect 14641 34035 14707 34038
rect 17217 34035 17283 34038
rect 19517 34035 19583 34038
rect 26325 34035 26391 34038
rect 11329 33962 11395 33965
rect 12433 33962 12499 33965
rect 11329 33960 12499 33962
rect 11329 33904 11334 33960
rect 11390 33904 12438 33960
rect 12494 33904 12499 33960
rect 11329 33902 12499 33904
rect 11329 33899 11395 33902
rect 12433 33899 12499 33902
rect 12065 33826 12131 33829
rect 17953 33826 18019 33829
rect 12065 33824 18019 33826
rect 12065 33768 12070 33824
rect 12126 33768 17958 33824
rect 18014 33768 18019 33824
rect 12065 33766 18019 33768
rect 12065 33763 12131 33766
rect 17953 33763 18019 33766
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 2865 33554 2931 33557
rect 26417 33554 26483 33557
rect 2730 33552 26483 33554
rect 2730 33496 2870 33552
rect 2926 33496 26422 33552
rect 26478 33496 26483 33552
rect 2730 33494 26483 33496
rect 200 33418 800 33448
rect 2730 33418 2790 33494
rect 2865 33491 2931 33494
rect 26417 33491 26483 33494
rect 200 33358 2790 33418
rect 13905 33418 13971 33421
rect 25865 33418 25931 33421
rect 13905 33416 25931 33418
rect 13905 33360 13910 33416
rect 13966 33360 25870 33416
rect 25926 33360 25931 33416
rect 13905 33358 25931 33360
rect 200 33328 800 33358
rect 13905 33355 13971 33358
rect 25865 33355 25931 33358
rect 38193 33418 38259 33421
rect 39200 33418 39800 33448
rect 38193 33416 39800 33418
rect 38193 33360 38198 33416
rect 38254 33360 39800 33416
rect 38193 33358 39800 33360
rect 38193 33355 38259 33358
rect 39200 33328 39800 33358
rect 2497 33284 2563 33285
rect 2446 33282 2452 33284
rect 2406 33222 2452 33282
rect 2516 33280 2563 33284
rect 2558 33224 2563 33280
rect 2446 33220 2452 33222
rect 2516 33220 2563 33224
rect 2497 33219 2563 33220
rect 10501 33282 10567 33285
rect 15377 33282 15443 33285
rect 10501 33280 15443 33282
rect 10501 33224 10506 33280
rect 10562 33224 15382 33280
rect 15438 33224 15443 33280
rect 10501 33222 15443 33224
rect 10501 33219 10567 33222
rect 15377 33219 15443 33222
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 5165 33146 5231 33149
rect 7281 33146 7347 33149
rect 5165 33144 7347 33146
rect 5165 33088 5170 33144
rect 5226 33088 7286 33144
rect 7342 33088 7347 33144
rect 5165 33086 7347 33088
rect 5165 33083 5231 33086
rect 7281 33083 7347 33086
rect 3325 33010 3391 33013
rect 3918 33010 3924 33012
rect 3325 33008 3924 33010
rect 3325 32952 3330 33008
rect 3386 32952 3924 33008
rect 3325 32950 3924 32952
rect 3325 32947 3391 32950
rect 3918 32948 3924 32950
rect 3988 32948 3994 33012
rect 3693 32874 3759 32877
rect 25681 32874 25747 32877
rect 3693 32872 25747 32874
rect 3693 32816 3698 32872
rect 3754 32816 25686 32872
rect 25742 32816 25747 32872
rect 3693 32814 25747 32816
rect 3693 32811 3759 32814
rect 25681 32811 25747 32814
rect 6361 32738 6427 32741
rect 11605 32738 11671 32741
rect 13261 32738 13327 32741
rect 18045 32738 18111 32741
rect 6361 32736 9690 32738
rect 6361 32680 6366 32736
rect 6422 32680 9690 32736
rect 6361 32678 9690 32680
rect 6361 32675 6427 32678
rect 3693 32602 3759 32605
rect 7281 32602 7347 32605
rect 3693 32600 7347 32602
rect 3693 32544 3698 32600
rect 3754 32544 7286 32600
rect 7342 32544 7347 32600
rect 3693 32542 7347 32544
rect 9630 32602 9690 32678
rect 11605 32736 13186 32738
rect 11605 32680 11610 32736
rect 11666 32680 13186 32736
rect 11605 32678 13186 32680
rect 11605 32675 11671 32678
rect 10174 32602 10180 32604
rect 9630 32542 10180 32602
rect 3693 32539 3759 32542
rect 7281 32539 7347 32542
rect 10174 32540 10180 32542
rect 10244 32602 10250 32604
rect 10593 32602 10659 32605
rect 10244 32600 10659 32602
rect 10244 32544 10598 32600
rect 10654 32544 10659 32600
rect 10244 32542 10659 32544
rect 10244 32540 10250 32542
rect 10593 32539 10659 32542
rect 11513 32602 11579 32605
rect 11973 32602 12039 32605
rect 11513 32600 12039 32602
rect 11513 32544 11518 32600
rect 11574 32544 11978 32600
rect 12034 32544 12039 32600
rect 11513 32542 12039 32544
rect 13126 32602 13186 32678
rect 13261 32736 18111 32738
rect 13261 32680 13266 32736
rect 13322 32680 18050 32736
rect 18106 32680 18111 32736
rect 13261 32678 18111 32680
rect 13261 32675 13327 32678
rect 18045 32675 18111 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 17953 32602 18019 32605
rect 13126 32600 18019 32602
rect 13126 32544 17958 32600
rect 18014 32544 18019 32600
rect 13126 32542 18019 32544
rect 11513 32539 11579 32542
rect 11973 32539 12039 32542
rect 17953 32539 18019 32542
rect 6545 32466 6611 32469
rect 12566 32466 12572 32468
rect 6545 32464 12572 32466
rect 6545 32408 6550 32464
rect 6606 32408 12572 32464
rect 6545 32406 12572 32408
rect 6545 32403 6611 32406
rect 12566 32404 12572 32406
rect 12636 32404 12642 32468
rect 17217 32466 17283 32469
rect 14920 32464 17283 32466
rect 14920 32408 17222 32464
rect 17278 32408 17283 32464
rect 14920 32406 17283 32408
rect 1669 32330 1735 32333
rect 2262 32330 2268 32332
rect 1669 32328 2268 32330
rect 1669 32272 1674 32328
rect 1730 32272 2268 32328
rect 1669 32270 2268 32272
rect 1669 32267 1735 32270
rect 2262 32268 2268 32270
rect 2332 32330 2338 32332
rect 3049 32330 3115 32333
rect 2332 32328 3115 32330
rect 2332 32272 3054 32328
rect 3110 32272 3115 32328
rect 2332 32270 3115 32272
rect 2332 32268 2338 32270
rect 3049 32267 3115 32270
rect 12065 32330 12131 32333
rect 13813 32330 13879 32333
rect 12065 32328 13879 32330
rect 12065 32272 12070 32328
rect 12126 32272 13818 32328
rect 13874 32272 13879 32328
rect 12065 32270 13879 32272
rect 12065 32267 12131 32270
rect 13813 32267 13879 32270
rect 10777 32194 10843 32197
rect 12801 32194 12867 32197
rect 14920 32194 14980 32406
rect 17217 32403 17283 32406
rect 16941 32332 17007 32333
rect 16941 32328 16988 32332
rect 17052 32330 17058 32332
rect 16941 32272 16946 32328
rect 16941 32268 16988 32272
rect 17052 32270 17098 32330
rect 17052 32268 17058 32270
rect 16941 32267 17007 32268
rect 10777 32192 12867 32194
rect 10777 32136 10782 32192
rect 10838 32136 12806 32192
rect 12862 32136 12867 32192
rect 10777 32134 12867 32136
rect 10777 32131 10843 32134
rect 12801 32131 12867 32134
rect 14046 32134 14980 32194
rect 15101 32194 15167 32197
rect 15561 32194 15627 32197
rect 15101 32192 15627 32194
rect 15101 32136 15106 32192
rect 15162 32136 15566 32192
rect 15622 32136 15627 32192
rect 15101 32134 15627 32136
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 6269 32058 6335 32061
rect 8201 32058 8267 32061
rect 14046 32058 14106 32134
rect 15101 32131 15167 32134
rect 15561 32131 15627 32134
rect 16021 32194 16087 32197
rect 18321 32194 18387 32197
rect 16021 32192 18387 32194
rect 16021 32136 16026 32192
rect 16082 32136 18326 32192
rect 18382 32136 18387 32192
rect 16021 32134 18387 32136
rect 16021 32131 16087 32134
rect 18321 32131 18387 32134
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 6269 32056 14106 32058
rect 6269 32000 6274 32056
rect 6330 32000 8206 32056
rect 8262 32000 14106 32056
rect 6269 31998 14106 32000
rect 14181 32058 14247 32061
rect 20805 32058 20871 32061
rect 14181 32056 20871 32058
rect 14181 32000 14186 32056
rect 14242 32000 20810 32056
rect 20866 32000 20871 32056
rect 14181 31998 20871 32000
rect 6269 31995 6335 31998
rect 8201 31995 8267 31998
rect 14181 31995 14247 31998
rect 20805 31995 20871 31998
rect 38193 32058 38259 32061
rect 39200 32058 39800 32088
rect 38193 32056 39800 32058
rect 38193 32000 38198 32056
rect 38254 32000 39800 32056
rect 38193 31998 39800 32000
rect 38193 31995 38259 31998
rect 39200 31968 39800 31998
rect 3877 31922 3943 31925
rect 7281 31922 7347 31925
rect 3877 31920 7347 31922
rect 3877 31864 3882 31920
rect 3938 31864 7286 31920
rect 7342 31864 7347 31920
rect 3877 31862 7347 31864
rect 3877 31859 3943 31862
rect 7281 31859 7347 31862
rect 11697 31922 11763 31925
rect 12065 31922 12131 31925
rect 11697 31920 12131 31922
rect 11697 31864 11702 31920
rect 11758 31864 12070 31920
rect 12126 31864 12131 31920
rect 11697 31862 12131 31864
rect 11697 31859 11763 31862
rect 12065 31859 12131 31862
rect 14273 31922 14339 31925
rect 17953 31922 18019 31925
rect 14273 31920 18019 31922
rect 14273 31864 14278 31920
rect 14334 31864 17958 31920
rect 18014 31864 18019 31920
rect 14273 31862 18019 31864
rect 14273 31859 14339 31862
rect 17953 31859 18019 31862
rect 2589 31788 2655 31789
rect 2589 31784 2636 31788
rect 2700 31786 2706 31788
rect 6729 31786 6795 31789
rect 9949 31786 10015 31789
rect 2589 31728 2594 31784
rect 2589 31724 2636 31728
rect 2700 31726 2746 31786
rect 6729 31784 10015 31786
rect 6729 31728 6734 31784
rect 6790 31728 9954 31784
rect 10010 31728 10015 31784
rect 6729 31726 10015 31728
rect 2700 31724 2706 31726
rect 2589 31723 2655 31724
rect 6729 31723 6795 31726
rect 9949 31723 10015 31726
rect 10593 31786 10659 31789
rect 27889 31786 27955 31789
rect 10593 31784 27955 31786
rect 10593 31728 10598 31784
rect 10654 31728 27894 31784
rect 27950 31728 27955 31784
rect 10593 31726 27955 31728
rect 10593 31723 10659 31726
rect 27889 31723 27955 31726
rect 13353 31650 13419 31653
rect 13670 31650 13676 31652
rect 13353 31648 13676 31650
rect 13353 31592 13358 31648
rect 13414 31592 13676 31648
rect 13353 31590 13676 31592
rect 13353 31587 13419 31590
rect 13670 31588 13676 31590
rect 13740 31588 13746 31652
rect 13813 31650 13879 31653
rect 17033 31650 17099 31653
rect 13813 31648 17099 31650
rect 13813 31592 13818 31648
rect 13874 31592 17038 31648
rect 17094 31592 17099 31648
rect 13813 31590 17099 31592
rect 13813 31587 13879 31590
rect 17033 31587 17099 31590
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 11697 31514 11763 31517
rect 12525 31514 12591 31517
rect 11697 31512 12591 31514
rect 11697 31456 11702 31512
rect 11758 31456 12530 31512
rect 12586 31456 12591 31512
rect 11697 31454 12591 31456
rect 11697 31451 11763 31454
rect 12525 31451 12591 31454
rect 15285 31514 15351 31517
rect 19333 31514 19399 31517
rect 15285 31512 19399 31514
rect 15285 31456 15290 31512
rect 15346 31456 19338 31512
rect 19394 31456 19399 31512
rect 15285 31454 19399 31456
rect 15285 31451 15351 31454
rect 19333 31451 19399 31454
rect 200 31378 800 31408
rect 1669 31378 1735 31381
rect 200 31376 1735 31378
rect 200 31320 1674 31376
rect 1730 31320 1735 31376
rect 200 31318 1735 31320
rect 200 31288 800 31318
rect 1669 31315 1735 31318
rect 19374 31316 19380 31380
rect 19444 31378 19450 31380
rect 20713 31378 20779 31381
rect 19444 31376 20779 31378
rect 19444 31320 20718 31376
rect 20774 31320 20779 31376
rect 19444 31318 20779 31320
rect 19444 31316 19450 31318
rect 20713 31315 20779 31318
rect 1853 31242 1919 31245
rect 18413 31242 18479 31245
rect 19241 31242 19307 31245
rect 1853 31240 19307 31242
rect 1853 31184 1858 31240
rect 1914 31184 18418 31240
rect 18474 31184 19246 31240
rect 19302 31184 19307 31240
rect 1853 31182 19307 31184
rect 1853 31179 1919 31182
rect 18413 31179 18479 31182
rect 19241 31179 19307 31182
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 5533 30970 5599 30973
rect 16798 30970 16804 30972
rect 5533 30968 16804 30970
rect 5533 30912 5538 30968
rect 5594 30912 16804 30968
rect 5533 30910 16804 30912
rect 5533 30907 5599 30910
rect 16798 30908 16804 30910
rect 16868 30908 16874 30972
rect 12341 30834 12407 30837
rect 13905 30834 13971 30837
rect 15193 30834 15259 30837
rect 12341 30832 13971 30834
rect 12341 30776 12346 30832
rect 12402 30776 13910 30832
rect 13966 30776 13971 30832
rect 12341 30774 13971 30776
rect 12341 30771 12407 30774
rect 13905 30771 13971 30774
rect 15150 30832 15259 30834
rect 15150 30776 15198 30832
rect 15254 30776 15259 30832
rect 15150 30771 15259 30776
rect 10593 30698 10659 30701
rect 15150 30698 15210 30771
rect 10593 30696 15210 30698
rect 10593 30640 10598 30696
rect 10654 30640 15210 30696
rect 10593 30638 15210 30640
rect 10593 30635 10659 30638
rect 12065 30562 12131 30565
rect 15929 30562 15995 30565
rect 12065 30560 15995 30562
rect 12065 30504 12070 30560
rect 12126 30504 15934 30560
rect 15990 30504 15995 30560
rect 12065 30502 15995 30504
rect 12065 30499 12131 30502
rect 15929 30499 15995 30502
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 12709 30426 12775 30429
rect 18781 30426 18847 30429
rect 12709 30424 18847 30426
rect 12709 30368 12714 30424
rect 12770 30368 18786 30424
rect 18842 30368 18847 30424
rect 12709 30366 18847 30368
rect 12709 30363 12775 30366
rect 18781 30363 18847 30366
rect 12566 30228 12572 30292
rect 12636 30290 12642 30292
rect 19609 30290 19675 30293
rect 12636 30288 19675 30290
rect 12636 30232 19614 30288
rect 19670 30232 19675 30288
rect 12636 30230 19675 30232
rect 12636 30228 12642 30230
rect 19609 30227 19675 30230
rect 1669 30154 1735 30157
rect 15142 30154 15148 30156
rect 1669 30152 15148 30154
rect 1669 30096 1674 30152
rect 1730 30096 15148 30152
rect 1669 30094 15148 30096
rect 1669 30091 1735 30094
rect 15142 30092 15148 30094
rect 15212 30092 15218 30156
rect 200 30018 800 30048
rect 1669 30018 1735 30021
rect 200 30016 1735 30018
rect 200 29960 1674 30016
rect 1730 29960 1735 30016
rect 200 29958 1735 29960
rect 200 29928 800 29958
rect 1669 29955 1735 29958
rect 13813 30018 13879 30021
rect 17861 30018 17927 30021
rect 13813 30016 17927 30018
rect 13813 29960 13818 30016
rect 13874 29960 17866 30016
rect 17922 29960 17927 30016
rect 13813 29958 17927 29960
rect 13813 29955 13879 29958
rect 17861 29955 17927 29958
rect 38193 30018 38259 30021
rect 39200 30018 39800 30048
rect 38193 30016 39800 30018
rect 38193 29960 38198 30016
rect 38254 29960 39800 30016
rect 38193 29958 39800 29960
rect 38193 29955 38259 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 39200 29928 39800 29958
rect 34930 29887 35246 29888
rect 9581 29882 9647 29885
rect 12525 29882 12591 29885
rect 9581 29880 12591 29882
rect 9581 29824 9586 29880
rect 9642 29824 12530 29880
rect 12586 29824 12591 29880
rect 9581 29822 12591 29824
rect 9581 29819 9647 29822
rect 12525 29819 12591 29822
rect 12985 29746 13051 29749
rect 13353 29746 13419 29749
rect 12985 29744 13419 29746
rect 12985 29688 12990 29744
rect 13046 29688 13358 29744
rect 13414 29688 13419 29744
rect 12985 29686 13419 29688
rect 12985 29683 13051 29686
rect 13353 29683 13419 29686
rect 15561 29746 15627 29749
rect 16982 29746 16988 29748
rect 15561 29744 16988 29746
rect 15561 29688 15566 29744
rect 15622 29688 16988 29744
rect 15561 29686 16988 29688
rect 15561 29683 15627 29686
rect 16982 29684 16988 29686
rect 17052 29684 17058 29748
rect 11513 29610 11579 29613
rect 17493 29610 17559 29613
rect 11513 29608 17559 29610
rect 11513 29552 11518 29608
rect 11574 29552 17498 29608
rect 17554 29552 17559 29608
rect 11513 29550 17559 29552
rect 11513 29547 11579 29550
rect 17493 29547 17559 29550
rect 9673 29474 9739 29477
rect 15193 29474 15259 29477
rect 9673 29472 15259 29474
rect 9673 29416 9678 29472
rect 9734 29416 15198 29472
rect 15254 29416 15259 29472
rect 9673 29414 15259 29416
rect 9673 29411 9739 29414
rect 15193 29411 15259 29414
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 8293 29338 8359 29341
rect 9397 29338 9463 29341
rect 8293 29336 9463 29338
rect 8293 29280 8298 29336
rect 8354 29280 9402 29336
rect 9458 29280 9463 29336
rect 8293 29278 9463 29280
rect 8293 29275 8359 29278
rect 9397 29275 9463 29278
rect 11145 29338 11211 29341
rect 14089 29338 14155 29341
rect 15837 29338 15903 29341
rect 11145 29336 15903 29338
rect 11145 29280 11150 29336
rect 11206 29280 14094 29336
rect 14150 29280 15842 29336
rect 15898 29280 15903 29336
rect 11145 29278 15903 29280
rect 11145 29275 11211 29278
rect 14089 29275 14155 29278
rect 15837 29275 15903 29278
rect 10777 29202 10843 29205
rect 16205 29202 16271 29205
rect 10777 29200 16271 29202
rect 10777 29144 10782 29200
rect 10838 29144 16210 29200
rect 16266 29144 16271 29200
rect 10777 29142 16271 29144
rect 10777 29139 10843 29142
rect 16205 29139 16271 29142
rect 1761 29068 1827 29069
rect 1710 29066 1716 29068
rect 1670 29006 1716 29066
rect 1780 29064 1827 29068
rect 1822 29008 1827 29064
rect 1710 29004 1716 29006
rect 1780 29004 1827 29008
rect 1761 29003 1827 29004
rect 13629 29066 13695 29069
rect 14089 29066 14155 29069
rect 13629 29064 14155 29066
rect 13629 29008 13634 29064
rect 13690 29008 14094 29064
rect 14150 29008 14155 29064
rect 13629 29006 14155 29008
rect 13629 29003 13695 29006
rect 14089 29003 14155 29006
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 38193 28658 38259 28661
rect 39200 28658 39800 28688
rect 38193 28656 39800 28658
rect 38193 28600 38198 28656
rect 38254 28600 39800 28656
rect 38193 28598 39800 28600
rect 38193 28595 38259 28598
rect 39200 28568 39800 28598
rect 5073 28522 5139 28525
rect 6821 28522 6887 28525
rect 9581 28522 9647 28525
rect 5073 28520 9647 28522
rect 5073 28464 5078 28520
rect 5134 28464 6826 28520
rect 6882 28464 9586 28520
rect 9642 28464 9647 28520
rect 5073 28462 9647 28464
rect 5073 28459 5139 28462
rect 6821 28459 6887 28462
rect 9581 28459 9647 28462
rect 5073 28386 5139 28389
rect 5441 28386 5507 28389
rect 5073 28384 5507 28386
rect 5073 28328 5078 28384
rect 5134 28328 5446 28384
rect 5502 28328 5507 28384
rect 5073 28326 5507 28328
rect 5073 28323 5139 28326
rect 5441 28323 5507 28326
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 7598 28188 7604 28252
rect 7668 28250 7674 28252
rect 14590 28250 14596 28252
rect 7668 28190 14596 28250
rect 7668 28188 7674 28190
rect 14590 28188 14596 28190
rect 14660 28188 14666 28252
rect 4521 28114 4587 28117
rect 5390 28114 5396 28116
rect 4521 28112 5396 28114
rect 4521 28056 4526 28112
rect 4582 28056 5396 28112
rect 4521 28054 5396 28056
rect 4521 28051 4587 28054
rect 5390 28052 5396 28054
rect 5460 28114 5466 28116
rect 8569 28114 8635 28117
rect 30741 28114 30807 28117
rect 5460 28112 8635 28114
rect 5460 28056 8574 28112
rect 8630 28056 8635 28112
rect 5460 28054 8635 28056
rect 5460 28052 5466 28054
rect 8569 28051 8635 28054
rect 12390 28112 30807 28114
rect 12390 28056 30746 28112
rect 30802 28056 30807 28112
rect 12390 28054 30807 28056
rect 200 27978 800 28008
rect 1669 27978 1735 27981
rect 200 27976 1735 27978
rect 200 27920 1674 27976
rect 1730 27920 1735 27976
rect 200 27918 1735 27920
rect 200 27888 800 27918
rect 1669 27915 1735 27918
rect 5758 27916 5764 27980
rect 5828 27978 5834 27980
rect 6177 27978 6243 27981
rect 12390 27978 12450 28054
rect 30741 28051 30807 28054
rect 5828 27976 12450 27978
rect 5828 27920 6182 27976
rect 6238 27920 12450 27976
rect 5828 27918 12450 27920
rect 5828 27916 5834 27918
rect 6177 27915 6243 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 9489 27706 9555 27709
rect 10174 27706 10180 27708
rect 9489 27704 10180 27706
rect 9489 27648 9494 27704
rect 9550 27648 10180 27704
rect 9489 27646 10180 27648
rect 9489 27643 9555 27646
rect 10174 27644 10180 27646
rect 10244 27644 10250 27708
rect 14549 27706 14615 27709
rect 17309 27706 17375 27709
rect 14549 27704 17375 27706
rect 14549 27648 14554 27704
rect 14610 27648 17314 27704
rect 17370 27648 17375 27704
rect 14549 27646 17375 27648
rect 14549 27643 14615 27646
rect 17309 27643 17375 27646
rect 7557 27570 7623 27573
rect 9305 27570 9371 27573
rect 7557 27568 9371 27570
rect 7557 27512 7562 27568
rect 7618 27512 9310 27568
rect 9366 27512 9371 27568
rect 7557 27510 9371 27512
rect 7557 27507 7623 27510
rect 9305 27507 9371 27510
rect 2446 27372 2452 27436
rect 2516 27434 2522 27436
rect 2865 27434 2931 27437
rect 2516 27432 2931 27434
rect 2516 27376 2870 27432
rect 2926 27376 2931 27432
rect 2516 27374 2931 27376
rect 2516 27372 2522 27374
rect 2865 27371 2931 27374
rect 5809 27434 5875 27437
rect 7833 27434 7899 27437
rect 5809 27432 7899 27434
rect 5809 27376 5814 27432
rect 5870 27376 7838 27432
rect 7894 27376 7899 27432
rect 5809 27374 7899 27376
rect 5809 27371 5875 27374
rect 7833 27371 7899 27374
rect 7557 27298 7623 27301
rect 8293 27298 8359 27301
rect 7557 27296 8359 27298
rect 7557 27240 7562 27296
rect 7618 27240 8298 27296
rect 8354 27240 8359 27296
rect 7557 27238 8359 27240
rect 7557 27235 7623 27238
rect 8293 27235 8359 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 6453 27162 6519 27165
rect 9213 27162 9279 27165
rect 6453 27160 9279 27162
rect 6453 27104 6458 27160
rect 6514 27104 9218 27160
rect 9274 27104 9279 27160
rect 6453 27102 9279 27104
rect 6453 27099 6519 27102
rect 9213 27099 9279 27102
rect 4889 27026 4955 27029
rect 7833 27026 7899 27029
rect 4889 27024 7899 27026
rect 4889 26968 4894 27024
rect 4950 26968 7838 27024
rect 7894 26968 7899 27024
rect 4889 26966 7899 26968
rect 4889 26963 4955 26966
rect 7833 26963 7899 26966
rect 4210 26688 4526 26689
rect 200 26618 800 26648
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 1669 26618 1735 26621
rect 200 26616 1735 26618
rect 200 26560 1674 26616
rect 1730 26560 1735 26616
rect 200 26558 1735 26560
rect 200 26528 800 26558
rect 1669 26555 1735 26558
rect 38193 26618 38259 26621
rect 39200 26618 39800 26648
rect 38193 26616 39800 26618
rect 38193 26560 38198 26616
rect 38254 26560 39800 26616
rect 38193 26558 39800 26560
rect 38193 26555 38259 26558
rect 39200 26528 39800 26558
rect 5073 26482 5139 26485
rect 5349 26482 5415 26485
rect 5073 26480 5415 26482
rect 5073 26424 5078 26480
rect 5134 26424 5354 26480
rect 5410 26424 5415 26480
rect 5073 26422 5415 26424
rect 5073 26419 5139 26422
rect 5349 26419 5415 26422
rect 10869 26482 10935 26485
rect 17493 26482 17559 26485
rect 10869 26480 17559 26482
rect 10869 26424 10874 26480
rect 10930 26424 17498 26480
rect 17554 26424 17559 26480
rect 10869 26422 17559 26424
rect 10869 26419 10935 26422
rect 17493 26419 17559 26422
rect 4061 26346 4127 26349
rect 4654 26346 4660 26348
rect 4061 26344 4660 26346
rect 4061 26288 4066 26344
rect 4122 26288 4660 26344
rect 4061 26286 4660 26288
rect 4061 26283 4127 26286
rect 4654 26284 4660 26286
rect 4724 26284 4730 26348
rect 5390 26284 5396 26348
rect 5460 26284 5466 26348
rect 6637 26346 6703 26349
rect 9673 26346 9739 26349
rect 6637 26344 9739 26346
rect 6637 26288 6642 26344
rect 6698 26288 9678 26344
rect 9734 26288 9739 26344
rect 6637 26286 9739 26288
rect 3918 26148 3924 26212
rect 3988 26210 3994 26212
rect 4797 26210 4863 26213
rect 3988 26208 4863 26210
rect 3988 26152 4802 26208
rect 4858 26152 4863 26208
rect 3988 26150 4863 26152
rect 3988 26148 3994 26150
rect 4797 26147 4863 26150
rect 5398 26077 5458 26284
rect 6637 26283 6703 26286
rect 9673 26283 9739 26286
rect 7373 26210 7439 26213
rect 8109 26210 8175 26213
rect 7373 26208 8175 26210
rect 7373 26152 7378 26208
rect 7434 26152 8114 26208
rect 8170 26152 8175 26208
rect 7373 26150 8175 26152
rect 7373 26147 7439 26150
rect 8109 26147 8175 26150
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 5398 26072 5507 26077
rect 5398 26016 5446 26072
rect 5502 26016 5507 26072
rect 5398 26014 5507 26016
rect 5441 26011 5507 26014
rect 4521 25938 4587 25941
rect 7281 25938 7347 25941
rect 9121 25938 9187 25941
rect 4521 25936 9187 25938
rect 4521 25880 4526 25936
rect 4582 25880 7286 25936
rect 7342 25880 9126 25936
rect 9182 25880 9187 25936
rect 4521 25878 9187 25880
rect 4521 25875 4587 25878
rect 7281 25875 7347 25878
rect 9121 25875 9187 25878
rect 9765 25938 9831 25941
rect 10961 25938 11027 25941
rect 9765 25936 11027 25938
rect 9765 25880 9770 25936
rect 9826 25880 10966 25936
rect 11022 25880 11027 25936
rect 9765 25878 11027 25880
rect 9765 25875 9831 25878
rect 10961 25875 11027 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 4613 25530 4679 25533
rect 14406 25530 14412 25532
rect 4613 25528 14412 25530
rect 4613 25472 4618 25528
rect 4674 25472 14412 25528
rect 4613 25470 14412 25472
rect 4613 25467 4679 25470
rect 14406 25468 14412 25470
rect 14476 25468 14482 25532
rect 7373 25394 7439 25397
rect 12617 25394 12683 25397
rect 7373 25392 12683 25394
rect 7373 25336 7378 25392
rect 7434 25336 12622 25392
rect 12678 25336 12683 25392
rect 7373 25334 12683 25336
rect 7373 25331 7439 25334
rect 12617 25331 12683 25334
rect 5809 25122 5875 25125
rect 10225 25122 10291 25125
rect 5809 25120 10291 25122
rect 5809 25064 5814 25120
rect 5870 25064 10230 25120
rect 10286 25064 10291 25120
rect 5809 25062 10291 25064
rect 5809 25059 5875 25062
rect 10225 25059 10291 25062
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 2814 24924 2820 24988
rect 2884 24986 2890 24988
rect 3693 24986 3759 24989
rect 2884 24984 3759 24986
rect 2884 24928 3698 24984
rect 3754 24928 3759 24984
rect 2884 24926 3759 24928
rect 2884 24924 2890 24926
rect 3693 24923 3759 24926
rect 1945 24714 2011 24717
rect 7598 24714 7604 24716
rect 1945 24712 7604 24714
rect 1945 24656 1950 24712
rect 2006 24656 7604 24712
rect 1945 24654 7604 24656
rect 1945 24651 2011 24654
rect 7598 24652 7604 24654
rect 7668 24652 7674 24716
rect 8845 24714 8911 24717
rect 11145 24714 11211 24717
rect 8845 24712 11211 24714
rect 8845 24656 8850 24712
rect 8906 24656 11150 24712
rect 11206 24656 11211 24712
rect 8845 24654 11211 24656
rect 8845 24651 8911 24654
rect 11145 24651 11211 24654
rect 200 24578 800 24608
rect 1669 24578 1735 24581
rect 200 24576 1735 24578
rect 200 24520 1674 24576
rect 1730 24520 1735 24576
rect 200 24518 1735 24520
rect 200 24488 800 24518
rect 1669 24515 1735 24518
rect 5349 24578 5415 24581
rect 8477 24578 8543 24581
rect 5349 24576 8543 24578
rect 5349 24520 5354 24576
rect 5410 24520 8482 24576
rect 8538 24520 8543 24576
rect 5349 24518 8543 24520
rect 5349 24515 5415 24518
rect 8477 24515 8543 24518
rect 38193 24578 38259 24581
rect 39200 24578 39800 24608
rect 38193 24576 39800 24578
rect 38193 24520 38198 24576
rect 38254 24520 39800 24576
rect 38193 24518 39800 24520
rect 38193 24515 38259 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 39200 24488 39800 24518
rect 34930 24447 35246 24448
rect 7741 24170 7807 24173
rect 10409 24170 10475 24173
rect 7741 24168 10475 24170
rect 7741 24112 7746 24168
rect 7802 24112 10414 24168
rect 10470 24112 10475 24168
rect 7741 24110 10475 24112
rect 7741 24107 7807 24110
rect 10409 24107 10475 24110
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 7741 23762 7807 23765
rect 16113 23762 16179 23765
rect 7741 23760 16179 23762
rect 7741 23704 7746 23760
rect 7802 23704 16118 23760
rect 16174 23704 16179 23760
rect 7741 23702 16179 23704
rect 7741 23699 7807 23702
rect 16113 23699 16179 23702
rect 7189 23626 7255 23629
rect 9213 23626 9279 23629
rect 7189 23624 9279 23626
rect 7189 23568 7194 23624
rect 7250 23568 9218 23624
rect 9274 23568 9279 23624
rect 7189 23566 9279 23568
rect 7189 23563 7255 23566
rect 9213 23563 9279 23566
rect 10409 23490 10475 23493
rect 10961 23490 11027 23493
rect 10409 23488 11027 23490
rect 10409 23432 10414 23488
rect 10470 23432 10966 23488
rect 11022 23432 11027 23488
rect 10409 23430 11027 23432
rect 10409 23427 10475 23430
rect 10961 23427 11027 23430
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 5717 23356 5783 23357
rect 5717 23354 5764 23356
rect 5672 23352 5764 23354
rect 5672 23296 5722 23352
rect 5672 23294 5764 23296
rect 5717 23292 5764 23294
rect 5828 23292 5834 23356
rect 5717 23291 5783 23292
rect 38193 23218 38259 23221
rect 39200 23218 39800 23248
rect 38193 23216 39800 23218
rect 38193 23160 38198 23216
rect 38254 23160 39800 23216
rect 38193 23158 39800 23160
rect 38193 23155 38259 23158
rect 39200 23128 39800 23158
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 200 22538 800 22568
rect 1669 22538 1735 22541
rect 200 22536 1735 22538
rect 200 22480 1674 22536
rect 1730 22480 1735 22536
rect 200 22478 1735 22480
rect 200 22448 800 22478
rect 1669 22475 1735 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 200 21178 800 21208
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 1577 21178 1643 21181
rect 200 21176 1643 21178
rect 200 21120 1582 21176
rect 1638 21120 1643 21176
rect 200 21118 1643 21120
rect 200 21088 800 21118
rect 1577 21115 1643 21118
rect 38193 21178 38259 21181
rect 39200 21178 39800 21208
rect 38193 21176 39800 21178
rect 38193 21120 38198 21176
rect 38254 21120 39800 21176
rect 38193 21118 39800 21120
rect 38193 21115 38259 21118
rect 39200 21088 39800 21118
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 1577 20634 1643 20637
rect 1710 20634 1716 20636
rect 1577 20632 1716 20634
rect 1577 20576 1582 20632
rect 1638 20576 1716 20632
rect 1577 20574 1716 20576
rect 1577 20571 1643 20574
rect 1710 20572 1716 20574
rect 1780 20572 1786 20636
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 2630 20028 2636 20092
rect 2700 20090 2706 20092
rect 3325 20090 3391 20093
rect 2700 20088 3391 20090
rect 2700 20032 3330 20088
rect 3386 20032 3391 20088
rect 2700 20030 3391 20032
rect 2700 20028 2706 20030
rect 3325 20027 3391 20030
rect 38285 19818 38351 19821
rect 39200 19818 39800 19848
rect 38285 19816 39800 19818
rect 38285 19760 38290 19816
rect 38346 19760 39800 19816
rect 38285 19758 39800 19760
rect 38285 19755 38351 19758
rect 39200 19728 39800 19758
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 200 19138 800 19168
rect 1577 19138 1643 19141
rect 200 19136 1643 19138
rect 200 19080 1582 19136
rect 1638 19080 1643 19136
rect 200 19078 1643 19080
rect 200 19048 800 19078
rect 1577 19075 1643 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 2221 19004 2287 19005
rect 2221 19002 2268 19004
rect 2176 19000 2268 19002
rect 2176 18944 2226 19000
rect 2176 18942 2268 18944
rect 2221 18940 2268 18942
rect 2332 18940 2338 19004
rect 2221 18939 2287 18940
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 200 17778 800 17808
rect 1669 17778 1735 17781
rect 200 17776 1735 17778
rect 200 17720 1674 17776
rect 1730 17720 1735 17776
rect 200 17718 1735 17720
rect 200 17688 800 17718
rect 1669 17715 1735 17718
rect 39200 17688 39800 17808
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 200 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 1669 15738 1735 15741
rect 200 15736 1735 15738
rect 200 15680 1674 15736
rect 1730 15680 1735 15736
rect 200 15678 1735 15680
rect 200 15648 800 15678
rect 1669 15675 1735 15678
rect 38285 15738 38351 15741
rect 39200 15738 39800 15768
rect 38285 15736 39800 15738
rect 38285 15680 38290 15736
rect 38346 15680 39800 15736
rect 38285 15678 39800 15680
rect 38285 15675 38351 15678
rect 39200 15648 39800 15678
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 38285 14378 38351 14381
rect 39200 14378 39800 14408
rect 38285 14376 39800 14378
rect 38285 14320 38290 14376
rect 38346 14320 39800 14376
rect 38285 14318 39800 14320
rect 38285 14315 38351 14318
rect 39200 14288 39800 14318
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 200 13698 800 13728
rect 1577 13698 1643 13701
rect 200 13696 1643 13698
rect 200 13640 1582 13696
rect 1638 13640 1643 13696
rect 200 13638 1643 13640
rect 200 13608 800 13638
rect 1577 13635 1643 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 200 12338 800 12368
rect 1669 12338 1735 12341
rect 200 12336 1735 12338
rect 200 12280 1674 12336
rect 1730 12280 1735 12336
rect 200 12278 1735 12280
rect 200 12248 800 12278
rect 1669 12275 1735 12278
rect 38193 12338 38259 12341
rect 39200 12338 39800 12368
rect 38193 12336 39800 12338
rect 38193 12280 38198 12336
rect 38254 12280 39800 12336
rect 38193 12278 39800 12280
rect 38193 12275 38259 12278
rect 39200 12248 39800 12278
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 38193 10978 38259 10981
rect 39200 10978 39800 11008
rect 38193 10976 39800 10978
rect 38193 10920 38198 10976
rect 38254 10920 39800 10976
rect 38193 10918 39800 10920
rect 38193 10915 38259 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 39200 10888 39800 10918
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 200 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 1669 10298 1735 10301
rect 200 10296 1735 10298
rect 200 10240 1674 10296
rect 1730 10240 1735 10296
rect 200 10238 1735 10240
rect 200 10208 800 10238
rect 1669 10235 1735 10238
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 200 8938 800 8968
rect 1669 8938 1735 8941
rect 200 8936 1735 8938
rect 200 8880 1674 8936
rect 1730 8880 1735 8936
rect 200 8878 1735 8880
rect 200 8848 800 8878
rect 1669 8875 1735 8878
rect 38193 8938 38259 8941
rect 39200 8938 39800 8968
rect 38193 8936 39800 8938
rect 38193 8880 38198 8936
rect 38254 8880 39800 8936
rect 38193 8878 39800 8880
rect 38193 8875 38259 8878
rect 39200 8848 39800 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 200 6898 800 6928
rect 1577 6898 1643 6901
rect 200 6896 1643 6898
rect 200 6840 1582 6896
rect 1638 6840 1643 6896
rect 200 6838 1643 6840
rect 200 6808 800 6838
rect 1577 6835 1643 6838
rect 38193 6898 38259 6901
rect 39200 6898 39800 6928
rect 38193 6896 39800 6898
rect 38193 6840 38198 6896
rect 38254 6840 39800 6896
rect 38193 6838 39800 6840
rect 38193 6835 38259 6838
rect 39200 6808 39800 6838
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 38193 5538 38259 5541
rect 39200 5538 39800 5568
rect 38193 5536 39800 5538
rect 38193 5480 38198 5536
rect 38254 5480 39800 5536
rect 38193 5478 39800 5480
rect 38193 5475 38259 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 39200 5448 39800 5478
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 200 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 1577 4858 1643 4861
rect 200 4856 1643 4858
rect 200 4800 1582 4856
rect 1638 4800 1643 4856
rect 200 4798 1643 4800
rect 200 4768 800 4798
rect 1577 4795 1643 4798
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 200 3498 800 3528
rect 1669 3498 1735 3501
rect 200 3496 1735 3498
rect 200 3440 1674 3496
rect 1730 3440 1735 3496
rect 200 3438 1735 3440
rect 200 3408 800 3438
rect 1669 3435 1735 3438
rect 38193 3498 38259 3501
rect 39200 3498 39800 3528
rect 38193 3496 39800 3498
rect 38193 3440 38198 3496
rect 38254 3440 39800 3496
rect 38193 3438 39800 3440
rect 38193 3435 38259 3438
rect 39200 3408 39800 3438
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 11973 2682 12039 2685
rect 13670 2682 13676 2684
rect 11973 2680 13676 2682
rect 11973 2624 11978 2680
rect 12034 2624 13676 2680
rect 11973 2622 13676 2624
rect 11973 2619 12039 2622
rect 13670 2620 13676 2622
rect 13740 2620 13746 2684
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 38193 2138 38259 2141
rect 39200 2138 39800 2168
rect 38193 2136 39800 2138
rect 38193 2080 38198 2136
rect 38254 2080 39800 2136
rect 38193 2078 39800 2080
rect 38193 2075 38259 2078
rect 39200 2048 39800 2078
rect 200 1458 800 1488
rect 1669 1458 1735 1461
rect 200 1456 1735 1458
rect 200 1400 1674 1456
rect 1730 1400 1735 1456
rect 200 1398 1735 1400
rect 200 1368 800 1398
rect 1669 1395 1735 1398
rect 37181 98 37247 101
rect 39200 98 39800 128
rect 37181 96 39800 98
rect 37181 40 37186 96
rect 37242 40 39800 96
rect 37181 38 39800 40
rect 37181 35 37247 38
rect 39200 8 39800 38
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19380 37164 19444 37228
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 2820 35940 2884 36004
rect 14596 35940 14660 36004
rect 15148 35940 15212 36004
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 14412 35532 14476 35596
rect 16804 35396 16868 35460
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4660 34640 4724 34644
rect 4660 34584 4674 34640
rect 4674 34584 4724 34640
rect 4660 34580 4724 34584
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 2452 33280 2516 33284
rect 2452 33224 2502 33280
rect 2502 33224 2516 33280
rect 2452 33220 2516 33224
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 3924 32948 3988 33012
rect 10180 32540 10244 32604
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 12572 32404 12636 32468
rect 2268 32268 2332 32332
rect 16988 32328 17052 32332
rect 16988 32272 17002 32328
rect 17002 32272 17052 32328
rect 16988 32268 17052 32272
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 2636 31784 2700 31788
rect 2636 31728 2650 31784
rect 2650 31728 2700 31784
rect 2636 31724 2700 31728
rect 13676 31588 13740 31652
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 19380 31316 19444 31380
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 16804 30908 16868 30972
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 12572 30228 12636 30292
rect 15148 30092 15212 30156
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 16988 29684 17052 29748
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 1716 29064 1780 29068
rect 1716 29008 1766 29064
rect 1766 29008 1780 29064
rect 1716 29004 1780 29008
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 7604 28188 7668 28252
rect 14596 28188 14660 28252
rect 5396 28052 5460 28116
rect 5764 27916 5828 27980
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 10180 27644 10244 27708
rect 2452 27372 2516 27436
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 4660 26284 4724 26348
rect 5396 26284 5460 26348
rect 3924 26148 3988 26212
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 14412 25468 14476 25532
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 2820 24924 2884 24988
rect 7604 24652 7668 24716
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 5764 23352 5828 23356
rect 5764 23296 5778 23352
rect 5778 23296 5828 23352
rect 5764 23292 5828 23296
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 1716 20572 1780 20636
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 2636 20028 2700 20092
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 2268 19000 2332 19004
rect 2268 18944 2282 19000
rect 2282 18944 2332 19000
rect 2268 18940 2332 18944
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 13676 2620 13740 2684
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 19379 37228 19445 37229
rect 19379 37164 19380 37228
rect 19444 37164 19445 37228
rect 19379 37163 19445 37164
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 2819 36004 2885 36005
rect 2819 35940 2820 36004
rect 2884 35940 2885 36004
rect 2819 35939 2885 35940
rect 2451 33284 2517 33285
rect 2451 33220 2452 33284
rect 2516 33220 2517 33284
rect 2451 33219 2517 33220
rect 2267 32332 2333 32333
rect 2267 32268 2268 32332
rect 2332 32268 2333 32332
rect 2267 32267 2333 32268
rect 1715 29068 1781 29069
rect 1715 29004 1716 29068
rect 1780 29004 1781 29068
rect 1715 29003 1781 29004
rect 1718 20637 1778 29003
rect 1715 20636 1781 20637
rect 1715 20572 1716 20636
rect 1780 20572 1781 20636
rect 1715 20571 1781 20572
rect 2270 19005 2330 32267
rect 2454 27437 2514 33219
rect 2635 31788 2701 31789
rect 2635 31724 2636 31788
rect 2700 31724 2701 31788
rect 2635 31723 2701 31724
rect 2451 27436 2517 27437
rect 2451 27372 2452 27436
rect 2516 27372 2517 27436
rect 2451 27371 2517 27372
rect 2638 20093 2698 31723
rect 2822 24989 2882 35939
rect 4208 35392 4528 36416
rect 14595 36004 14661 36005
rect 14595 35940 14596 36004
rect 14660 35940 14661 36004
rect 14595 35939 14661 35940
rect 15147 36004 15213 36005
rect 15147 35940 15148 36004
rect 15212 35940 15213 36004
rect 15147 35939 15213 35940
rect 14411 35596 14477 35597
rect 14411 35532 14412 35596
rect 14476 35532 14477 35596
rect 14411 35531 14477 35532
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4659 34644 4725 34645
rect 4659 34580 4660 34644
rect 4724 34580 4725 34644
rect 4659 34579 4725 34580
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 3923 33012 3989 33013
rect 3923 32948 3924 33012
rect 3988 32948 3989 33012
rect 3923 32947 3989 32948
rect 3926 26213 3986 32947
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 3923 26212 3989 26213
rect 3923 26148 3924 26212
rect 3988 26148 3989 26212
rect 3923 26147 3989 26148
rect 4208 25600 4528 26624
rect 4662 26349 4722 34579
rect 10179 32604 10245 32605
rect 10179 32540 10180 32604
rect 10244 32540 10245 32604
rect 10179 32539 10245 32540
rect 7603 28252 7669 28253
rect 7603 28188 7604 28252
rect 7668 28188 7669 28252
rect 7603 28187 7669 28188
rect 5395 28116 5461 28117
rect 5395 28052 5396 28116
rect 5460 28052 5461 28116
rect 5395 28051 5461 28052
rect 5398 26349 5458 28051
rect 5763 27980 5829 27981
rect 5763 27916 5764 27980
rect 5828 27916 5829 27980
rect 5763 27915 5829 27916
rect 4659 26348 4725 26349
rect 4659 26284 4660 26348
rect 4724 26284 4725 26348
rect 4659 26283 4725 26284
rect 5395 26348 5461 26349
rect 5395 26284 5396 26348
rect 5460 26284 5461 26348
rect 5395 26283 5461 26284
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 2819 24988 2885 24989
rect 2819 24924 2820 24988
rect 2884 24924 2885 24988
rect 2819 24923 2885 24924
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 5766 23357 5826 27915
rect 7606 24717 7666 28187
rect 10182 27709 10242 32539
rect 12571 32468 12637 32469
rect 12571 32404 12572 32468
rect 12636 32404 12637 32468
rect 12571 32403 12637 32404
rect 12574 30293 12634 32403
rect 13675 31652 13741 31653
rect 13675 31588 13676 31652
rect 13740 31588 13741 31652
rect 13675 31587 13741 31588
rect 12571 30292 12637 30293
rect 12571 30228 12572 30292
rect 12636 30228 12637 30292
rect 12571 30227 12637 30228
rect 10179 27708 10245 27709
rect 10179 27644 10180 27708
rect 10244 27644 10245 27708
rect 10179 27643 10245 27644
rect 7603 24716 7669 24717
rect 7603 24652 7604 24716
rect 7668 24652 7669 24716
rect 7603 24651 7669 24652
rect 5763 23356 5829 23357
rect 5763 23292 5764 23356
rect 5828 23292 5829 23356
rect 5763 23291 5829 23292
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 2635 20092 2701 20093
rect 2635 20028 2636 20092
rect 2700 20028 2701 20092
rect 2635 20027 2701 20028
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 2267 19004 2333 19005
rect 2267 18940 2268 19004
rect 2332 18940 2333 19004
rect 2267 18939 2333 18940
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 13678 2685 13738 31587
rect 14414 25533 14474 35531
rect 14598 28253 14658 35939
rect 15150 30157 15210 35939
rect 16803 35460 16869 35461
rect 16803 35396 16804 35460
rect 16868 35396 16869 35460
rect 16803 35395 16869 35396
rect 16806 30973 16866 35395
rect 16987 32332 17053 32333
rect 16987 32268 16988 32332
rect 17052 32268 17053 32332
rect 16987 32267 17053 32268
rect 16803 30972 16869 30973
rect 16803 30908 16804 30972
rect 16868 30908 16869 30972
rect 16803 30907 16869 30908
rect 15147 30156 15213 30157
rect 15147 30092 15148 30156
rect 15212 30092 15213 30156
rect 15147 30091 15213 30092
rect 16990 29749 17050 32267
rect 19382 31381 19442 37163
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19379 31380 19445 31381
rect 19379 31316 19380 31380
rect 19444 31316 19445 31380
rect 19379 31315 19445 31316
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 16987 29748 17053 29749
rect 16987 29684 16988 29748
rect 17052 29684 17053 29748
rect 16987 29683 17053 29684
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 14595 28252 14661 28253
rect 14595 28188 14596 28252
rect 14660 28188 14661 28252
rect 14595 28187 14661 28188
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 14411 25532 14477 25533
rect 14411 25468 14412 25532
rect 14476 25468 14477 25532
rect 14411 25467 14477 25468
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 13675 2684 13741 2685
rect 13675 2620 13676 2684
rect 13740 2620 13741 2684
rect 13675 2619 13741 2620
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__224__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14996 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__A
timestamp 1667941163
transform 1 0 19412 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__A
timestamp 1667941163
transform 1 0 20884 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__232__A
timestamp 1667941163
transform 1 0 20792 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__A
timestamp 1667941163
transform 1 0 18032 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__A
timestamp 1667941163
transform -1 0 18492 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A
timestamp 1667941163
transform 1 0 17848 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__A
timestamp 1667941163
transform -1 0 12880 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__A
timestamp 1667941163
transform -1 0 17020 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__A
timestamp 1667941163
transform 1 0 16928 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__A
timestamp 1667941163
transform 1 0 21344 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__248__A
timestamp 1667941163
transform -1 0 18492 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__A
timestamp 1667941163
transform 1 0 8464 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__A
timestamp 1667941163
transform 1 0 21896 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__A
timestamp 1667941163
transform 1 0 21344 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__A
timestamp 1667941163
transform 1 0 21712 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__A
timestamp 1667941163
transform -1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__A
timestamp 1667941163
transform -1 0 6716 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__A
timestamp 1667941163
transform -1 0 1748 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__A
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__A
timestamp 1667941163
transform 1 0 22816 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__A
timestamp 1667941163
transform -1 0 3956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__A
timestamp 1667941163
transform -1 0 4692 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__A
timestamp 1667941163
transform 1 0 22540 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__A
timestamp 1667941163
transform 1 0 20608 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__A
timestamp 1667941163
transform -1 0 22724 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__287__A
timestamp 1667941163
transform 1 0 22264 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__288__A
timestamp 1667941163
transform 1 0 20884 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__A
timestamp 1667941163
transform -1 0 2392 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__A
timestamp 1667941163
transform -1 0 7360 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__A
timestamp 1667941163
transform -1 0 21436 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__293__A
timestamp 1667941163
transform 1 0 20700 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__294__A
timestamp 1667941163
transform -1 0 22172 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__A
timestamp 1667941163
transform 1 0 13616 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__296__A
timestamp 1667941163
transform 1 0 21988 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__298__A
timestamp 1667941163
transform -1 0 22080 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__299__A
timestamp 1667941163
transform 1 0 21620 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__300__A
timestamp 1667941163
transform -1 0 22172 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__303__A
timestamp 1667941163
transform -1 0 22172 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__304__A
timestamp 1667941163
transform 1 0 22264 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__307__A
timestamp 1667941163
transform -1 0 7912 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__308__A
timestamp 1667941163
transform 1 0 11960 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__311__A
timestamp 1667941163
transform 1 0 9384 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__312__A
timestamp 1667941163
transform 1 0 10580 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__315__A
timestamp 1667941163
transform -1 0 13432 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__316__A
timestamp 1667941163
transform -1 0 13708 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__330__A
timestamp 1667941163
transform 1 0 16192 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__331__A
timestamp 1667941163
transform 1 0 20700 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__332__A
timestamp 1667941163
transform 1 0 20700 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__333__A
timestamp 1667941163
transform -1 0 5244 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__A
timestamp 1667941163
transform -1 0 6716 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__337__A
timestamp 1667941163
transform 1 0 3956 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__A
timestamp 1667941163
transform 1 0 4968 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__A
timestamp 1667941163
transform -1 0 21896 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__A
timestamp 1667941163
transform 1 0 3128 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__344__A
timestamp 1667941163
transform -1 0 20884 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__346__A
timestamp 1667941163
transform 1 0 16468 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__347__A
timestamp 1667941163
transform 1 0 5612 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__A
timestamp 1667941163
transform 1 0 22816 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__A
timestamp 1667941163
transform 1 0 5336 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__350__A
timestamp 1667941163
transform -1 0 21528 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__352__A
timestamp 1667941163
transform -1 0 4140 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__353__A
timestamp 1667941163
transform 1 0 20148 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__354__A
timestamp 1667941163
transform 1 0 12972 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__A
timestamp 1667941163
transform 1 0 14260 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__356__A
timestamp 1667941163
transform 1 0 25208 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__357__A
timestamp 1667941163
transform 1 0 4692 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__359__A
timestamp 1667941163
transform 1 0 12328 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__360__A
timestamp 1667941163
transform 1 0 20332 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__361__A
timestamp 1667941163
transform -1 0 16284 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__363__A
timestamp 1667941163
transform -1 0 7360 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__364__A
timestamp 1667941163
transform 1 0 11132 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__366__A
timestamp 1667941163
transform -1 0 20240 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__367__A
timestamp 1667941163
transform -1 0 21896 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__368__A
timestamp 1667941163
transform 1 0 25944 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__369__A
timestamp 1667941163
transform 1 0 21068 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__A
timestamp 1667941163
transform 1 0 21344 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__371__A
timestamp 1667941163
transform 1 0 4784 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__374__A
timestamp 1667941163
transform 1 0 9752 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__376__A
timestamp 1667941163
transform 1 0 4784 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__377__A
timestamp 1667941163
transform -1 0 11592 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__378__A
timestamp 1667941163
transform -1 0 16928 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__380__A
timestamp 1667941163
transform 1 0 13892 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__381__A
timestamp 1667941163
transform 1 0 19688 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__382__A
timestamp 1667941163
transform -1 0 31188 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__383__A
timestamp 1667941163
transform -1 0 20240 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__A
timestamp 1667941163
transform -1 0 19780 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__388__A
timestamp 1667941163
transform -1 0 5428 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__389__A
timestamp 1667941163
transform -1 0 22724 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__390__A
timestamp 1667941163
transform 1 0 29992 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__393__A
timestamp 1667941163
transform 1 0 2484 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__394__A
timestamp 1667941163
transform 1 0 20792 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__395__A
timestamp 1667941163
transform 1 0 4600 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__396__A
timestamp 1667941163
transform -1 0 25484 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__397__A
timestamp 1667941163
transform 1 0 24564 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__398__A
timestamp 1667941163
transform 1 0 21068 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__399__A
timestamp 1667941163
transform 1 0 4508 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__400__A
timestamp 1667941163
transform 1 0 3128 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__401__A
timestamp 1667941163
transform -1 0 2760 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__402__A
timestamp 1667941163
transform 1 0 25116 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__404__A
timestamp 1667941163
transform 1 0 4232 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__405__A
timestamp 1667941163
transform 1 0 26404 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__406__A
timestamp 1667941163
transform -1 0 3404 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__407__A
timestamp 1667941163
transform -1 0 2484 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__408__A
timestamp 1667941163
transform 1 0 2116 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__409__A
timestamp 1667941163
transform 1 0 22540 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__410__A
timestamp 1667941163
transform 1 0 22816 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__411__A
timestamp 1667941163
transform 1 0 23092 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__412__A
timestamp 1667941163
transform 1 0 23092 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__413__A
timestamp 1667941163
transform -1 0 29164 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__415__A
timestamp 1667941163
transform -1 0 23828 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__416__A
timestamp 1667941163
transform 1 0 7544 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__417__A
timestamp 1667941163
transform 1 0 23092 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__418__A
timestamp 1667941163
transform -1 0 4784 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__419__A
timestamp 1667941163
transform 1 0 3312 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__420__A
timestamp 1667941163
transform -1 0 1748 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__421__A
timestamp 1667941163
transform 1 0 3404 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__A
timestamp 1667941163
transform 1 0 5612 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__423__A
timestamp 1667941163
transform 1 0 23368 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__424__A
timestamp 1667941163
transform -1 0 23828 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__426__A
timestamp 1667941163
transform 1 0 2576 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__427__A
timestamp 1667941163
transform 1 0 2944 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__428__A
timestamp 1667941163
transform -1 0 2300 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__429__A
timestamp 1667941163
transform 1 0 3956 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__430__A
timestamp 1667941163
transform 1 0 3956 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__431__A
timestamp 1667941163
transform 1 0 2760 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__432__A
timestamp 1667941163
transform 1 0 3956 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__433__A
timestamp 1667941163
transform 1 0 22632 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__434__A
timestamp 1667941163
transform 1 0 3220 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__435__A
timestamp 1667941163
transform -1 0 25484 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__464__CLK
timestamp 1667941163
transform 1 0 28520 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__464__D
timestamp 1667941163
transform -1 0 29808 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__465__CLK
timestamp 1667941163
transform 1 0 25116 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__465__D
timestamp 1667941163
transform -1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__466__CLK
timestamp 1667941163
transform 1 0 3956 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__466__D
timestamp 1667941163
transform -1 0 5060 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__467__CLK
timestamp 1667941163
transform 1 0 24564 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__468__CLK
timestamp 1667941163
transform 1 0 24196 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__468__D
timestamp 1667941163
transform -1 0 23828 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__469__CLK
timestamp 1667941163
transform 1 0 24748 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__469__D
timestamp 1667941163
transform -1 0 24380 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__470__CLK
timestamp 1667941163
transform 1 0 5152 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__471__CLK
timestamp 1667941163
transform 1 0 28796 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__472__CLK
timestamp 1667941163
transform 1 0 4048 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__473__CLK
timestamp 1667941163
transform 1 0 23368 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__474__CLK
timestamp 1667941163
transform 1 0 25852 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__475__CLK
timestamp 1667941163
transform 1 0 25668 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__476__CLK
timestamp 1667941163
transform 1 0 5060 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__477__CLK
timestamp 1667941163
transform 1 0 3956 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__478__CLK
timestamp 1667941163
transform 1 0 5888 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__478__D
timestamp 1667941163
transform 1 0 5704 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__479__CLK
timestamp 1667941163
transform 1 0 22540 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__480__CLK
timestamp 1667941163
transform 1 0 22448 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__480__D
timestamp 1667941163
transform 1 0 9752 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__481__CLK
timestamp 1667941163
transform 1 0 25944 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__482__CLK
timestamp 1667941163
transform 1 0 28428 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__483__CLK
timestamp 1667941163
transform 1 0 27876 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__483__D
timestamp 1667941163
transform -1 0 29164 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__484__CLK
timestamp 1667941163
transform 1 0 26772 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__484__D
timestamp 1667941163
transform -1 0 25300 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__485__CLK
timestamp 1667941163
transform 1 0 21252 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__486__CLK
timestamp 1667941163
transform 1 0 5888 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__486__D
timestamp 1667941163
transform -1 0 7176 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__487__CLK
timestamp 1667941163
transform 1 0 5060 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__488__CLK
timestamp 1667941163
transform 1 0 28244 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__489__CLK
timestamp 1667941163
transform 1 0 27324 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__490__CLK
timestamp 1667941163
transform 1 0 4324 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__490__D
timestamp 1667941163
transform -1 0 5520 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__491__CLK
timestamp 1667941163
transform 1 0 6440 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__491__D
timestamp 1667941163
transform 1 0 5888 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__492__CLK
timestamp 1667941163
transform 1 0 23736 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__492__D
timestamp 1667941163
transform -1 0 23368 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__493__CLK
timestamp 1667941163
transform 1 0 27968 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__493__D
timestamp 1667941163
transform -1 0 27508 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__494__CLK
timestamp 1667941163
transform 1 0 26220 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__494__D
timestamp 1667941163
transform -1 0 26036 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__495__CLK
timestamp 1667941163
transform 1 0 24564 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__495__D
timestamp 1667941163
transform -1 0 23920 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__495__RESET_B
timestamp 1667941163
transform -1 0 24012 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__496__CLK
timestamp 1667941163
transform 1 0 3496 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__497__CLK
timestamp 1667941163
transform 1 0 24288 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__498__CLK
timestamp 1667941163
transform 1 0 23920 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__498__D
timestamp 1667941163
transform -1 0 24932 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__499__CLK
timestamp 1667941163
transform 1 0 4508 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__500__CLK
timestamp 1667941163
transform 1 0 27140 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__501__CLK
timestamp 1667941163
transform 1 0 27692 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__501__D
timestamp 1667941163
transform -1 0 27324 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__502__CLK
timestamp 1667941163
transform 1 0 23368 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__502__D
timestamp 1667941163
transform -1 0 22724 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__502__RESET_B
timestamp 1667941163
transform -1 0 23368 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__503__CLK
timestamp 1667941163
transform 1 0 6532 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__504__CLK
timestamp 1667941163
transform 1 0 14260 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__505__CLK
timestamp 1667941163
transform 1 0 23092 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__506__CLK
timestamp 1667941163
transform 1 0 25668 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__507__CLK
timestamp 1667941163
transform 1 0 24564 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__507__D
timestamp 1667941163
transform -1 0 23552 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__508__CLK
timestamp 1667941163
transform 1 0 29072 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__508__D
timestamp 1667941163
transform -1 0 28060 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__509__CLK
timestamp 1667941163
transform 1 0 22264 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__510__CLK
timestamp 1667941163
transform 1 0 5888 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__511__CLK
timestamp 1667941163
transform 1 0 23920 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__512__CLK
timestamp 1667941163
transform 1 0 21988 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__513__CLK
timestamp 1667941163
transform 1 0 24288 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__514__CLK
timestamp 1667941163
transform 1 0 25392 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__514__D
timestamp 1667941163
transform -1 0 24748 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__515__CLK
timestamp 1667941163
transform 1 0 22264 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__515__D
timestamp 1667941163
transform -1 0 8648 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__516__CLK
timestamp 1667941163
transform 1 0 22540 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__517__CLK
timestamp 1667941163
transform 1 0 26220 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__518__CLK
timestamp 1667941163
transform 1 0 24840 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__519__CLK
timestamp 1667941163
transform 1 0 27876 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__520__CLK
timestamp 1667941163
transform 1 0 28428 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__520__D
timestamp 1667941163
transform -1 0 26956 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__521__CLK
timestamp 1667941163
transform 1 0 3036 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__522__CLK
timestamp 1667941163
transform 1 0 21988 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__523__CLK
timestamp 1667941163
transform 1 0 21988 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__524__CLK
timestamp 1667941163
transform 1 0 25116 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__525__CLK
timestamp 1667941163
transform 1 0 26496 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__526__CLK
timestamp 1667941163
transform 1 0 26220 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__527__CLK
timestamp 1667941163
transform 1 0 7820 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__528__CLK
timestamp 1667941163
transform 1 0 9108 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__529__CLK
timestamp 1667941163
transform 1 0 22632 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__542__A
timestamp 1667941163
transform 1 0 29624 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__543__A
timestamp 1667941163
transform -1 0 19504 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__544__A
timestamp 1667941163
transform -1 0 38272 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__545__A
timestamp 1667941163
transform -1 0 15548 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__546__A
timestamp 1667941163
transform -1 0 26680 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__548__A
timestamp 1667941163
transform -1 0 16744 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__549__A
timestamp 1667941163
transform -1 0 2576 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__550__A
timestamp 1667941163
transform -1 0 6072 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__551__A
timestamp 1667941163
transform -1 0 35052 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__552__A
timestamp 1667941163
transform 1 0 22816 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__554__A
timestamp 1667941163
transform 1 0 4876 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__555__A
timestamp 1667941163
transform 1 0 2392 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__556__A
timestamp 1667941163
transform -1 0 10120 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__557__A
timestamp 1667941163
transform -1 0 31740 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__558__A
timestamp 1667941163
transform -1 0 22172 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__559__A
timestamp 1667941163
transform 1 0 2760 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__560__A
timestamp 1667941163
transform 1 0 37260 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__561__A
timestamp 1667941163
transform -1 0 14444 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__562__A
timestamp 1667941163
transform -1 0 25208 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__563__A
timestamp 1667941163
transform 1 0 27232 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__564__A
timestamp 1667941163
transform 1 0 15180 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__565__A
timestamp 1667941163
transform 1 0 10764 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__566__A
timestamp 1667941163
transform -1 0 10488 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__567__A
timestamp 1667941163
transform 1 0 24196 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__569__A
timestamp 1667941163
transform 1 0 17756 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__570__A
timestamp 1667941163
transform -1 0 23460 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__571__A
timestamp 1667941163
transform -1 0 31556 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__574__A
timestamp 1667941163
transform -1 0 23184 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__575__A
timestamp 1667941163
transform 1 0 12696 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__576__A
timestamp 1667941163
transform -1 0 16928 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__577__A
timestamp 1667941163
transform 1 0 2668 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__578__A
timestamp 1667941163
transform -1 0 20332 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__613__A
timestamp 1667941163
transform 1 0 16192 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__619__A
timestamp 1667941163
transform -1 0 21528 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__621__A
timestamp 1667941163
transform 1 0 19136 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__628__A
timestamp 1667941163
transform -1 0 6808 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__691__A
timestamp 1667941163
transform 1 0 20424 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__693__A
timestamp 1667941163
transform 1 0 17756 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1667941163
transform -1 0 37628 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1667941163
transform 1 0 38180 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1667941163
transform -1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1667941163
transform -1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1667941163
transform -1 0 35144 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1667941163
transform -1 0 1748 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1667941163
transform -1 0 1748 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1667941163
transform -1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1667941163
transform -1 0 37628 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1667941163
transform -1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1667941163
transform -1 0 25852 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1667941163
transform -1 0 37628 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1667941163
transform -1 0 14536 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1667941163
transform -1 0 1748 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1667941163
transform -1 0 37628 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1667941163
transform -1 0 22172 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1667941163
transform -1 0 2300 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1667941163
transform -1 0 26588 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1667941163
transform -1 0 37628 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1667941163
transform -1 0 9384 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1667941163
transform -1 0 1748 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1667941163
transform -1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1667941163
transform -1 0 38364 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1667941163
transform -1 0 4600 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1667941163
transform -1 0 1748 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1667941163
transform -1 0 2484 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1667941163
transform -1 0 28060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1667941163
transform -1 0 1748 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1667941163
transform -1 0 25300 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1667941163
transform -1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1667941163
transform -1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1667941163
transform -1 0 33212 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1667941163
transform -1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1667941163
transform -1 0 37628 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1667941163
transform -1 0 1748 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1667941163
transform -1 0 3036 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1667941163
transform -1 0 36432 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1667941163
transform -1 0 1748 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1667941163
transform -1 0 37628 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1667941163
transform -1 0 31280 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output41_A
timestamp 1667941163
transform 1 0 37444 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output48_A
timestamp 1667941163
transform -1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output56_A
timestamp 1667941163
transform -1 0 26680 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output57_A
timestamp 1667941163
transform 1 0 34684 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output59_A
timestamp 1667941163
transform 1 0 37444 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output74_A
timestamp 1667941163
transform 1 0 2300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output75_A
timestamp 1667941163
transform -1 0 36984 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output79_A
timestamp 1667941163
transform -1 0 37628 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output88_A
timestamp 1667941163
transform -1 0 25852 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2668 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1667941163
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34
timestamp 1667941163
transform 1 0 4232 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4968 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1667941163
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63
timestamp 1667941163
transform 1 0 6900 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_75 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1667941163
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90
timestamp 1667941163
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_104
timestamp 1667941163
transform 1 0 10672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1667941163
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 12052 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_127
timestamp 1667941163
transform 1 0 12788 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_133
timestamp 1667941163
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1667941163
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1667941163
transform 1 0 14536 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154
timestamp 1667941163
transform 1 0 15272 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1667941163
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_175
timestamp 1667941163
transform 1 0 17204 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_183
timestamp 1667941163
transform 1 0 17940 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_189
timestamp 1667941163
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1667941163
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_205
timestamp 1667941163
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_210
timestamp 1667941163
transform 1 0 20424 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1667941163
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_231
timestamp 1667941163
transform 1 0 22356 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_239
timestamp 1667941163
transform 1 0 23092 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_245
timestamp 1667941163
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1667941163
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_261
timestamp 1667941163
transform 1 0 25116 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_266
timestamp 1667941163
transform 1 0 25576 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1667941163
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_287
timestamp 1667941163
transform 1 0 27508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_293
timestamp 1667941163
transform 1 0 28060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1667941163
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1667941163
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_315
timestamp 1667941163
transform 1 0 30084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_327
timestamp 1667941163
transform 1 0 31188 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_331
timestamp 1667941163
transform 1 0 31556 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_334
timestamp 1667941163
transform 1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_343
timestamp 1667941163
transform 1 0 32660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_349
timestamp 1667941163
transform 1 0 33212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_357
timestamp 1667941163
transform 1 0 33948 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1667941163
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_371
timestamp 1667941163
transform 1 0 35236 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_377
timestamp 1667941163
transform 1 0 35788 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_382
timestamp 1667941163
transform 1 0 36248 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1667941163
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_405
timestamp 1667941163
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1667941163
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1667941163
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_27
timestamp 1667941163
transform 1 0 3588 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_35
timestamp 1667941163
transform 1 0 4324 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_38
timestamp 1667941163
transform 1 0 4600 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_50
timestamp 1667941163
transform 1 0 5704 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_69
timestamp 1667941163
transform 1 0 7452 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_77
timestamp 1667941163
transform 1 0 8188 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_83
timestamp 1667941163
transform 1 0 8740 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_95
timestamp 1667941163
transform 1 0 9844 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_107
timestamp 1667941163
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1667941163
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_122
timestamp 1667941163
transform 1 0 12328 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_128
timestamp 1667941163
transform 1 0 12880 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_140
timestamp 1667941163
transform 1 0 13984 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_152
timestamp 1667941163
transform 1 0 15088 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1667941163
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_181
timestamp 1667941163
transform 1 0 17756 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_189
timestamp 1667941163
transform 1 0 18492 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_194
timestamp 1667941163
transform 1 0 18952 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_200
timestamp 1667941163
transform 1 0 19504 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_212
timestamp 1667941163
transform 1 0 20608 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1667941163
transform 1 0 20884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1667941163
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1667941163
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1667941163
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1667941163
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1667941163
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1667941163
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_293
timestamp 1667941163
transform 1 0 28060 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_301
timestamp 1667941163
transform 1 0 28796 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_306
timestamp 1667941163
transform 1 0 29256 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_312
timestamp 1667941163
transform 1 0 29808 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_324
timestamp 1667941163
transform 1 0 30912 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1667941163
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_361
timestamp 1667941163
transform 1 0 34316 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_367
timestamp 1667941163
transform 1 0 34868 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_379
timestamp 1667941163
transform 1 0 35972 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_384
timestamp 1667941163
transform 1 0 36432 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1667941163
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_397
timestamp 1667941163
transform 1 0 37628 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_9
timestamp 1667941163
transform 1 0 1932 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_21
timestamp 1667941163
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1667941163
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1667941163
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1667941163
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1667941163
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1667941163
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1667941163
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1667941163
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1667941163
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1667941163
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1667941163
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1667941163
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1667941163
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1667941163
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1667941163
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1667941163
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1667941163
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1667941163
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1667941163
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1667941163
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1667941163
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1667941163
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1667941163
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1667941163
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1667941163
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1667941163
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1667941163
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1667941163
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1667941163
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1667941163
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1667941163
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1667941163
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_389
timestamp 1667941163
transform 1 0 36892 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_397
timestamp 1667941163
transform 1 0 37628 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_405
timestamp 1667941163
transform 1 0 38364 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7
timestamp 1667941163
transform 1 0 1748 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_19
timestamp 1667941163
transform 1 0 2852 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_31
timestamp 1667941163
transform 1 0 3956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_43
timestamp 1667941163
transform 1 0 5060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1667941163
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1667941163
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1667941163
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1667941163
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1667941163
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1667941163
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1667941163
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1667941163
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1667941163
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1667941163
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1667941163
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1667941163
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1667941163
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1667941163
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1667941163
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1667941163
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1667941163
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1667941163
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1667941163
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1667941163
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1667941163
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1667941163
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1667941163
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1667941163
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1667941163
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1667941163
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1667941163
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1667941163
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1667941163
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1667941163
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_401
timestamp 1667941163
transform 1 0 37996 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7
timestamp 1667941163
transform 1 0 1748 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_19
timestamp 1667941163
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1667941163
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1667941163
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1667941163
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1667941163
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1667941163
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1667941163
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1667941163
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1667941163
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1667941163
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1667941163
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1667941163
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1667941163
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1667941163
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1667941163
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1667941163
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1667941163
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1667941163
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1667941163
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1667941163
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1667941163
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1667941163
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1667941163
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1667941163
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1667941163
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1667941163
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1667941163
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1667941163
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1667941163
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1667941163
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1667941163
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1667941163
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_401
timestamp 1667941163
transform 1 0 37996 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_9
timestamp 1667941163
transform 1 0 1932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_21
timestamp 1667941163
transform 1 0 3036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_33
timestamp 1667941163
transform 1 0 4140 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_45
timestamp 1667941163
transform 1 0 5244 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1667941163
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1667941163
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1667941163
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1667941163
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1667941163
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1667941163
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1667941163
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1667941163
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1667941163
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1667941163
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1667941163
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1667941163
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1667941163
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1667941163
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1667941163
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1667941163
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1667941163
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1667941163
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1667941163
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1667941163
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1667941163
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1667941163
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1667941163
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1667941163
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1667941163
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1667941163
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1667941163
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1667941163
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1667941163
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1667941163
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1667941163
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1667941163
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1667941163
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1667941163
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1667941163
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1667941163
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1667941163
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1667941163
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1667941163
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1667941163
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1667941163
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1667941163
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1667941163
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1667941163
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1667941163
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1667941163
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1667941163
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1667941163
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1667941163
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1667941163
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1667941163
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1667941163
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1667941163
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1667941163
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1667941163
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1667941163
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1667941163
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1667941163
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1667941163
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1667941163
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1667941163
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1667941163
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1667941163
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1667941163
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1667941163
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_389
timestamp 1667941163
transform 1 0 36892 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_397
timestamp 1667941163
transform 1 0 37628 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_405
timestamp 1667941163
transform 1 0 38364 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1667941163
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1667941163
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1667941163
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1667941163
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1667941163
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1667941163
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1667941163
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1667941163
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1667941163
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1667941163
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1667941163
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1667941163
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1667941163
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1667941163
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1667941163
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1667941163
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1667941163
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1667941163
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1667941163
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1667941163
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1667941163
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_249
timestamp 1667941163
transform 1 0 24012 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_256
timestamp 1667941163
transform 1 0 24656 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_262
timestamp 1667941163
transform 1 0 25208 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_274
timestamp 1667941163
transform 1 0 26312 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1667941163
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1667941163
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1667941163
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1667941163
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1667941163
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1667941163
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1667941163
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1667941163
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1667941163
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1667941163
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7
timestamp 1667941163
transform 1 0 1748 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_19
timestamp 1667941163
transform 1 0 2852 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1667941163
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1667941163
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1667941163
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1667941163
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1667941163
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1667941163
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1667941163
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1667941163
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1667941163
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1667941163
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1667941163
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1667941163
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1667941163
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1667941163
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1667941163
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1667941163
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1667941163
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1667941163
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1667941163
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1667941163
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1667941163
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1667941163
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1667941163
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1667941163
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1667941163
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1667941163
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1667941163
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1667941163
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1667941163
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1667941163
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1667941163
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1667941163
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_401
timestamp 1667941163
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1667941163
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1667941163
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1667941163
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1667941163
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1667941163
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1667941163
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1667941163
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1667941163
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1667941163
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1667941163
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1667941163
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1667941163
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1667941163
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1667941163
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1667941163
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1667941163
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1667941163
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1667941163
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1667941163
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1667941163
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_234
timestamp 1667941163
transform 1 0 22632 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_240
timestamp 1667941163
transform 1 0 23184 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_252
timestamp 1667941163
transform 1 0 24288 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_264
timestamp 1667941163
transform 1 0 25392 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 1667941163
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1667941163
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1667941163
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1667941163
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1667941163
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1667941163
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1667941163
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1667941163
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1667941163
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1667941163
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_397
timestamp 1667941163
transform 1 0 37628 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1667941163
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1667941163
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1667941163
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1667941163
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1667941163
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1667941163
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1667941163
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1667941163
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1667941163
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1667941163
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1667941163
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1667941163
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1667941163
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1667941163
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1667941163
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1667941163
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1667941163
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1667941163
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1667941163
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1667941163
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1667941163
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1667941163
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1667941163
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1667941163
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1667941163
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1667941163
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1667941163
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1667941163
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1667941163
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1667941163
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1667941163
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1667941163
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1667941163
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_401
timestamp 1667941163
transform 1 0 37996 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_7
timestamp 1667941163
transform 1 0 1748 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_19
timestamp 1667941163
transform 1 0 2852 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_31
timestamp 1667941163
transform 1 0 3956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_43
timestamp 1667941163
transform 1 0 5060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1667941163
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1667941163
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1667941163
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1667941163
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1667941163
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1667941163
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1667941163
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1667941163
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1667941163
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1667941163
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1667941163
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1667941163
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1667941163
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1667941163
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1667941163
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1667941163
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1667941163
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1667941163
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1667941163
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1667941163
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1667941163
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1667941163
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1667941163
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1667941163
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1667941163
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1667941163
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1667941163
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1667941163
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1667941163
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_9
timestamp 1667941163
transform 1 0 1932 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_21
timestamp 1667941163
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1667941163
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1667941163
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1667941163
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1667941163
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1667941163
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1667941163
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1667941163
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1667941163
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1667941163
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1667941163
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1667941163
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_147
timestamp 1667941163
transform 1 0 14628 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_151
timestamp 1667941163
transform 1 0 14996 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_157
timestamp 1667941163
transform 1 0 15548 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_166
timestamp 1667941163
transform 1 0 16376 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_172
timestamp 1667941163
transform 1 0 16928 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_184
timestamp 1667941163
transform 1 0 18032 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1667941163
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1667941163
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1667941163
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1667941163
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1667941163
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1667941163
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1667941163
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1667941163
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1667941163
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1667941163
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1667941163
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1667941163
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1667941163
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1667941163
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1667941163
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1667941163
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_405
timestamp 1667941163
transform 1 0 38364 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1667941163
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1667941163
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1667941163
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1667941163
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1667941163
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1667941163
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1667941163
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1667941163
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1667941163
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1667941163
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1667941163
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1667941163
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1667941163
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1667941163
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1667941163
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1667941163
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1667941163
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1667941163
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1667941163
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1667941163
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1667941163
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1667941163
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1667941163
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1667941163
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1667941163
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1667941163
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1667941163
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1667941163
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1667941163
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1667941163
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1667941163
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1667941163
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1667941163
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1667941163
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1667941163
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1667941163
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1667941163
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1667941163
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1667941163
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1667941163
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1667941163
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1667941163
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1667941163
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1667941163
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1667941163
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1667941163
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_153
timestamp 1667941163
transform 1 0 15180 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_161
timestamp 1667941163
transform 1 0 15916 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_166
timestamp 1667941163
transform 1 0 16376 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_172
timestamp 1667941163
transform 1 0 16928 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_184
timestamp 1667941163
transform 1 0 18032 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1667941163
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1667941163
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1667941163
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1667941163
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1667941163
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1667941163
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1667941163
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1667941163
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1667941163
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1667941163
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1667941163
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1667941163
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1667941163
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1667941163
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1667941163
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1667941163
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_401
timestamp 1667941163
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_9
timestamp 1667941163
transform 1 0 1932 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_21
timestamp 1667941163
transform 1 0 3036 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_33
timestamp 1667941163
transform 1 0 4140 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_45
timestamp 1667941163
transform 1 0 5244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1667941163
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1667941163
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_81
timestamp 1667941163
transform 1 0 8556 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_87
timestamp 1667941163
transform 1 0 9108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_99
timestamp 1667941163
transform 1 0 10212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1667941163
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1667941163
transform 1 0 11960 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_124
timestamp 1667941163
transform 1 0 12512 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_136
timestamp 1667941163
transform 1 0 13616 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_148
timestamp 1667941163
transform 1 0 14720 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_160
timestamp 1667941163
transform 1 0 15824 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1667941163
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_193
timestamp 1667941163
transform 1 0 18860 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_197
timestamp 1667941163
transform 1 0 19228 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_203
timestamp 1667941163
transform 1 0 19780 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_215
timestamp 1667941163
transform 1 0 20884 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1667941163
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1667941163
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1667941163
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_261
timestamp 1667941163
transform 1 0 25116 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_266
timestamp 1667941163
transform 1 0 25576 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_272
timestamp 1667941163
transform 1 0 26128 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1667941163
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1667941163
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1667941163
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1667941163
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1667941163
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1667941163
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1667941163
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1667941163
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1667941163
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1667941163
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1667941163
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1667941163
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1667941163
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1667941163
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1667941163
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1667941163
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_97
timestamp 1667941163
transform 1 0 10028 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_108
timestamp 1667941163
transform 1 0 11040 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_114
timestamp 1667941163
transform 1 0 11592 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_126
timestamp 1667941163
transform 1 0 12696 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1667941163
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1667941163
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1667941163
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1667941163
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1667941163
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1667941163
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1667941163
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1667941163
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1667941163
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1667941163
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1667941163
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1667941163
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1667941163
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1667941163
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1667941163
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1667941163
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1667941163
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1667941163
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1667941163
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1667941163
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_389
timestamp 1667941163
transform 1 0 36892 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_397
timestamp 1667941163
transform 1 0 37628 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_405
timestamp 1667941163
transform 1 0 38364 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1667941163
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1667941163
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1667941163
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1667941163
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1667941163
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1667941163
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1667941163
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1667941163
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1667941163
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1667941163
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1667941163
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1667941163
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1667941163
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1667941163
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1667941163
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1667941163
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1667941163
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1667941163
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1667941163
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1667941163
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1667941163
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1667941163
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1667941163
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1667941163
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1667941163
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1667941163
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1667941163
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1667941163
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1667941163
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1667941163
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1667941163
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1667941163
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1667941163
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1667941163
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1667941163
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1667941163
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1667941163
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1667941163
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1667941163
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1667941163
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1667941163
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1667941163
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1667941163
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1667941163
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1667941163
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1667941163
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1667941163
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_153
timestamp 1667941163
transform 1 0 15180 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_159
timestamp 1667941163
transform 1 0 15732 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1667941163
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1667941163
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1667941163
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1667941163
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1667941163
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1667941163
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1667941163
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1667941163
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1667941163
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1667941163
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1667941163
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1667941163
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1667941163
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1667941163
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1667941163
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1667941163
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1667941163
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1667941163
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1667941163
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_389
timestamp 1667941163
transform 1 0 36892 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_397
timestamp 1667941163
transform 1 0 37628 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_402
timestamp 1667941163
transform 1 0 38088 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_406
timestamp 1667941163
transform 1 0 38456 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_9
timestamp 1667941163
transform 1 0 1932 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_21
timestamp 1667941163
transform 1 0 3036 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_33
timestamp 1667941163
transform 1 0 4140 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_45
timestamp 1667941163
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1667941163
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1667941163
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1667941163
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1667941163
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1667941163
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1667941163
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1667941163
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1667941163
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1667941163
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1667941163
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1667941163
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1667941163
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1667941163
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1667941163
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1667941163
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1667941163
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1667941163
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1667941163
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1667941163
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1667941163
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1667941163
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1667941163
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1667941163
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1667941163
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1667941163
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1667941163
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1667941163
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1667941163
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1667941163
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1667941163
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_397
timestamp 1667941163
transform 1 0 37628 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1667941163
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_7
timestamp 1667941163
transform 1 0 1748 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_19
timestamp 1667941163
transform 1 0 2852 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1667941163
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1667941163
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1667941163
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1667941163
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1667941163
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1667941163
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1667941163
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1667941163
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1667941163
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1667941163
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1667941163
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1667941163
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1667941163
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1667941163
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1667941163
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1667941163
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1667941163
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1667941163
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1667941163
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1667941163
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1667941163
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1667941163
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1667941163
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1667941163
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1667941163
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1667941163
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1667941163
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1667941163
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1667941163
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1667941163
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1667941163
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_401
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_9
timestamp 1667941163
transform 1 0 1932 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_16
timestamp 1667941163
transform 1 0 2576 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_28
timestamp 1667941163
transform 1 0 3680 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_40
timestamp 1667941163
transform 1 0 4784 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1667941163
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1667941163
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1667941163
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1667941163
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1667941163
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1667941163
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1667941163
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1667941163
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1667941163
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1667941163
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1667941163
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1667941163
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1667941163
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1667941163
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1667941163
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1667941163
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1667941163
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1667941163
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1667941163
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1667941163
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1667941163
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1667941163
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1667941163
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1667941163
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1667941163
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1667941163
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1667941163
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1667941163
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_401
timestamp 1667941163
transform 1 0 37996 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_10
timestamp 1667941163
transform 1 0 2024 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_16
timestamp 1667941163
transform 1 0 2576 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1667941163
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1667941163
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1667941163
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1667941163
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1667941163
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1667941163
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1667941163
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1667941163
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1667941163
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1667941163
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1667941163
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1667941163
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1667941163
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1667941163
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1667941163
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1667941163
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1667941163
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1667941163
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1667941163
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1667941163
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1667941163
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1667941163
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1667941163
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1667941163
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1667941163
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1667941163
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1667941163
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1667941163
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1667941163
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1667941163
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1667941163
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_389
timestamp 1667941163
transform 1 0 36892 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_405
timestamp 1667941163
transform 1 0 38364 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1667941163
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1667941163
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1667941163
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1667941163
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1667941163
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1667941163
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1667941163
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1667941163
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1667941163
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1667941163
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1667941163
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1667941163
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1667941163
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1667941163
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1667941163
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1667941163
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1667941163
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1667941163
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1667941163
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1667941163
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1667941163
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1667941163
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1667941163
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1667941163
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1667941163
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1667941163
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1667941163
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1667941163
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1667941163
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1667941163
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1667941163
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1667941163
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1667941163
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1667941163
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1667941163
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1667941163
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1667941163
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1667941163
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_53
timestamp 1667941163
transform 1 0 5980 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_61
timestamp 1667941163
transform 1 0 6716 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_66
timestamp 1667941163
transform 1 0 7176 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_78
timestamp 1667941163
transform 1 0 8280 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1667941163
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1667941163
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1667941163
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1667941163
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1667941163
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1667941163
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1667941163
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1667941163
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1667941163
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1667941163
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1667941163
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1667941163
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1667941163
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1667941163
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1667941163
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1667941163
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1667941163
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1667941163
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1667941163
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1667941163
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1667941163
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1667941163
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1667941163
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1667941163
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1667941163
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1667941163
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_401
timestamp 1667941163
transform 1 0 37996 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_405
timestamp 1667941163
transform 1 0 38364 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_9
timestamp 1667941163
transform 1 0 1932 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_21
timestamp 1667941163
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_33
timestamp 1667941163
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1667941163
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1667941163
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1667941163
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1667941163
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1667941163
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1667941163
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1667941163
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1667941163
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1667941163
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1667941163
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1667941163
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1667941163
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1667941163
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1667941163
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1667941163
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1667941163
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1667941163
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1667941163
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1667941163
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1667941163
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1667941163
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1667941163
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1667941163
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1667941163
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1667941163
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1667941163
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1667941163
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1667941163
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1667941163
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1667941163
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1667941163
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1667941163
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1667941163
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1667941163
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1667941163
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1667941163
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1667941163
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1667941163
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1667941163
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1667941163
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1667941163
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1667941163
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1667941163
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1667941163
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1667941163
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1667941163
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1667941163
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1667941163
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1667941163
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1667941163
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1667941163
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1667941163
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1667941163
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1667941163
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1667941163
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1667941163
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1667941163
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1667941163
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1667941163
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1667941163
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1667941163
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1667941163
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1667941163
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1667941163
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1667941163
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_401
timestamp 1667941163
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1667941163
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1667941163
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1667941163
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1667941163
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1667941163
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_63
timestamp 1667941163
transform 1 0 6900 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_75
timestamp 1667941163
transform 1 0 8004 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_87
timestamp 1667941163
transform 1 0 9108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_99
timestamp 1667941163
transform 1 0 10212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1667941163
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1667941163
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1667941163
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1667941163
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1667941163
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1667941163
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1667941163
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_193
timestamp 1667941163
transform 1 0 18860 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_201
timestamp 1667941163
transform 1 0 19596 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_205
timestamp 1667941163
transform 1 0 19964 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_211
timestamp 1667941163
transform 1 0 20516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1667941163
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1667941163
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1667941163
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1667941163
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1667941163
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1667941163
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1667941163
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1667941163
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1667941163
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1667941163
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1667941163
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1667941163
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1667941163
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1667941163
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1667941163
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1667941163
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1667941163
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1667941163
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1667941163
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1667941163
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1667941163
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1667941163
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1667941163
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1667941163
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1667941163
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1667941163
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1667941163
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1667941163
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1667941163
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1667941163
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1667941163
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1667941163
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1667941163
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1667941163
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1667941163
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1667941163
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1667941163
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1667941163
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1667941163
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1667941163
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1667941163
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1667941163
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1667941163
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1667941163
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1667941163
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1667941163
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1667941163
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1667941163
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1667941163
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1667941163
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1667941163
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_9
timestamp 1667941163
transform 1 0 1932 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_21
timestamp 1667941163
transform 1 0 3036 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_33
timestamp 1667941163
transform 1 0 4140 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_45
timestamp 1667941163
transform 1 0 5244 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp 1667941163
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1667941163
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1667941163
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1667941163
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1667941163
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1667941163
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1667941163
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1667941163
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1667941163
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1667941163
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1667941163
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1667941163
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1667941163
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1667941163
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1667941163
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1667941163
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1667941163
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1667941163
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1667941163
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1667941163
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1667941163
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1667941163
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_305
timestamp 1667941163
transform 1 0 29164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_309
timestamp 1667941163
transform 1 0 29532 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_321
timestamp 1667941163
transform 1 0 30636 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_333
timestamp 1667941163
transform 1 0 31740 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1667941163
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1667941163
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1667941163
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1667941163
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1667941163
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_7
timestamp 1667941163
transform 1 0 1748 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_13
timestamp 1667941163
transform 1 0 2300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_25
timestamp 1667941163
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_33
timestamp 1667941163
transform 1 0 4140 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_37
timestamp 1667941163
transform 1 0 4508 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_43
timestamp 1667941163
transform 1 0 5060 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_55
timestamp 1667941163
transform 1 0 6164 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_67
timestamp 1667941163
transform 1 0 7268 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_79
timestamp 1667941163
transform 1 0 8372 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1667941163
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1667941163
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1667941163
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1667941163
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_133
timestamp 1667941163
transform 1 0 13340 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_137
timestamp 1667941163
transform 1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1667941163
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1667941163
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1667941163
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1667941163
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1667941163
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_202
timestamp 1667941163
transform 1 0 19688 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_208
timestamp 1667941163
transform 1 0 20240 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_220
timestamp 1667941163
transform 1 0 21344 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_232
timestamp 1667941163
transform 1 0 22448 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_244
timestamp 1667941163
transform 1 0 23552 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1667941163
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1667941163
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1667941163
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1667941163
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1667941163
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1667941163
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1667941163
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1667941163
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1667941163
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1667941163
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1667941163
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1667941163
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_401
timestamp 1667941163
transform 1 0 37996 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_9
timestamp 1667941163
transform 1 0 1932 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_15
timestamp 1667941163
transform 1 0 2484 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_21
timestamp 1667941163
transform 1 0 3036 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_33
timestamp 1667941163
transform 1 0 4140 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_45
timestamp 1667941163
transform 1 0 5244 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1667941163
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1667941163
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1667941163
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1667941163
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1667941163
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_117
timestamp 1667941163
transform 1 0 11868 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_120
timestamp 1667941163
transform 1 0 12144 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_128
timestamp 1667941163
transform 1 0 12880 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_134
timestamp 1667941163
transform 1 0 13432 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_138
timestamp 1667941163
transform 1 0 13800 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_141
timestamp 1667941163
transform 1 0 14076 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_145
timestamp 1667941163
transform 1 0 14444 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_149
timestamp 1667941163
transform 1 0 14812 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_155
timestamp 1667941163
transform 1 0 15364 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_163
timestamp 1667941163
transform 1 0 16100 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1667941163
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1667941163
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1667941163
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1667941163
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1667941163
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1667941163
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1667941163
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1667941163
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1667941163
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1667941163
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1667941163
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1667941163
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1667941163
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1667941163
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1667941163
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1667941163
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1667941163
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1667941163
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1667941163
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1667941163
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1667941163
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_401
timestamp 1667941163
transform 1 0 37996 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1667941163
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_7
timestamp 1667941163
transform 1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_11
timestamp 1667941163
transform 1 0 2116 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_14
timestamp 1667941163
transform 1 0 2392 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_20
timestamp 1667941163
transform 1 0 2944 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1667941163
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_33
timestamp 1667941163
transform 1 0 4140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_45
timestamp 1667941163
transform 1 0 5244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_57
timestamp 1667941163
transform 1 0 6348 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_69
timestamp 1667941163
transform 1 0 7452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_81
timestamp 1667941163
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_97
timestamp 1667941163
transform 1 0 10028 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_105
timestamp 1667941163
transform 1 0 10764 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_111
timestamp 1667941163
transform 1 0 11316 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_119
timestamp 1667941163
transform 1 0 12052 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_123
timestamp 1667941163
transform 1 0 12420 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_127
timestamp 1667941163
transform 1 0 12788 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_131
timestamp 1667941163
transform 1 0 13156 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1667941163
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_146
timestamp 1667941163
transform 1 0 14536 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_154
timestamp 1667941163
transform 1 0 15272 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_164
timestamp 1667941163
transform 1 0 16192 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_170
timestamp 1667941163
transform 1 0 16744 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_182
timestamp 1667941163
transform 1 0 17848 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1667941163
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1667941163
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1667941163
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1667941163
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1667941163
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1667941163
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1667941163
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1667941163
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1667941163
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1667941163
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1667941163
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1667941163
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1667941163
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1667941163
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1667941163
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1667941163
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_389
timestamp 1667941163
transform 1 0 36892 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_405
timestamp 1667941163
transform 1 0 38364 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_7
timestamp 1667941163
transform 1 0 1748 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_13
timestamp 1667941163
transform 1 0 2300 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_19
timestamp 1667941163
transform 1 0 2852 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_25
timestamp 1667941163
transform 1 0 3404 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_28
timestamp 1667941163
transform 1 0 3680 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_34
timestamp 1667941163
transform 1 0 4232 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_40
timestamp 1667941163
transform 1 0 4784 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_46
timestamp 1667941163
transform 1 0 5336 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1667941163
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1667941163
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1667941163
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_93
timestamp 1667941163
transform 1 0 9660 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_96
timestamp 1667941163
transform 1 0 9936 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_103
timestamp 1667941163
transform 1 0 10580 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1667941163
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_124
timestamp 1667941163
transform 1 0 12512 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_133
timestamp 1667941163
transform 1 0 13340 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_140
timestamp 1667941163
transform 1 0 13984 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_152
timestamp 1667941163
transform 1 0 15088 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1667941163
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_173
timestamp 1667941163
transform 1 0 17020 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_185
timestamp 1667941163
transform 1 0 18124 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_197
timestamp 1667941163
transform 1 0 19228 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_209
timestamp 1667941163
transform 1 0 20332 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_221
timestamp 1667941163
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1667941163
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1667941163
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1667941163
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1667941163
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1667941163
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1667941163
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1667941163
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1667941163
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1667941163
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1667941163
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1667941163
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1667941163
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1667941163
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1667941163
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1667941163
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_7
timestamp 1667941163
transform 1 0 1748 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_15
timestamp 1667941163
transform 1 0 2484 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_18
timestamp 1667941163
transform 1 0 2760 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_24
timestamp 1667941163
transform 1 0 3312 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_33
timestamp 1667941163
transform 1 0 4140 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_39
timestamp 1667941163
transform 1 0 4692 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_45
timestamp 1667941163
transform 1 0 5244 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_51
timestamp 1667941163
transform 1 0 5796 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_63
timestamp 1667941163
transform 1 0 6900 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_75
timestamp 1667941163
transform 1 0 8004 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1667941163
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_97
timestamp 1667941163
transform 1 0 10028 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_102
timestamp 1667941163
transform 1 0 10488 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_109
timestamp 1667941163
transform 1 0 11132 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_116
timestamp 1667941163
transform 1 0 11776 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_124
timestamp 1667941163
transform 1 0 12512 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1667941163
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_152
timestamp 1667941163
transform 1 0 15088 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_160
timestamp 1667941163
transform 1 0 15824 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_171
timestamp 1667941163
transform 1 0 16836 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_178
timestamp 1667941163
transform 1 0 17480 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_184
timestamp 1667941163
transform 1 0 18032 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1667941163
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1667941163
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1667941163
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1667941163
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1667941163
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1667941163
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1667941163
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1667941163
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1667941163
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1667941163
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1667941163
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1667941163
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1667941163
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1667941163
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1667941163
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1667941163
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_401
timestamp 1667941163
transform 1 0 37996 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_9
timestamp 1667941163
transform 1 0 1932 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_15
timestamp 1667941163
transform 1 0 2484 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_25
timestamp 1667941163
transform 1 0 3404 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_31
timestamp 1667941163
transform 1 0 3956 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_37
timestamp 1667941163
transform 1 0 4508 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_43
timestamp 1667941163
transform 1 0 5060 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_49
timestamp 1667941163
transform 1 0 5612 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_52
timestamp 1667941163
transform 1 0 5888 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_61
timestamp 1667941163
transform 1 0 6716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_73
timestamp 1667941163
transform 1 0 7820 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_85
timestamp 1667941163
transform 1 0 8924 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_89
timestamp 1667941163
transform 1 0 9292 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_92
timestamp 1667941163
transform 1 0 9568 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_98
timestamp 1667941163
transform 1 0 10120 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1667941163
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_119
timestamp 1667941163
transform 1 0 12052 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_128
timestamp 1667941163
transform 1 0 12880 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_137
timestamp 1667941163
transform 1 0 13708 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_145
timestamp 1667941163
transform 1 0 14444 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1667941163
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1667941163
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_179
timestamp 1667941163
transform 1 0 17572 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_191
timestamp 1667941163
transform 1 0 18676 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_203
timestamp 1667941163
transform 1 0 19780 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_215
timestamp 1667941163
transform 1 0 20884 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1667941163
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1667941163
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1667941163
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1667941163
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1667941163
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1667941163
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1667941163
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1667941163
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1667941163
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1667941163
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1667941163
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1667941163
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1667941163
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1667941163
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1667941163
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1667941163
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_7
timestamp 1667941163
transform 1 0 1748 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_13
timestamp 1667941163
transform 1 0 2300 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_17
timestamp 1667941163
transform 1 0 2668 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_20
timestamp 1667941163
transform 1 0 2944 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1667941163
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_33
timestamp 1667941163
transform 1 0 4140 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_39
timestamp 1667941163
transform 1 0 4692 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_45
timestamp 1667941163
transform 1 0 5244 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_51
timestamp 1667941163
transform 1 0 5796 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_54
timestamp 1667941163
transform 1 0 6072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_60
timestamp 1667941163
transform 1 0 6624 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_66
timestamp 1667941163
transform 1 0 7176 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_72
timestamp 1667941163
transform 1 0 7728 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1667941163
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_89
timestamp 1667941163
transform 1 0 9292 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_93
timestamp 1667941163
transform 1 0 9660 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_106
timestamp 1667941163
transform 1 0 10856 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_119
timestamp 1667941163
transform 1 0 12052 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1667941163
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1667941163
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_145
timestamp 1667941163
transform 1 0 14444 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_154
timestamp 1667941163
transform 1 0 15272 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_161
timestamp 1667941163
transform 1 0 15916 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_168
timestamp 1667941163
transform 1 0 16560 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_174
timestamp 1667941163
transform 1 0 17112 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_180
timestamp 1667941163
transform 1 0 17664 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_183
timestamp 1667941163
transform 1 0 17940 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1667941163
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1667941163
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1667941163
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1667941163
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1667941163
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1667941163
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1667941163
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1667941163
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1667941163
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1667941163
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1667941163
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1667941163
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1667941163
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1667941163
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1667941163
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1667941163
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1667941163
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1667941163
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1667941163
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_401
timestamp 1667941163
transform 1 0 37996 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_9
timestamp 1667941163
transform 1 0 1932 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_15
timestamp 1667941163
transform 1 0 2484 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_18
timestamp 1667941163
transform 1 0 2760 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_24
timestamp 1667941163
transform 1 0 3312 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_27
timestamp 1667941163
transform 1 0 3588 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_33
timestamp 1667941163
transform 1 0 4140 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_39
timestamp 1667941163
transform 1 0 4692 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_42
timestamp 1667941163
transform 1 0 4968 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_48
timestamp 1667941163
transform 1 0 5520 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1667941163
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_61
timestamp 1667941163
transform 1 0 6716 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_65
timestamp 1667941163
transform 1 0 7084 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_68
timestamp 1667941163
transform 1 0 7360 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_74
timestamp 1667941163
transform 1 0 7912 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_81
timestamp 1667941163
transform 1 0 8556 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_88
timestamp 1667941163
transform 1 0 9200 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_95
timestamp 1667941163
transform 1 0 9844 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_102
timestamp 1667941163
transform 1 0 10488 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1667941163
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_123
timestamp 1667941163
transform 1 0 12420 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_136
timestamp 1667941163
transform 1 0 13616 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_149
timestamp 1667941163
transform 1 0 14812 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1667941163
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1667941163
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_181
timestamp 1667941163
transform 1 0 17756 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_190
timestamp 1667941163
transform 1 0 18584 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_203
timestamp 1667941163
transform 1 0 19780 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_215
timestamp 1667941163
transform 1 0 20884 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1667941163
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1667941163
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1667941163
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1667941163
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1667941163
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1667941163
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1667941163
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1667941163
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1667941163
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1667941163
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1667941163
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1667941163
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1667941163
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1667941163
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1667941163
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1667941163
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_10
timestamp 1667941163
transform 1 0 2024 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_16
timestamp 1667941163
transform 1 0 2576 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_22
timestamp 1667941163
transform 1 0 3128 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_33
timestamp 1667941163
transform 1 0 4140 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_39
timestamp 1667941163
transform 1 0 4692 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_45
timestamp 1667941163
transform 1 0 5244 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_51
timestamp 1667941163
transform 1 0 5796 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_59
timestamp 1667941163
transform 1 0 6532 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_62
timestamp 1667941163
transform 1 0 6808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_68
timestamp 1667941163
transform 1 0 7360 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_75
timestamp 1667941163
transform 1 0 8004 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1667941163
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_91
timestamp 1667941163
transform 1 0 9476 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_95
timestamp 1667941163
transform 1 0 9844 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_108
timestamp 1667941163
transform 1 0 11040 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_115
timestamp 1667941163
transform 1 0 11684 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_127
timestamp 1667941163
transform 1 0 12788 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_131
timestamp 1667941163
transform 1 0 13156 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_135
timestamp 1667941163
transform 1 0 13524 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1667941163
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_152
timestamp 1667941163
transform 1 0 15088 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_160
timestamp 1667941163
transform 1 0 15824 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_170
timestamp 1667941163
transform 1 0 16744 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_177
timestamp 1667941163
transform 1 0 17388 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_183
timestamp 1667941163
transform 1 0 17940 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1667941163
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1667941163
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1667941163
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1667941163
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1667941163
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1667941163
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1667941163
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1667941163
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_277
timestamp 1667941163
transform 1 0 26588 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_283
timestamp 1667941163
transform 1 0 27140 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_286
timestamp 1667941163
transform 1 0 27416 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_294
timestamp 1667941163
transform 1 0 28152 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_306
timestamp 1667941163
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1667941163
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1667941163
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1667941163
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1667941163
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1667941163
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1667941163
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1667941163
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 1667941163
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_7
timestamp 1667941163
transform 1 0 1748 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_11
timestamp 1667941163
transform 1 0 2116 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_17
timestamp 1667941163
transform 1 0 2668 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_25
timestamp 1667941163
transform 1 0 3404 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_33
timestamp 1667941163
transform 1 0 4140 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_36
timestamp 1667941163
transform 1 0 4416 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_44
timestamp 1667941163
transform 1 0 5152 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1667941163
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_61
timestamp 1667941163
transform 1 0 6716 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_68
timestamp 1667941163
transform 1 0 7360 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_75
timestamp 1667941163
transform 1 0 8004 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_82
timestamp 1667941163
transform 1 0 8648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_94
timestamp 1667941163
transform 1 0 9752 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_39_109
timestamp 1667941163
transform 1 0 11132 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_123
timestamp 1667941163
transform 1 0 12420 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_131
timestamp 1667941163
transform 1 0 13156 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_141
timestamp 1667941163
transform 1 0 14076 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_148
timestamp 1667941163
transform 1 0 14720 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1667941163
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1667941163
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_174
timestamp 1667941163
transform 1 0 17112 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_182
timestamp 1667941163
transform 1 0 17848 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_192
timestamp 1667941163
transform 1 0 18768 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_198
timestamp 1667941163
transform 1 0 19320 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_204
timestamp 1667941163
transform 1 0 19872 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_216
timestamp 1667941163
transform 1 0 20976 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1667941163
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1667941163
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1667941163
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1667941163
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1667941163
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1667941163
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1667941163
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1667941163
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1667941163
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1667941163
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1667941163
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1667941163
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1667941163
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1667941163
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1667941163
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_7
timestamp 1667941163
transform 1 0 1748 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_11
timestamp 1667941163
transform 1 0 2116 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_18
timestamp 1667941163
transform 1 0 2760 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_24
timestamp 1667941163
transform 1 0 3312 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_33
timestamp 1667941163
transform 1 0 4140 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_39
timestamp 1667941163
transform 1 0 4692 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_42
timestamp 1667941163
transform 1 0 4968 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_48
timestamp 1667941163
transform 1 0 5520 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_54
timestamp 1667941163
transform 1 0 6072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_61
timestamp 1667941163
transform 1 0 6716 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_68
timestamp 1667941163
transform 1 0 7360 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_75
timestamp 1667941163
transform 1 0 8004 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1667941163
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_96
timestamp 1667941163
transform 1 0 9936 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_112
timestamp 1667941163
transform 1 0 11408 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_120
timestamp 1667941163
transform 1 0 12144 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_129
timestamp 1667941163
transform 1 0 12972 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1667941163
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_147
timestamp 1667941163
transform 1 0 14628 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_153
timestamp 1667941163
transform 1 0 15180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_166
timestamp 1667941163
transform 1 0 16376 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_173
timestamp 1667941163
transform 1 0 17020 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_180
timestamp 1667941163
transform 1 0 17664 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_186
timestamp 1667941163
transform 1 0 18216 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_193
timestamp 1667941163
transform 1 0 18860 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_203
timestamp 1667941163
transform 1 0 19780 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1667941163
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1667941163
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1667941163
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1667941163
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1667941163
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1667941163
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1667941163
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1667941163
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1667941163
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1667941163
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1667941163
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1667941163
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1667941163
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1667941163
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1667941163
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1667941163
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1667941163
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_401
timestamp 1667941163
transform 1 0 37996 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_9
timestamp 1667941163
transform 1 0 1932 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_16
timestamp 1667941163
transform 1 0 2576 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_23
timestamp 1667941163
transform 1 0 3220 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_30
timestamp 1667941163
transform 1 0 3864 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_38
timestamp 1667941163
transform 1 0 4600 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_41
timestamp 1667941163
transform 1 0 4876 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_47
timestamp 1667941163
transform 1 0 5428 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_54
timestamp 1667941163
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_62
timestamp 1667941163
transform 1 0 6808 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_69
timestamp 1667941163
transform 1 0 7452 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_76
timestamp 1667941163
transform 1 0 8096 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_83
timestamp 1667941163
transform 1 0 8740 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_95
timestamp 1667941163
transform 1 0 9844 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1667941163
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_119
timestamp 1667941163
transform 1 0 12052 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_129
timestamp 1667941163
transform 1 0 12972 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_133
timestamp 1667941163
transform 1 0 13340 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_137
timestamp 1667941163
transform 1 0 13708 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_149
timestamp 1667941163
transform 1 0 14812 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1667941163
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_174
timestamp 1667941163
transform 1 0 17112 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_182
timestamp 1667941163
transform 1 0 17848 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_186
timestamp 1667941163
transform 1 0 18216 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_193
timestamp 1667941163
transform 1 0 18860 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_206
timestamp 1667941163
transform 1 0 20056 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_212
timestamp 1667941163
transform 1 0 20608 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1667941163
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1667941163
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1667941163
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1667941163
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1667941163
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1667941163
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1667941163
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1667941163
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1667941163
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1667941163
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1667941163
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1667941163
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1667941163
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1667941163
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1667941163
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_7
timestamp 1667941163
transform 1 0 1748 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_11
timestamp 1667941163
transform 1 0 2116 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_18
timestamp 1667941163
transform 1 0 2760 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_25
timestamp 1667941163
transform 1 0 3404 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_34
timestamp 1667941163
transform 1 0 4232 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_43
timestamp 1667941163
transform 1 0 5060 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_50
timestamp 1667941163
transform 1 0 5704 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_57
timestamp 1667941163
transform 1 0 6348 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_64
timestamp 1667941163
transform 1 0 6992 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_76
timestamp 1667941163
transform 1 0 8096 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1667941163
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_91
timestamp 1667941163
transform 1 0 9476 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_101
timestamp 1667941163
transform 1 0 10396 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_107
timestamp 1667941163
transform 1 0 10948 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_119
timestamp 1667941163
transform 1 0 12052 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_132
timestamp 1667941163
transform 1 0 13248 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1667941163
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_152
timestamp 1667941163
transform 1 0 15088 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_158
timestamp 1667941163
transform 1 0 15640 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_167
timestamp 1667941163
transform 1 0 16468 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_174
timestamp 1667941163
transform 1 0 17112 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_181
timestamp 1667941163
transform 1 0 17756 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1667941163
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_212
timestamp 1667941163
transform 1 0 20608 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_219
timestamp 1667941163
transform 1 0 21252 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_225
timestamp 1667941163
transform 1 0 21804 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_237
timestamp 1667941163
transform 1 0 22908 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_249
timestamp 1667941163
transform 1 0 24012 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1667941163
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1667941163
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_289
timestamp 1667941163
transform 1 0 27692 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_295
timestamp 1667941163
transform 1 0 28244 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_299
timestamp 1667941163
transform 1 0 28612 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1667941163
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_314
timestamp 1667941163
transform 1 0 29992 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_326
timestamp 1667941163
transform 1 0 31096 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_338
timestamp 1667941163
transform 1 0 32200 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_350
timestamp 1667941163
transform 1 0 33304 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_362
timestamp 1667941163
transform 1 0 34408 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_389
timestamp 1667941163
transform 1 0 36892 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_397
timestamp 1667941163
transform 1 0 37628 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_402
timestamp 1667941163
transform 1 0 38088 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_406
timestamp 1667941163
transform 1 0 38456 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_7
timestamp 1667941163
transform 1 0 1748 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_11
timestamp 1667941163
transform 1 0 2116 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_18
timestamp 1667941163
transform 1 0 2760 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_25
timestamp 1667941163
transform 1 0 3404 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_34
timestamp 1667941163
transform 1 0 4232 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_40
timestamp 1667941163
transform 1 0 4784 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_47
timestamp 1667941163
transform 1 0 5428 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_54
timestamp 1667941163
transform 1 0 6072 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_63
timestamp 1667941163
transform 1 0 6900 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_76
timestamp 1667941163
transform 1 0 8096 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_89
timestamp 1667941163
transform 1 0 9292 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_102
timestamp 1667941163
transform 1 0 10488 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_106
timestamp 1667941163
transform 1 0 10856 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1667941163
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_120
timestamp 1667941163
transform 1 0 12144 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_133
timestamp 1667941163
transform 1 0 13340 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_145
timestamp 1667941163
transform 1 0 14444 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_152
timestamp 1667941163
transform 1 0 15088 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_159
timestamp 1667941163
transform 1 0 15732 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_166
timestamp 1667941163
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_173
timestamp 1667941163
transform 1 0 17020 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_177
timestamp 1667941163
transform 1 0 17388 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_189
timestamp 1667941163
transform 1 0 18492 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_198
timestamp 1667941163
transform 1 0 19320 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_212
timestamp 1667941163
transform 1 0 20608 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_219
timestamp 1667941163
transform 1 0 21252 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1667941163
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_229
timestamp 1667941163
transform 1 0 22172 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_235
timestamp 1667941163
transform 1 0 22724 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_247
timestamp 1667941163
transform 1 0 23828 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_259
timestamp 1667941163
transform 1 0 24932 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_271
timestamp 1667941163
transform 1 0 26036 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1667941163
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1667941163
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1667941163
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1667941163
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1667941163
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1667941163
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1667941163
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1667941163
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1667941163
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1667941163
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_402
timestamp 1667941163
transform 1 0 38088 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_406
timestamp 1667941163
transform 1 0 38456 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_7
timestamp 1667941163
transform 1 0 1748 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_11
timestamp 1667941163
transform 1 0 2116 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_18
timestamp 1667941163
transform 1 0 2760 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_22
timestamp 1667941163
transform 1 0 3128 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_26
timestamp 1667941163
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_34
timestamp 1667941163
transform 1 0 4232 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_48
timestamp 1667941163
transform 1 0 5520 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_55
timestamp 1667941163
transform 1 0 6164 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_62
timestamp 1667941163
transform 1 0 6808 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_69
timestamp 1667941163
transform 1 0 7452 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_82
timestamp 1667941163
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_99
timestamp 1667941163
transform 1 0 10212 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_111
timestamp 1667941163
transform 1 0 11316 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_123
timestamp 1667941163
transform 1 0 12420 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1667941163
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_145
timestamp 1667941163
transform 1 0 14444 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_157
timestamp 1667941163
transform 1 0 15548 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_164
timestamp 1667941163
transform 1 0 16192 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_175
timestamp 1667941163
transform 1 0 17204 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_182
timestamp 1667941163
transform 1 0 17848 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1667941163
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_44_208
timestamp 1667941163
transform 1 0 20240 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_216
timestamp 1667941163
transform 1 0 20976 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_222
timestamp 1667941163
transform 1 0 21528 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_228
timestamp 1667941163
transform 1 0 22080 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_240
timestamp 1667941163
transform 1 0 23184 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1667941163
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1667941163
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1667941163
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1667941163
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1667941163
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_314
timestamp 1667941163
transform 1 0 29992 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_321
timestamp 1667941163
transform 1 0 30636 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_327
timestamp 1667941163
transform 1 0 31188 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_339
timestamp 1667941163
transform 1 0 32292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_351
timestamp 1667941163
transform 1 0 33396 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1667941163
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1667941163
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1667941163
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_401
timestamp 1667941163
transform 1 0 37996 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_404
timestamp 1667941163
transform 1 0 38272 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_9
timestamp 1667941163
transform 1 0 1932 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_16
timestamp 1667941163
transform 1 0 2576 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_23
timestamp 1667941163
transform 1 0 3220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_29
timestamp 1667941163
transform 1 0 3772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_33
timestamp 1667941163
transform 1 0 4140 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_40
timestamp 1667941163
transform 1 0 4784 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_47
timestamp 1667941163
transform 1 0 5428 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1667941163
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_61
timestamp 1667941163
transform 1 0 6716 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_65
timestamp 1667941163
transform 1 0 7084 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_78
timestamp 1667941163
transform 1 0 8280 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_95
timestamp 1667941163
transform 1 0 9844 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_108
timestamp 1667941163
transform 1 0 11040 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_128
timestamp 1667941163
transform 1 0 12880 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_134
timestamp 1667941163
transform 1 0 13432 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_138
timestamp 1667941163
transform 1 0 13800 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_151
timestamp 1667941163
transform 1 0 14996 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_158
timestamp 1667941163
transform 1 0 15640 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_162
timestamp 1667941163
transform 1 0 16008 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1667941163
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_180
timestamp 1667941163
transform 1 0 17664 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_189
timestamp 1667941163
transform 1 0 18492 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_202
timestamp 1667941163
transform 1 0 19688 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_211
timestamp 1667941163
transform 1 0 20516 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1667941163
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1667941163
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_229
timestamp 1667941163
transform 1 0 22172 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_235
timestamp 1667941163
transform 1 0 22724 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_243
timestamp 1667941163
transform 1 0 23460 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_247
timestamp 1667941163
transform 1 0 23828 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_253
timestamp 1667941163
transform 1 0 24380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_265
timestamp 1667941163
transform 1 0 25484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_277
timestamp 1667941163
transform 1 0 26588 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1667941163
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1667941163
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1667941163
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1667941163
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1667941163
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1667941163
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1667941163
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1667941163
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1667941163
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1667941163
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_397
timestamp 1667941163
transform 1 0 37628 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1667941163
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_7
timestamp 1667941163
transform 1 0 1748 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_11
timestamp 1667941163
transform 1 0 2116 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_15
timestamp 1667941163
transform 1 0 2484 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_19
timestamp 1667941163
transform 1 0 2852 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_26
timestamp 1667941163
transform 1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_33
timestamp 1667941163
transform 1 0 4140 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_40
timestamp 1667941163
transform 1 0 4784 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_47
timestamp 1667941163
transform 1 0 5428 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_54
timestamp 1667941163
transform 1 0 6072 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_61
timestamp 1667941163
transform 1 0 6716 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_68
timestamp 1667941163
transform 1 0 7360 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_75
timestamp 1667941163
transform 1 0 8004 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_82
timestamp 1667941163
transform 1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_95
timestamp 1667941163
transform 1 0 9844 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_112
timestamp 1667941163
transform 1 0 11408 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_131
timestamp 1667941163
transform 1 0 13156 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1667941163
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_145
timestamp 1667941163
transform 1 0 14444 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_155
timestamp 1667941163
transform 1 0 15364 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_172
timestamp 1667941163
transform 1 0 16928 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_178
timestamp 1667941163
transform 1 0 17480 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_182
timestamp 1667941163
transform 1 0 17848 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1667941163
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_203
timestamp 1667941163
transform 1 0 19780 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_213
timestamp 1667941163
transform 1 0 20700 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_220
timestamp 1667941163
transform 1 0 21344 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_226
timestamp 1667941163
transform 1 0 21896 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_232
timestamp 1667941163
transform 1 0 22448 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_238
timestamp 1667941163
transform 1 0 23000 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_250
timestamp 1667941163
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_258
timestamp 1667941163
transform 1 0 24840 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_264
timestamp 1667941163
transform 1 0 25392 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_276
timestamp 1667941163
transform 1 0 26496 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_288
timestamp 1667941163
transform 1 0 27600 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_300
timestamp 1667941163
transform 1 0 28704 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1667941163
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1667941163
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1667941163
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1667941163
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1667941163
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1667941163
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_401
timestamp 1667941163
transform 1 0 37996 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_9
timestamp 1667941163
transform 1 0 1932 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_18
timestamp 1667941163
transform 1 0 2760 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_25
timestamp 1667941163
transform 1 0 3404 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_32
timestamp 1667941163
transform 1 0 4048 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_40
timestamp 1667941163
transform 1 0 4784 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_47
timestamp 1667941163
transform 1 0 5428 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_54
timestamp 1667941163
transform 1 0 6072 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_66
timestamp 1667941163
transform 1 0 7176 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_79
timestamp 1667941163
transform 1 0 8372 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_87
timestamp 1667941163
transform 1 0 9108 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_97
timestamp 1667941163
transform 1 0 10028 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_110
timestamp 1667941163
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_122
timestamp 1667941163
transform 1 0 12328 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_135
timestamp 1667941163
transform 1 0 13524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_150
timestamp 1667941163
transform 1 0 14904 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_157
timestamp 1667941163
transform 1 0 15548 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_166
timestamp 1667941163
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_180
timestamp 1667941163
transform 1 0 17664 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_184
timestamp 1667941163
transform 1 0 18032 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_188
timestamp 1667941163
transform 1 0 18400 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_201
timestamp 1667941163
transform 1 0 19596 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_213
timestamp 1667941163
transform 1 0 20700 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_219
timestamp 1667941163
transform 1 0 21252 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1667941163
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_229
timestamp 1667941163
transform 1 0 22172 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_241
timestamp 1667941163
transform 1 0 23276 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_253
timestamp 1667941163
transform 1 0 24380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_265
timestamp 1667941163
transform 1 0 25484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_277
timestamp 1667941163
transform 1 0 26588 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1667941163
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1667941163
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1667941163
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1667941163
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1667941163
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1667941163
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1667941163
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1667941163
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1667941163
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1667941163
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1667941163
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_12
timestamp 1667941163
transform 1 0 2208 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_19
timestamp 1667941163
transform 1 0 2852 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_26
timestamp 1667941163
transform 1 0 3496 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_40
timestamp 1667941163
transform 1 0 4784 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_46
timestamp 1667941163
transform 1 0 5336 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_60
timestamp 1667941163
transform 1 0 6624 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_69
timestamp 1667941163
transform 1 0 7452 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_82
timestamp 1667941163
transform 1 0 8648 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_98
timestamp 1667941163
transform 1 0 10120 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_115
timestamp 1667941163
transform 1 0 11684 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_136
timestamp 1667941163
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_152
timestamp 1667941163
transform 1 0 15088 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_167
timestamp 1667941163
transform 1 0 16468 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_180
timestamp 1667941163
transform 1 0 17664 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_184
timestamp 1667941163
transform 1 0 18032 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_194
timestamp 1667941163
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_202
timestamp 1667941163
transform 1 0 19688 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_209
timestamp 1667941163
transform 1 0 20332 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_216
timestamp 1667941163
transform 1 0 20976 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_222
timestamp 1667941163
transform 1 0 21528 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_234
timestamp 1667941163
transform 1 0 22632 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_246
timestamp 1667941163
transform 1 0 23736 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1667941163
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1667941163
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1667941163
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1667941163
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1667941163
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_321
timestamp 1667941163
transform 1 0 30636 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_325
timestamp 1667941163
transform 1 0 31004 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_331
timestamp 1667941163
transform 1 0 31556 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_343
timestamp 1667941163
transform 1 0 32660 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_355
timestamp 1667941163
transform 1 0 33764 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_360
timestamp 1667941163
transform 1 0 34224 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_369
timestamp 1667941163
transform 1 0 35052 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_381
timestamp 1667941163
transform 1 0 36156 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_393
timestamp 1667941163
transform 1 0 37260 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_405
timestamp 1667941163
transform 1 0 38364 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_9
timestamp 1667941163
transform 1 0 1932 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_15
timestamp 1667941163
transform 1 0 2484 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_19
timestamp 1667941163
transform 1 0 2852 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_43
timestamp 1667941163
transform 1 0 5060 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_54
timestamp 1667941163
transform 1 0 6072 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_71
timestamp 1667941163
transform 1 0 7636 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_84
timestamp 1667941163
transform 1 0 8832 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_97
timestamp 1667941163
transform 1 0 10028 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_110
timestamp 1667941163
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_135
timestamp 1667941163
transform 1 0 13524 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_139
timestamp 1667941163
transform 1 0 13892 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_149
timestamp 1667941163
transform 1 0 14812 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_162
timestamp 1667941163
transform 1 0 16008 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_181
timestamp 1667941163
transform 1 0 17756 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_194
timestamp 1667941163
transform 1 0 18952 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_198
timestamp 1667941163
transform 1 0 19320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_202
timestamp 1667941163
transform 1 0 19688 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_209
timestamp 1667941163
transform 1 0 20332 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_216
timestamp 1667941163
transform 1 0 20976 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 1667941163
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_229
timestamp 1667941163
transform 1 0 22172 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_241
timestamp 1667941163
transform 1 0 23276 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_253
timestamp 1667941163
transform 1 0 24380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_265
timestamp 1667941163
transform 1 0 25484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_277
timestamp 1667941163
transform 1 0 26588 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1667941163
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1667941163
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1667941163
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1667941163
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1667941163
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1667941163
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1667941163
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1667941163
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_26
timestamp 1667941163
transform 1 0 3496 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_51
timestamp 1667941163
transform 1 0 5796 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_59
timestamp 1667941163
transform 1 0 6532 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_81
timestamp 1667941163
transform 1 0 8556 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_96
timestamp 1667941163
transform 1 0 9936 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_102
timestamp 1667941163
transform 1 0 10488 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_124
timestamp 1667941163
transform 1 0 12512 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_50_137
timestamp 1667941163
transform 1 0 13708 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_158
timestamp 1667941163
transform 1 0 15640 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_50_175
timestamp 1667941163
transform 1 0 17204 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_183
timestamp 1667941163
transform 1 0 17940 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_193
timestamp 1667941163
transform 1 0 18860 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_202
timestamp 1667941163
transform 1 0 19688 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_209
timestamp 1667941163
transform 1 0 20332 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_216
timestamp 1667941163
transform 1 0 20976 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_222
timestamp 1667941163
transform 1 0 21528 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_228
timestamp 1667941163
transform 1 0 22080 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_234
timestamp 1667941163
transform 1 0 22632 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_246
timestamp 1667941163
transform 1 0 23736 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1667941163
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1667941163
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1667941163
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1667941163
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1667941163
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1667941163
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1667941163
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1667941163
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1667941163
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1667941163
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1667941163
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_389
timestamp 1667941163
transform 1 0 36892 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_395
timestamp 1667941163
transform 1 0 37444 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_402
timestamp 1667941163
transform 1 0 38088 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_406
timestamp 1667941163
transform 1 0 38456 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_26
timestamp 1667941163
transform 1 0 3496 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_50
timestamp 1667941163
transform 1 0 5704 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_63
timestamp 1667941163
transform 1 0 6900 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_85
timestamp 1667941163
transform 1 0 8924 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1667941163
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_135
timestamp 1667941163
transform 1 0 13524 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_143
timestamp 1667941163
transform 1 0 14260 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_153
timestamp 1667941163
transform 1 0 15180 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1667941163
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_180
timestamp 1667941163
transform 1 0 17664 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_187
timestamp 1667941163
transform 1 0 18308 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_191
timestamp 1667941163
transform 1 0 18676 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_195
timestamp 1667941163
transform 1 0 19044 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_202
timestamp 1667941163
transform 1 0 19688 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_209
timestamp 1667941163
transform 1 0 20332 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_215
timestamp 1667941163
transform 1 0 20884 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_51_221
timestamp 1667941163
transform 1 0 21436 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_229
timestamp 1667941163
transform 1 0 22172 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_235
timestamp 1667941163
transform 1 0 22724 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_247
timestamp 1667941163
transform 1 0 23828 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_259
timestamp 1667941163
transform 1 0 24932 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_271
timestamp 1667941163
transform 1 0 26036 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1667941163
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1667941163
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_305
timestamp 1667941163
transform 1 0 29164 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_310
timestamp 1667941163
transform 1 0 29624 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_316
timestamp 1667941163
transform 1 0 30176 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_328
timestamp 1667941163
transform 1 0 31280 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1667941163
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1667941163
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1667941163
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1667941163
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1667941163
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_26
timestamp 1667941163
transform 1 0 3496 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_54
timestamp 1667941163
transform 1 0 6072 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_58
timestamp 1667941163
transform 1 0 6440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_82
timestamp 1667941163
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_89
timestamp 1667941163
transform 1 0 9292 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_96
timestamp 1667941163
transform 1 0 9936 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_103
timestamp 1667941163
transform 1 0 10580 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_130
timestamp 1667941163
transform 1 0 13064 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_134
timestamp 1667941163
transform 1 0 13432 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1667941163
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_146
timestamp 1667941163
transform 1 0 14536 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_159
timestamp 1667941163
transform 1 0 15732 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_172
timestamp 1667941163
transform 1 0 16928 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_185
timestamp 1667941163
transform 1 0 18124 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_193
timestamp 1667941163
transform 1 0 18860 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_202
timestamp 1667941163
transform 1 0 19688 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_209
timestamp 1667941163
transform 1 0 20332 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_215
timestamp 1667941163
transform 1 0 20884 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_226
timestamp 1667941163
transform 1 0 21896 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1667941163
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1667941163
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1667941163
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1667941163
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1667941163
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1667941163
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1667941163
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1667941163
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_321
timestamp 1667941163
transform 1 0 30636 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_327
timestamp 1667941163
transform 1 0 31188 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1667941163
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1667941163
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1667941163
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1667941163
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1667941163
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1667941163
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_401
timestamp 1667941163
transform 1 0 37996 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_9
timestamp 1667941163
transform 1 0 1932 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_16
timestamp 1667941163
transform 1 0 2576 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_43
timestamp 1667941163
transform 1 0 5060 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_54
timestamp 1667941163
transform 1 0 6072 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_64
timestamp 1667941163
transform 1 0 6992 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_91
timestamp 1667941163
transform 1 0 9476 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_99
timestamp 1667941163
transform 1 0 10212 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_103
timestamp 1667941163
transform 1 0 10580 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 1667941163
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_136
timestamp 1667941163
transform 1 0 13616 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_145
timestamp 1667941163
transform 1 0 14444 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_158
timestamp 1667941163
transform 1 0 15640 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_165
timestamp 1667941163
transform 1 0 16284 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_173
timestamp 1667941163
transform 1 0 17020 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_183
timestamp 1667941163
transform 1 0 17940 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_196
timestamp 1667941163
transform 1 0 19136 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_203
timestamp 1667941163
transform 1 0 19780 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_210
timestamp 1667941163
transform 1 0 20424 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1667941163
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1667941163
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_229
timestamp 1667941163
transform 1 0 22172 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_235
timestamp 1667941163
transform 1 0 22724 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_241
timestamp 1667941163
transform 1 0 23276 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_253
timestamp 1667941163
transform 1 0 24380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_265
timestamp 1667941163
transform 1 0 25484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_277
timestamp 1667941163
transform 1 0 26588 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1667941163
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1667941163
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1667941163
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1667941163
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1667941163
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1667941163
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1667941163
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1667941163
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1667941163
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1667941163
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1667941163
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_26
timestamp 1667941163
transform 1 0 3496 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_35
timestamp 1667941163
transform 1 0 4324 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_42
timestamp 1667941163
transform 1 0 4968 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_69
timestamp 1667941163
transform 1 0 7452 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_75
timestamp 1667941163
transform 1 0 8004 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_82
timestamp 1667941163
transform 1 0 8648 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_89
timestamp 1667941163
transform 1 0 9292 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_93
timestamp 1667941163
transform 1 0 9660 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_100
timestamp 1667941163
transform 1 0 10304 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_125
timestamp 1667941163
transform 1 0 12604 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_131
timestamp 1667941163
transform 1 0 13156 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_138
timestamp 1667941163
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_146
timestamp 1667941163
transform 1 0 14536 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_161
timestamp 1667941163
transform 1 0 15916 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_174
timestamp 1667941163
transform 1 0 17112 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_187
timestamp 1667941163
transform 1 0 18308 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_194
timestamp 1667941163
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_202
timestamp 1667941163
transform 1 0 19688 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_209
timestamp 1667941163
transform 1 0 20332 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_220
timestamp 1667941163
transform 1 0 21344 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_226
timestamp 1667941163
transform 1 0 21896 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_232
timestamp 1667941163
transform 1 0 22448 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_238
timestamp 1667941163
transform 1 0 23000 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_244
timestamp 1667941163
transform 1 0 23552 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1667941163
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1667941163
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1667941163
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1667941163
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1667941163
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1667941163
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1667941163
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1667941163
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1667941163
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1667941163
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_401
timestamp 1667941163
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_9
timestamp 1667941163
transform 1 0 1932 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_17
timestamp 1667941163
transform 1 0 2668 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_23
timestamp 1667941163
transform 1 0 3220 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_48
timestamp 1667941163
transform 1 0 5520 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_54
timestamp 1667941163
transform 1 0 6072 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_84
timestamp 1667941163
transform 1 0 8832 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_110
timestamp 1667941163
transform 1 0 11224 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_136
timestamp 1667941163
transform 1 0 13616 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1667941163
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1667941163
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_180
timestamp 1667941163
transform 1 0 17664 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_195
timestamp 1667941163
transform 1 0 19044 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_202
timestamp 1667941163
transform 1 0 19688 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_209
timestamp 1667941163
transform 1 0 20332 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_215
timestamp 1667941163
transform 1 0 20884 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_221
timestamp 1667941163
transform 1 0 21436 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_230
timestamp 1667941163
transform 1 0 22264 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_236
timestamp 1667941163
transform 1 0 22816 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_242
timestamp 1667941163
transform 1 0 23368 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_248
timestamp 1667941163
transform 1 0 23920 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_254
timestamp 1667941163
transform 1 0 24472 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_266
timestamp 1667941163
transform 1 0 25576 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_278
timestamp 1667941163
transform 1 0 26680 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1667941163
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1667941163
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1667941163
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1667941163
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1667941163
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1667941163
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1667941163
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1667941163
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1667941163
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1667941163
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_26
timestamp 1667941163
transform 1 0 3496 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_33
timestamp 1667941163
transform 1 0 4140 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_37
timestamp 1667941163
transform 1 0 4508 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_64
timestamp 1667941163
transform 1 0 6992 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_56_73
timestamp 1667941163
transform 1 0 7820 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_82
timestamp 1667941163
transform 1 0 8648 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_90
timestamp 1667941163
transform 1 0 9384 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_94
timestamp 1667941163
transform 1 0 9752 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_98
timestamp 1667941163
transform 1 0 10120 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_102
timestamp 1667941163
transform 1 0 10488 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_106
timestamp 1667941163
transform 1 0 10856 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1667941163
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1667941163
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_145
timestamp 1667941163
transform 1 0 14444 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_158
timestamp 1667941163
transform 1 0 15640 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_166
timestamp 1667941163
transform 1 0 16376 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_180
timestamp 1667941163
transform 1 0 17664 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_186
timestamp 1667941163
transform 1 0 18216 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_190
timestamp 1667941163
transform 1 0 18584 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_202
timestamp 1667941163
transform 1 0 19688 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_208
timestamp 1667941163
transform 1 0 20240 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_214
timestamp 1667941163
transform 1 0 20792 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_222
timestamp 1667941163
transform 1 0 21528 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_226
timestamp 1667941163
transform 1 0 21896 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_232
timestamp 1667941163
transform 1 0 22448 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_238
timestamp 1667941163
transform 1 0 23000 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_244
timestamp 1667941163
transform 1 0 23552 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1667941163
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_257
timestamp 1667941163
transform 1 0 24748 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_263
timestamp 1667941163
transform 1 0 25300 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_269
timestamp 1667941163
transform 1 0 25852 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_281
timestamp 1667941163
transform 1 0 26956 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_293
timestamp 1667941163
transform 1 0 28060 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_305
timestamp 1667941163
transform 1 0 29164 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1667941163
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1667941163
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1667941163
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1667941163
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1667941163
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_401
timestamp 1667941163
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_15
timestamp 1667941163
transform 1 0 2484 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_23
timestamp 1667941163
transform 1 0 3220 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_27
timestamp 1667941163
transform 1 0 3588 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_49
timestamp 1667941163
transform 1 0 5612 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1667941163
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_63
timestamp 1667941163
transform 1 0 6900 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_85
timestamp 1667941163
transform 1 0 8924 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_110
timestamp 1667941163
transform 1 0 11224 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_138
timestamp 1667941163
transform 1 0 13800 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_144
timestamp 1667941163
transform 1 0 14352 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_148
timestamp 1667941163
transform 1 0 14720 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_165
timestamp 1667941163
transform 1 0 16284 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_174
timestamp 1667941163
transform 1 0 17112 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_182
timestamp 1667941163
transform 1 0 17848 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_186
timestamp 1667941163
transform 1 0 18216 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_195
timestamp 1667941163
transform 1 0 19044 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_202
timestamp 1667941163
transform 1 0 19688 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_213
timestamp 1667941163
transform 1 0 20700 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_219
timestamp 1667941163
transform 1 0 21252 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1667941163
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_229
timestamp 1667941163
transform 1 0 22172 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_235
timestamp 1667941163
transform 1 0 22724 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_241
timestamp 1667941163
transform 1 0 23276 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_247
timestamp 1667941163
transform 1 0 23828 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_253
timestamp 1667941163
transform 1 0 24380 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_259
timestamp 1667941163
transform 1 0 24932 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_265
timestamp 1667941163
transform 1 0 25484 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_271
timestamp 1667941163
transform 1 0 26036 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_57_277
timestamp 1667941163
transform 1 0 26588 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1667941163
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1667941163
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1667941163
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1667941163
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1667941163
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1667941163
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1667941163
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_397
timestamp 1667941163
transform 1 0 37628 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_26
timestamp 1667941163
transform 1 0 3496 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_34
timestamp 1667941163
transform 1 0 4232 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_42
timestamp 1667941163
transform 1 0 4968 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_69
timestamp 1667941163
transform 1 0 7452 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_76
timestamp 1667941163
transform 1 0 8096 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_82
timestamp 1667941163
transform 1 0 8648 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_90
timestamp 1667941163
transform 1 0 9384 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_96
timestamp 1667941163
transform 1 0 9936 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_121
timestamp 1667941163
transform 1 0 12236 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_129
timestamp 1667941163
transform 1 0 12972 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1667941163
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1667941163
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_150
timestamp 1667941163
transform 1 0 14904 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_163
timestamp 1667941163
transform 1 0 16100 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_169
timestamp 1667941163
transform 1 0 16652 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_176
timestamp 1667941163
transform 1 0 17296 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_193
timestamp 1667941163
transform 1 0 18860 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_201
timestamp 1667941163
transform 1 0 19596 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_211
timestamp 1667941163
transform 1 0 20516 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_217
timestamp 1667941163
transform 1 0 21068 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_223
timestamp 1667941163
transform 1 0 21620 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_229
timestamp 1667941163
transform 1 0 22172 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_235
timestamp 1667941163
transform 1 0 22724 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_241
timestamp 1667941163
transform 1 0 23276 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_247
timestamp 1667941163
transform 1 0 23828 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1667941163
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_257
timestamp 1667941163
transform 1 0 24748 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_263
timestamp 1667941163
transform 1 0 25300 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_269
timestamp 1667941163
transform 1 0 25852 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_275
timestamp 1667941163
transform 1 0 26404 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_287
timestamp 1667941163
transform 1 0 27508 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_299
timestamp 1667941163
transform 1 0 28612 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1667941163
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1667941163
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1667941163
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1667941163
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1667941163
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1667941163
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1667941163
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1667941163
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 1667941163
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_9
timestamp 1667941163
transform 1 0 1932 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_20
timestamp 1667941163
transform 1 0 2944 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_59_49
timestamp 1667941163
transform 1 0 5612 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1667941163
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_62
timestamp 1667941163
transform 1 0 6808 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_89
timestamp 1667941163
transform 1 0 9292 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_96
timestamp 1667941163
transform 1 0 9936 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_103
timestamp 1667941163
transform 1 0 10580 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_110
timestamp 1667941163
transform 1 0 11224 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_135
timestamp 1667941163
transform 1 0 13524 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_142
timestamp 1667941163
transform 1 0 14168 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_146
timestamp 1667941163
transform 1 0 14536 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_150
timestamp 1667941163
transform 1 0 14904 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_154
timestamp 1667941163
transform 1 0 15272 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_158
timestamp 1667941163
transform 1 0 15640 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_165
timestamp 1667941163
transform 1 0 16284 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_180
timestamp 1667941163
transform 1 0 17664 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_184
timestamp 1667941163
transform 1 0 18032 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_188
timestamp 1667941163
transform 1 0 18400 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_195
timestamp 1667941163
transform 1 0 19044 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_203
timestamp 1667941163
transform 1 0 19780 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_210
timestamp 1667941163
transform 1 0 20424 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_216
timestamp 1667941163
transform 1 0 20976 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_222
timestamp 1667941163
transform 1 0 21528 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_229
timestamp 1667941163
transform 1 0 22172 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_235
timestamp 1667941163
transform 1 0 22724 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_241
timestamp 1667941163
transform 1 0 23276 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_247
timestamp 1667941163
transform 1 0 23828 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_253
timestamp 1667941163
transform 1 0 24380 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_259
timestamp 1667941163
transform 1 0 24932 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_265
timestamp 1667941163
transform 1 0 25484 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_271
timestamp 1667941163
transform 1 0 26036 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_277
timestamp 1667941163
transform 1 0 26588 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_285
timestamp 1667941163
transform 1 0 27324 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_297
timestamp 1667941163
transform 1 0 28428 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_309
timestamp 1667941163
transform 1 0 29532 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_321
timestamp 1667941163
transform 1 0 30636 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_333
timestamp 1667941163
transform 1 0 31740 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1667941163
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1667941163
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1667941163
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1667941163
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1667941163
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_26
timestamp 1667941163
transform 1 0 3496 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_34
timestamp 1667941163
transform 1 0 4232 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_58
timestamp 1667941163
transform 1 0 6440 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_82
timestamp 1667941163
transform 1 0 8648 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_103
timestamp 1667941163
transform 1 0 10580 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_125
timestamp 1667941163
transform 1 0 12604 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1667941163
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1667941163
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_145
timestamp 1667941163
transform 1 0 14444 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_152
timestamp 1667941163
transform 1 0 15088 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_159
timestamp 1667941163
transform 1 0 15732 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_166
timestamp 1667941163
transform 1 0 16376 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_174
timestamp 1667941163
transform 1 0 17112 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_178
timestamp 1667941163
transform 1 0 17480 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_185
timestamp 1667941163
transform 1 0 18124 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_60_194
timestamp 1667941163
transform 1 0 18952 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_203
timestamp 1667941163
transform 1 0 19780 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_210
timestamp 1667941163
transform 1 0 20424 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_220
timestamp 1667941163
transform 1 0 21344 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_226
timestamp 1667941163
transform 1 0 21896 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_232
timestamp 1667941163
transform 1 0 22448 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_238
timestamp 1667941163
transform 1 0 23000 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_244
timestamp 1667941163
transform 1 0 23552 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 1667941163
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_257
timestamp 1667941163
transform 1 0 24748 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_263
timestamp 1667941163
transform 1 0 25300 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_269
timestamp 1667941163
transform 1 0 25852 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_275
timestamp 1667941163
transform 1 0 26404 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_281
timestamp 1667941163
transform 1 0 26956 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_287
timestamp 1667941163
transform 1 0 27508 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_293
timestamp 1667941163
transform 1 0 28060 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_305
timestamp 1667941163
transform 1 0 29164 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1667941163
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1667941163
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1667941163
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1667941163
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1667941163
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1667941163
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1667941163
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_401
timestamp 1667941163
transform 1 0 37996 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_9
timestamp 1667941163
transform 1 0 1932 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_30
timestamp 1667941163
transform 1 0 3864 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1667941163
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_61
timestamp 1667941163
transform 1 0 6716 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_66
timestamp 1667941163
transform 1 0 7176 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_135
timestamp 1667941163
transform 1 0 13524 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_159
timestamp 1667941163
transform 1 0 15732 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_166
timestamp 1667941163
transform 1 0 16376 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_174
timestamp 1667941163
transform 1 0 17112 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_182
timestamp 1667941163
transform 1 0 17848 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_186
timestamp 1667941163
transform 1 0 18216 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_193
timestamp 1667941163
transform 1 0 18860 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_199
timestamp 1667941163
transform 1 0 19412 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_203
timestamp 1667941163
transform 1 0 19780 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_210
timestamp 1667941163
transform 1 0 20424 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1667941163
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1667941163
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_230
timestamp 1667941163
transform 1 0 22264 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_236
timestamp 1667941163
transform 1 0 22816 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_242
timestamp 1667941163
transform 1 0 23368 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_248
timestamp 1667941163
transform 1 0 23920 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_254
timestamp 1667941163
transform 1 0 24472 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_260
timestamp 1667941163
transform 1 0 25024 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_266
timestamp 1667941163
transform 1 0 25576 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_272
timestamp 1667941163
transform 1 0 26128 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_278
timestamp 1667941163
transform 1 0 26680 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_285
timestamp 1667941163
transform 1 0 27324 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_291
timestamp 1667941163
transform 1 0 27876 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_297
timestamp 1667941163
transform 1 0 28428 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_303
timestamp 1667941163
transform 1 0 28980 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_315
timestamp 1667941163
transform 1 0 30084 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_327
timestamp 1667941163
transform 1 0 31188 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1667941163
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1667941163
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1667941163
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1667941163
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1667941163
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1667941163
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_397
timestamp 1667941163
transform 1 0 37628 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_26
timestamp 1667941163
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_34
timestamp 1667941163
transform 1 0 4232 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_58
timestamp 1667941163
transform 1 0 6440 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_82
timestamp 1667941163
transform 1 0 8648 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_107
timestamp 1667941163
transform 1 0 10948 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_131
timestamp 1667941163
transform 1 0 13156 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_138
timestamp 1667941163
transform 1 0 13800 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_163
timestamp 1667941163
transform 1 0 16100 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_167
timestamp 1667941163
transform 1 0 16468 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_171
timestamp 1667941163
transform 1 0 16836 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_178
timestamp 1667941163
transform 1 0 17480 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_185
timestamp 1667941163
transform 1 0 18124 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_62_194
timestamp 1667941163
transform 1 0 18952 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_202
timestamp 1667941163
transform 1 0 19688 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_212
timestamp 1667941163
transform 1 0 20608 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_220
timestamp 1667941163
transform 1 0 21344 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_224
timestamp 1667941163
transform 1 0 21712 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_237
timestamp 1667941163
transform 1 0 22908 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_243
timestamp 1667941163
transform 1 0 23460 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_249
timestamp 1667941163
transform 1 0 24012 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_257
timestamp 1667941163
transform 1 0 24748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_263
timestamp 1667941163
transform 1 0 25300 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_269
timestamp 1667941163
transform 1 0 25852 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_275
timestamp 1667941163
transform 1 0 26404 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_281
timestamp 1667941163
transform 1 0 26956 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_287
timestamp 1667941163
transform 1 0 27508 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_293
timestamp 1667941163
transform 1 0 28060 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_299
timestamp 1667941163
transform 1 0 28612 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_305
timestamp 1667941163
transform 1 0 29164 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1667941163
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1667941163
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1667941163
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1667941163
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1667941163
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_389
timestamp 1667941163
transform 1 0 36892 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_397
timestamp 1667941163
transform 1 0 37628 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_405
timestamp 1667941163
transform 1 0 38364 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_9
timestamp 1667941163
transform 1 0 1932 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_30
timestamp 1667941163
transform 1 0 3864 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_54
timestamp 1667941163
transform 1 0 6072 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_61
timestamp 1667941163
transform 1 0 6716 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_85
timestamp 1667941163
transform 1 0 8924 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_110
timestamp 1667941163
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_136
timestamp 1667941163
transform 1 0 13616 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_160
timestamp 1667941163
transform 1 0 15824 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_166
timestamp 1667941163
transform 1 0 16376 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_175
timestamp 1667941163
transform 1 0 17204 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_182
timestamp 1667941163
transform 1 0 17848 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_188
timestamp 1667941163
transform 1 0 18400 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_192
timestamp 1667941163
transform 1 0 18768 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_202
timestamp 1667941163
transform 1 0 19688 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_212
timestamp 1667941163
transform 1 0 20608 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_218
timestamp 1667941163
transform 1 0 21160 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 1667941163
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_230
timestamp 1667941163
transform 1 0 22264 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_237
timestamp 1667941163
transform 1 0 22908 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_244
timestamp 1667941163
transform 1 0 23552 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_251
timestamp 1667941163
transform 1 0 24196 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_257
timestamp 1667941163
transform 1 0 24748 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_263
timestamp 1667941163
transform 1 0 25300 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_272
timestamp 1667941163
transform 1 0 26128 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_278
timestamp 1667941163
transform 1 0 26680 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_288
timestamp 1667941163
transform 1 0 27600 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_294
timestamp 1667941163
transform 1 0 28152 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_300
timestamp 1667941163
transform 1 0 28704 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_306
timestamp 1667941163
transform 1 0 29256 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_312
timestamp 1667941163
transform 1 0 29808 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_324
timestamp 1667941163
transform 1 0 30912 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1667941163
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1667941163
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1667941163
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1667941163
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1667941163
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_397
timestamp 1667941163
transform 1 0 37628 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1667941163
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_26
timestamp 1667941163
transform 1 0 3496 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_33
timestamp 1667941163
transform 1 0 4140 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_54
timestamp 1667941163
transform 1 0 6072 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_61
timestamp 1667941163
transform 1 0 6716 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_82
timestamp 1667941163
transform 1 0 8648 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_89
timestamp 1667941163
transform 1 0 9292 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_110
timestamp 1667941163
transform 1 0 11224 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_135
timestamp 1667941163
transform 1 0 13524 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1667941163
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_163
timestamp 1667941163
transform 1 0 16100 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_167
timestamp 1667941163
transform 1 0 16468 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_175
timestamp 1667941163
transform 1 0 17204 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_182
timestamp 1667941163
transform 1 0 17848 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1667941163
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1667941163
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_203
timestamp 1667941163
transform 1 0 19780 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_209
timestamp 1667941163
transform 1 0 20332 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_216
timestamp 1667941163
transform 1 0 20976 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_222
timestamp 1667941163
transform 1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_231
timestamp 1667941163
transform 1 0 22356 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_238
timestamp 1667941163
transform 1 0 23000 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_244
timestamp 1667941163
transform 1 0 23552 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_250
timestamp 1667941163
transform 1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_259
timestamp 1667941163
transform 1 0 24932 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_267
timestamp 1667941163
transform 1 0 25668 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_275
timestamp 1667941163
transform 1 0 26404 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_278
timestamp 1667941163
transform 1 0 26680 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_287
timestamp 1667941163
transform 1 0 27508 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_293
timestamp 1667941163
transform 1 0 28060 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_299
timestamp 1667941163
transform 1 0 28612 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_305
timestamp 1667941163
transform 1 0 29164 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_315
timestamp 1667941163
transform 1 0 30084 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_322
timestamp 1667941163
transform 1 0 30728 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_328
timestamp 1667941163
transform 1 0 31280 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_343
timestamp 1667941163
transform 1 0 32660 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_351
timestamp 1667941163
transform 1 0 33396 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1667941163
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1667941163
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_370
timestamp 1667941163
transform 1 0 35144 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_384
timestamp 1667941163
transform 1 0 36432 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_390
timestamp 1667941163
transform 1 0 36984 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_393
timestamp 1667941163
transform 1 0 37260 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_399
timestamp 1667941163
transform 1 0 37812 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_405
timestamp 1667941163
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _213_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17848 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _214_
timestamp 1667941163
transform -1 0 15548 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _215_
timestamp 1667941163
transform 1 0 14260 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _216_
timestamp 1667941163
transform 1 0 13524 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _217_
timestamp 1667941163
transform 1 0 22724 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _218_
timestamp 1667941163
transform 1 0 17940 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _219_
timestamp 1667941163
transform 1 0 16008 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 1667941163
transform 1 0 14168 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _221_
timestamp 1667941163
transform 1 0 20700 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1667941163
transform 1 0 17020 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _223_
timestamp 1667941163
transform -1 0 17112 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _224_
timestamp 1667941163
transform -1 0 17020 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _225_
timestamp 1667941163
transform -1 0 17388 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _226_
timestamp 1667941163
transform 1 0 18308 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _227_
timestamp 1667941163
transform 1 0 19504 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1667941163
transform -1 0 20516 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _229_
timestamp 1667941163
transform 1 0 18584 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _230_
timestamp 1667941163
transform 1 0 17204 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _231_
timestamp 1667941163
transform 1 0 18308 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _232_
timestamp 1667941163
transform -1 0 21252 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _233_
timestamp 1667941163
transform 1 0 18584 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _234_
timestamp 1667941163
transform 1 0 10948 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1667941163
transform 1 0 11868 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _236_
timestamp 1667941163
transform -1 0 17664 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _237_
timestamp 1667941163
transform -1 0 15916 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _238_
timestamp 1667941163
transform -1 0 7452 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 1667941163
transform -1 0 13524 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 1667941163
transform -1 0 17480 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _241_
timestamp 1667941163
transform -1 0 13800 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _242_
timestamp 1667941163
transform 1 0 14260 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1667941163
transform 1 0 14444 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _244_
timestamp 1667941163
transform 1 0 16560 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _245_
timestamp 1667941163
transform -1 0 16560 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _246_
timestamp 1667941163
transform -1 0 20332 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _247_
timestamp 1667941163
transform -1 0 6808 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1667941163
transform -1 0 16376 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 1667941163
transform -1 0 12328 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _250_
timestamp 1667941163
transform 1 0 19412 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1667941163
transform 1 0 11408 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1667941163
transform 1 0 13432 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1667941163
transform 1 0 16836 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1667941163
transform 1 0 19412 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1667941163
transform 1 0 7728 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp 1667941163
transform -1 0 16192 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 1667941163
transform -1 0 15640 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 1667941163
transform -1 0 20976 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1667941163
transform -1 0 14904 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp 1667941163
transform 1 0 10304 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _261_
timestamp 1667941163
transform 1 0 10028 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp 1667941163
transform 1 0 7728 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _263_
timestamp 1667941163
transform -1 0 6072 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1667941163
transform 1 0 9568 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1667941163
transform -1 0 6808 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 1667941163
transform 1 0 6440 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _267_
timestamp 1667941163
transform 1 0 6900 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _268_
timestamp 1667941163
transform 1 0 8372 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _269_
timestamp 1667941163
transform 1 0 7820 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1667941163
transform 1 0 2576 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1667941163
transform 1 0 15456 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _272_
timestamp 1667941163
transform 1 0 10580 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1667941163
transform 1 0 8924 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _274_
timestamp 1667941163
transform -1 0 3404 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _275_
timestamp 1667941163
transform 1 0 8372 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _276_
timestamp 1667941163
transform 1 0 6072 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _277_
timestamp 1667941163
transform 1 0 8280 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _278_
timestamp 1667941163
transform 1 0 3220 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _279_
timestamp 1667941163
transform -1 0 4048 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1667941163
transform 1 0 4508 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _281_
timestamp 1667941163
transform -1 0 3496 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _282_
timestamp 1667941163
transform 1 0 9844 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _283_
timestamp 1667941163
transform 1 0 16100 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _284_
timestamp 1667941163
transform -1 0 20332 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _285_
timestamp 1667941163
transform 1 0 18032 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _286_
timestamp 1667941163
transform -1 0 2852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _287_
timestamp 1667941163
transform 1 0 16560 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _288_
timestamp 1667941163
transform -1 0 15640 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _289_
timestamp 1667941163
transform -1 0 2208 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _290_
timestamp 1667941163
transform 1 0 4600 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _291_
timestamp 1667941163
transform 1 0 7728 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _292_
timestamp 1667941163
transform -1 0 20332 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _293_
timestamp 1667941163
transform -1 0 20332 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _294_
timestamp 1667941163
transform -1 0 19688 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1667941163
transform -1 0 17112 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1667941163
transform 1 0 16100 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1667941163
transform 1 0 17940 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1667941163
transform -1 0 19044 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1667941163
transform -1 0 21252 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _300_
timestamp 1667941163
transform 1 0 18216 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _301_
timestamp 1667941163
transform 1 0 17572 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _302_
timestamp 1667941163
transform 1 0 17940 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _303_
timestamp 1667941163
transform -1 0 19320 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _304_
timestamp 1667941163
transform 1 0 17572 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _305_
timestamp 1667941163
transform 1 0 17112 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _306_
timestamp 1667941163
transform 1 0 5152 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _307_
timestamp 1667941163
transform 1 0 9568 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _308_
timestamp 1667941163
transform -1 0 12420 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _309_
timestamp 1667941163
transform -1 0 13156 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1667941163
transform 1 0 5796 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _311_
timestamp 1667941163
transform 1 0 10212 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _312_
timestamp 1667941163
transform -1 0 11224 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _313_
timestamp 1667941163
transform 1 0 11500 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _314_
timestamp 1667941163
transform 1 0 5888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _315_
timestamp 1667941163
transform 1 0 13432 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _316_
timestamp 1667941163
transform 1 0 13708 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _317_
timestamp 1667941163
transform 1 0 13064 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _318_
timestamp 1667941163
transform 1 0 3864 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _319_
timestamp 1667941163
transform 1 0 10304 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _320_
timestamp 1667941163
transform 1 0 7084 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _321_
timestamp 1667941163
transform 1 0 8372 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _322_
timestamp 1667941163
transform 1 0 4508 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _323_
timestamp 1667941163
transform 1 0 5796 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _324_
timestamp 1667941163
transform 1 0 7084 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _325_
timestamp 1667941163
transform 1 0 7084 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _326_
timestamp 1667941163
transform 1 0 4784 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _327_
timestamp 1667941163
transform 1 0 7176 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _328_
timestamp 1667941163
transform 1 0 8372 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _329_
timestamp 1667941163
transform 1 0 10948 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _330_
timestamp 1667941163
transform -1 0 17112 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _331_
timestamp 1667941163
transform -1 0 20332 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _332_
timestamp 1667941163
transform -1 0 20332 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _333_
timestamp 1667941163
transform 1 0 5152 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _334_
timestamp 1667941163
transform 1 0 9384 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _335_
timestamp 1667941163
transform 1 0 5796 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _336_
timestamp 1667941163
transform 1 0 6624 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _337_
timestamp 1667941163
transform 1 0 6808 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _338_
timestamp 1667941163
transform 1 0 9660 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp 1667941163
transform 1 0 5152 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _340_
timestamp 1667941163
transform 1 0 13064 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _341_
timestamp 1667941163
transform -1 0 16376 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _342_
timestamp 1667941163
transform 1 0 2576 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _343_
timestamp 1667941163
transform -1 0 14904 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _344_
timestamp 1667941163
transform 1 0 21252 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1667941163
transform 1 0 8832 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp 1667941163
transform -1 0 14720 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1667941163
transform 1 0 5796 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _348_
timestamp 1667941163
transform -1 0 15088 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _349_
timestamp 1667941163
transform 1 0 5796 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _350_
timestamp 1667941163
transform -1 0 16376 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _351_
timestamp 1667941163
transform -1 0 6900 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _352_
timestamp 1667941163
transform 1 0 3956 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _353_
timestamp 1667941163
transform -1 0 15088 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _354_
timestamp 1667941163
transform -1 0 13800 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _355_
timestamp 1667941163
transform -1 0 13800 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _356_
timestamp 1667941163
transform -1 0 24840 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _357_
timestamp 1667941163
transform 1 0 6716 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _358_
timestamp 1667941163
transform -1 0 2576 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _359_
timestamp 1667941163
transform -1 0 11960 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _360_
timestamp 1667941163
transform -1 0 19964 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _361_
timestamp 1667941163
transform -1 0 15732 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _362_
timestamp 1667941163
transform -1 0 29532 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _363_
timestamp 1667941163
transform 1 0 8372 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _364_
timestamp 1667941163
transform 1 0 10856 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp 1667941163
transform 1 0 29716 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _366_
timestamp 1667941163
transform -1 0 19688 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _367_
timestamp 1667941163
transform -1 0 21344 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _368_
timestamp 1667941163
transform -1 0 25576 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _369_
timestamp 1667941163
transform -1 0 18400 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _370_
timestamp 1667941163
transform -1 0 20976 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _371_
timestamp 1667941163
transform 1 0 5244 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _372_
timestamp 1667941163
transform -1 0 7176 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _373_
timestamp 1667941163
transform -1 0 17848 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _374_
timestamp 1667941163
transform -1 0 10580 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _375_
timestamp 1667941163
transform 1 0 17848 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _376_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 4784 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _377_
timestamp 1667941163
transform 1 0 10764 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _378_
timestamp 1667941163
transform 1 0 16100 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _379_
timestamp 1667941163
transform 1 0 28336 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _380_
timestamp 1667941163
transform -1 0 14444 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _381_
timestamp 1667941163
transform 1 0 13524 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _382_
timestamp 1667941163
transform -1 0 30636 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _383_
timestamp 1667941163
transform -1 0 18860 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _384_
timestamp 1667941163
transform 1 0 18952 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _385_
timestamp 1667941163
transform 1 0 27324 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _386_
timestamp 1667941163
transform 1 0 23920 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _387_
timestamp 1667941163
transform -1 0 29992 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _388_
timestamp 1667941163
transform 1 0 8464 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _389_
timestamp 1667941163
transform -1 0 15732 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _390_
timestamp 1667941163
transform -1 0 29624 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _391_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 20608 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _392_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19872 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _393_
timestamp 1667941163
transform -1 0 2116 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _394_
timestamp 1667941163
transform -1 0 21068 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _395_
timestamp 1667941163
transform -1 0 4232 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _396_
timestamp 1667941163
transform 1 0 3956 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _397_
timestamp 1667941163
transform 1 0 7820 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _398_
timestamp 1667941163
transform -1 0 19688 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _399_
timestamp 1667941163
transform 1 0 2484 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _400_
timestamp 1667941163
transform 1 0 2484 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _401_
timestamp 1667941163
transform -1 0 2576 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _402_
timestamp 1667941163
transform 1 0 4232 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _403_
timestamp 1667941163
transform 1 0 20792 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _404_
timestamp 1667941163
transform 1 0 3956 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _405_
timestamp 1667941163
transform 1 0 3956 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _406_
timestamp 1667941163
transform 1 0 2944 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _407_
timestamp 1667941163
transform 1 0 1840 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _408_
timestamp 1667941163
transform 1 0 1840 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _409_
timestamp 1667941163
transform -1 0 8648 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _410_
timestamp 1667941163
transform 1 0 9108 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _411_
timestamp 1667941163
transform -1 0 10580 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _412_
timestamp 1667941163
transform -1 0 11224 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _413_
timestamp 1667941163
transform 1 0 3956 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _414_
timestamp 1667941163
transform 1 0 19964 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _415_
timestamp 1667941163
transform -1 0 9384 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _416_
timestamp 1667941163
transform 1 0 6716 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _417_
timestamp 1667941163
transform 1 0 5796 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _418_
timestamp 1667941163
transform -1 0 4324 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _419_
timestamp 1667941163
transform 1 0 2484 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _420_
timestamp 1667941163
transform 1 0 1840 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _421_
timestamp 1667941163
transform 1 0 3128 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _422_
timestamp 1667941163
transform 1 0 4692 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _423_
timestamp 1667941163
transform -1 0 7820 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _424_
timestamp 1667941163
transform -1 0 9936 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _425_
timestamp 1667941163
transform 1 0 19872 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _426_
timestamp 1667941163
transform 1 0 2300 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _427_
timestamp 1667941163
transform 1 0 1840 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _428_
timestamp 1667941163
transform 1 0 1840 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _429_
timestamp 1667941163
transform 1 0 3128 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _430_
timestamp 1667941163
transform 1 0 3220 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _431_
timestamp 1667941163
transform 1 0 2484 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _432_
timestamp 1667941163
transform -1 0 3864 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _433_
timestamp 1667941163
transform -1 0 22264 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _434_
timestamp 1667941163
transform 1 0 2944 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _435_
timestamp 1667941163
transform 1 0 6532 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _436_
timestamp 1667941163
transform -1 0 19688 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _437_
timestamp 1667941163
transform -1 0 19688 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _438_
timestamp 1667941163
transform -1 0 19688 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _439_
timestamp 1667941163
transform -1 0 18952 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _440_
timestamp 1667941163
transform -1 0 19688 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _441_
timestamp 1667941163
transform -1 0 18768 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _442_
timestamp 1667941163
transform -1 0 20424 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _443_
timestamp 1667941163
transform 1 0 20792 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _444_
timestamp 1667941163
transform -1 0 18400 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _445_
timestamp 1667941163
transform -1 0 19044 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _446_
timestamp 1667941163
transform -1 0 19044 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _447_
timestamp 1667941163
transform 1 0 20056 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _448_
timestamp 1667941163
transform -1 0 20700 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _449_
timestamp 1667941163
transform -1 0 22264 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _450_
timestamp 1667941163
transform -1 0 21896 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _451_
timestamp 1667941163
transform -1 0 22264 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _452_
timestamp 1667941163
transform -1 0 21528 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _453_
timestamp 1667941163
transform -1 0 21712 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _454_
timestamp 1667941163
transform 1 0 22632 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _455_
timestamp 1667941163
transform -1 0 22540 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _456_
timestamp 1667941163
transform -1 0 21896 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _457_
timestamp 1667941163
transform -1 0 21344 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _458_
timestamp 1667941163
transform -1 0 20424 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _459_
timestamp 1667941163
transform -1 0 19780 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _460_
timestamp 1667941163
transform -1 0 18952 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _461_
timestamp 1667941163
transform -1 0 18952 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _462_
timestamp 1667941163
transform -1 0 19780 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _463_
timestamp 1667941163
transform -1 0 19688 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _464_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 3864 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _465_
timestamp 1667941163
transform 1 0 14260 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _466_
timestamp 1667941163
transform 1 0 1656 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _467_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 6992 0 1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _468_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6992 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _469_
timestamp 1667941163
transform -1 0 9292 0 -1 34816
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _470_
timestamp 1667941163
transform 1 0 1656 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _471_
timestamp 1667941163
transform 1 0 1656 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _472_
timestamp 1667941163
transform -1 0 3496 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _473_
timestamp 1667941163
transform -1 0 7452 0 1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _474_
timestamp 1667941163
transform -1 0 5612 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _475_
timestamp 1667941163
transform -1 0 7452 0 1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _476_
timestamp 1667941163
transform -1 0 5060 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _477_
timestamp 1667941163
transform -1 0 3496 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _478_
timestamp 1667941163
transform -1 0 5704 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _479_
timestamp 1667941163
transform -1 0 9476 0 -1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _480_
timestamp 1667941163
transform -1 0 11224 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _481_
timestamp 1667941163
transform -1 0 9660 0 -1 35904
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _482_
timestamp 1667941163
transform 1 0 4600 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _483_
timestamp 1667941163
transform -1 0 6072 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _484_
timestamp 1667941163
transform 1 0 4600 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _485_
timestamp 1667941163
transform -1 0 13616 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _486_
timestamp 1667941163
transform 1 0 6992 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _487_
timestamp 1667941163
transform 1 0 2944 0 -1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _488_
timestamp 1667941163
transform 1 0 2024 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _489_
timestamp 1667941163
transform -1 0 3496 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _490_
timestamp 1667941163
transform -1 0 5796 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _491_
timestamp 1667941163
transform -1 0 8556 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _492_
timestamp 1667941163
transform -1 0 8832 0 -1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _493_
timestamp 1667941163
transform 1 0 6808 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _494_
timestamp 1667941163
transform 1 0 1656 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _495_
timestamp 1667941163
transform -1 0 16100 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _496_
timestamp 1667941163
transform -1 0 3496 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _497_
timestamp 1667941163
transform -1 0 5520 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _498_
timestamp 1667941163
transform -1 0 5612 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _499_
timestamp 1667941163
transform 1 0 3956 0 1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _500_
timestamp 1667941163
transform 1 0 1656 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _501_
timestamp 1667941163
transform -1 0 6072 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _502_
timestamp 1667941163
transform -1 0 15732 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _503_
timestamp 1667941163
transform -1 0 8648 0 1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _504_
timestamp 1667941163
transform -1 0 15916 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _505_
timestamp 1667941163
transform 1 0 9292 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _506_
timestamp 1667941163
transform -1 0 13524 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _507_
timestamp 1667941163
transform 1 0 13984 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _508_
timestamp 1667941163
transform 1 0 4232 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _509_
timestamp 1667941163
transform -1 0 12604 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _510_
timestamp 1667941163
transform 1 0 10580 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _511_
timestamp 1667941163
transform 1 0 10672 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _512_
timestamp 1667941163
transform -1 0 13524 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _513_
timestamp 1667941163
transform 1 0 11684 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _514_
timestamp 1667941163
transform 1 0 9108 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _515_
timestamp 1667941163
transform 1 0 11224 0 1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _516_
timestamp 1667941163
transform -1 0 12236 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _517_
timestamp 1667941163
transform 1 0 9292 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _518_
timestamp 1667941163
transform 1 0 11684 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _519_
timestamp 1667941163
transform 1 0 9384 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _520_
timestamp 1667941163
transform 1 0 6808 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _521_
timestamp 1667941163
transform -1 0 13064 0 1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _522_
timestamp 1667941163
transform -1 0 13616 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _523_
timestamp 1667941163
transform 1 0 11684 0 -1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _524_
timestamp 1667941163
transform 1 0 11316 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _525_
timestamp 1667941163
transform 1 0 6808 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _526_
timestamp 1667941163
transform -1 0 8648 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _527_
timestamp 1667941163
transform -1 0 13524 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _528_
timestamp 1667941163
transform 1 0 11684 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _529_
timestamp 1667941163
transform 1 0 9384 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _541_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 38088 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _542_
timestamp 1667941163
transform -1 0 29256 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _543_
timestamp 1667941163
transform -1 0 18952 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _544_
timestamp 1667941163
transform 1 0 37812 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _545_
timestamp 1667941163
transform -1 0 14996 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _546_
timestamp 1667941163
transform -1 0 26128 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _547_
timestamp 1667941163
transform -1 0 17848 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _548_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 15824 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _549_
timestamp 1667941163
transform 1 0 1748 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _550_
timestamp 1667941163
transform 1 0 6440 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _551_
timestamp 1667941163
transform 1 0 33948 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _552_
timestamp 1667941163
transform 1 0 13524 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _553_
timestamp 1667941163
transform 1 0 8464 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _554_
timestamp 1667941163
transform 1 0 4232 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _555_
timestamp 1667941163
transform 1 0 1748 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _556_
timestamp 1667941163
transform -1 0 11224 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _557_
timestamp 1667941163
transform -1 0 31188 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _558_
timestamp 1667941163
transform -1 0 19688 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _559_
timestamp 1667941163
transform 1 0 2300 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _560_
timestamp 1667941163
transform -1 0 38088 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _561_
timestamp 1667941163
transform -1 0 17204 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _562_
timestamp 1667941163
transform -1 0 24656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _563_
timestamp 1667941163
transform 1 0 27784 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _564_
timestamp 1667941163
transform 1 0 14260 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _565_
timestamp 1667941163
transform 1 0 14260 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _566_
timestamp 1667941163
transform 1 0 12144 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _567_
timestamp 1667941163
transform -1 0 23828 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _568_
timestamp 1667941163
transform -1 0 38088 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _569_
timestamp 1667941163
transform 1 0 17480 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _570_
timestamp 1667941163
transform -1 0 17480 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _571_
timestamp 1667941163
transform -1 0 31004 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _572_
timestamp 1667941163
transform -1 0 18860 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _573_
timestamp 1667941163
transform 1 0 13524 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _574_
timestamp 1667941163
transform -1 0 22632 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _575_
timestamp 1667941163
transform 1 0 12052 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _576_
timestamp 1667941163
transform -1 0 16376 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _577_
timestamp 1667941163
transform -1 0 2760 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _578_
timestamp 1667941163
transform 1 0 18216 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _579_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 15272 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _580_
timestamp 1667941163
transform 1 0 16836 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _581_
timestamp 1667941163
transform 1 0 9108 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _582_
timestamp 1667941163
transform 1 0 12880 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _583__91 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 5428 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _583_
timestamp 1667941163
transform 1 0 10212 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _584_
timestamp 1667941163
transform 1 0 9660 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _585_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 12420 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _586_
timestamp 1667941163
transform 1 0 14444 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _587_
timestamp 1667941163
transform 1 0 14812 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _588_
timestamp 1667941163
transform 1 0 9200 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _589_
timestamp 1667941163
transform 1 0 9292 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _590_
timestamp 1667941163
transform 1 0 16468 0 1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _591_
timestamp 1667941163
transform -1 0 9292 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _592_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 9016 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _592__92
timestamp 1667941163
transform -1 0 8004 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _593_
timestamp 1667941163
transform 1 0 9108 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _594_
timestamp 1667941163
transform 1 0 7820 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _595_
timestamp 1667941163
transform 1 0 12696 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _596_
timestamp 1667941163
transform 1 0 10396 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _597_
timestamp 1667941163
transform 1 0 12144 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _598_
timestamp 1667941163
transform -1 0 13248 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _599_
timestamp 1667941163
transform -1 0 8280 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _600_
timestamp 1667941163
transform 1 0 7360 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _601_
timestamp 1667941163
transform -1 0 13340 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _602_
timestamp 1667941163
transform -1 0 15088 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _603_
timestamp 1667941163
transform -1 0 10856 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _604_
timestamp 1667941163
transform -1 0 12512 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _605_
timestamp 1667941163
transform -1 0 12880 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _606__93
timestamp 1667941163
transform -1 0 9660 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _606_
timestamp 1667941163
transform 1 0 10488 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _607_
timestamp 1667941163
transform -1 0 15088 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _608_
timestamp 1667941163
transform -1 0 16284 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _609_
timestamp 1667941163
transform -1 0 12788 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _610_
timestamp 1667941163
transform 1 0 10672 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _611_
timestamp 1667941163
transform 1 0 11224 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _612_
timestamp 1667941163
transform 1 0 11684 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _613_
timestamp 1667941163
transform -1 0 16192 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _614_
timestamp 1667941163
transform -1 0 12420 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _615_
timestamp 1667941163
transform 1 0 18768 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _616_
timestamp 1667941163
transform -1 0 18952 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _617_
timestamp 1667941163
transform 1 0 17756 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _618__94
timestamp 1667941163
transform -1 0 19688 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _618_
timestamp 1667941163
transform 1 0 19964 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _619_
timestamp 1667941163
transform -1 0 20240 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _620_
timestamp 1667941163
transform 1 0 18216 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _621_
timestamp 1667941163
transform 1 0 17940 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _622_
timestamp 1667941163
transform 1 0 16836 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _623_
timestamp 1667941163
transform 1 0 18124 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _624_
timestamp 1667941163
transform 1 0 19872 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _625_
timestamp 1667941163
transform 1 0 18216 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _626_
timestamp 1667941163
transform 1 0 15548 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _627_
timestamp 1667941163
transform -1 0 11408 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _628_
timestamp 1667941163
transform 1 0 5428 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _629_
timestamp 1667941163
transform 1 0 3956 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _630__95
timestamp 1667941163
transform 1 0 16008 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _630_
timestamp 1667941163
transform -1 0 15916 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _631_
timestamp 1667941163
transform -1 0 16468 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _632_
timestamp 1667941163
transform -1 0 17112 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _633_
timestamp 1667941163
transform 1 0 18032 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _634_
timestamp 1667941163
transform -1 0 17664 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _635_
timestamp 1667941163
transform -1 0 11684 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _636_
timestamp 1667941163
transform -1 0 17664 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _637_
timestamp 1667941163
transform 1 0 10304 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _638_
timestamp 1667941163
transform 1 0 16836 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _639_
timestamp 1667941163
transform 1 0 7544 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _640_
timestamp 1667941163
transform 1 0 8004 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _641_
timestamp 1667941163
transform 1 0 9108 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _642_
timestamp 1667941163
transform 1 0 7268 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _642__96
timestamp 1667941163
transform -1 0 5704 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _643_
timestamp 1667941163
transform -1 0 10212 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _644_
timestamp 1667941163
transform 1 0 6900 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _645_
timestamp 1667941163
transform 1 0 10212 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _646_
timestamp 1667941163
transform 1 0 14812 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _647_
timestamp 1667941163
transform 1 0 7820 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _648_
timestamp 1667941163
transform 1 0 9200 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _649_
timestamp 1667941163
transform 1 0 9108 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _650_
timestamp 1667941163
transform -1 0 16284 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _651_
timestamp 1667941163
transform 1 0 11960 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _652_
timestamp 1667941163
transform 1 0 11684 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _653_
timestamp 1667941163
transform 1 0 9568 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _654_
timestamp 1667941163
transform 1 0 10396 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _654__97
timestamp 1667941163
transform -1 0 7452 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _655_
timestamp 1667941163
transform -1 0 14444 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _656_
timestamp 1667941163
transform 1 0 11684 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _657_
timestamp 1667941163
transform 1 0 10396 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _658_
timestamp 1667941163
transform 1 0 14904 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _659_
timestamp 1667941163
transform 1 0 15732 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _660_
timestamp 1667941163
transform 1 0 9016 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _661_
timestamp 1667941163
transform 1 0 10580 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _662_
timestamp 1667941163
transform -1 0 15180 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _663_
timestamp 1667941163
transform 1 0 16836 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _664_
timestamp 1667941163
transform -1 0 17756 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _665_
timestamp 1667941163
transform -1 0 18124 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _666__98
timestamp 1667941163
transform 1 0 16836 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _666_
timestamp 1667941163
transform -1 0 15916 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _667_
timestamp 1667941163
transform -1 0 15548 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _668_
timestamp 1667941163
transform -1 0 14812 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _669_
timestamp 1667941163
transform 1 0 14168 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _670_
timestamp 1667941163
transform 1 0 14260 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _671_
timestamp 1667941163
transform 1 0 16376 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _672_
timestamp 1667941163
transform 1 0 13984 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _673_
timestamp 1667941163
transform 1 0 11316 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _674_
timestamp 1667941163
transform 1 0 12972 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _675_
timestamp 1667941163
transform -1 0 15088 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _676_
timestamp 1667941163
transform 1 0 12788 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _677_
timestamp 1667941163
transform 1 0 12880 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _678_
timestamp 1667941163
transform -1 0 15088 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _678__99
timestamp 1667941163
transform -1 0 14812 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _679_
timestamp 1667941163
transform -1 0 15916 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _680_
timestamp 1667941163
transform -1 0 17572 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _681_
timestamp 1667941163
transform -1 0 15272 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _682_
timestamp 1667941163
transform -1 0 16468 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _683_
timestamp 1667941163
transform 1 0 13248 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _684_
timestamp 1667941163
transform 1 0 12604 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _685_
timestamp 1667941163
transform 1 0 15180 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _686_
timestamp 1667941163
transform 1 0 12236 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _687_
timestamp 1667941163
transform 1 0 17112 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _688_
timestamp 1667941163
transform 1 0 18308 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _689_
timestamp 1667941163
transform 1 0 18124 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _690__100
timestamp 1667941163
transform 1 0 20056 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _690_
timestamp 1667941163
transform 1 0 19872 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _691_
timestamp 1667941163
transform -1 0 20056 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _692_
timestamp 1667941163
transform -1 0 19688 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _693_
timestamp 1667941163
transform 1 0 16928 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _694_
timestamp 1667941163
transform 1 0 15916 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _695_
timestamp 1667941163
transform 1 0 17480 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _696_
timestamp 1667941163
transform 1 0 19780 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _697_
timestamp 1667941163
transform 1 0 18952 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _698_
timestamp 1667941163
transform 1 0 15548 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _699_
timestamp 1667941163
transform 1 0 18032 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _700__101
timestamp 1667941163
transform 1 0 23276 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _700_
timestamp 1667941163
transform -1 0 22908 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _701_
timestamp 1667941163
transform -1 0 16928 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _702_
timestamp 1667941163
transform -1 0 16376 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _703_
timestamp 1667941163
transform 1 0 13984 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _704_
timestamp 1667941163
transform 1 0 14076 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _705_
timestamp 1667941163
transform 1 0 18216 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _706_
timestamp 1667941163
transform 1 0 15180 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _707_
timestamp 1667941163
transform -1 0 15364 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1667941163
transform -1 0 38364 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1667941163
transform -1 0 38364 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 38364 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1667941163
transform -1 0 38364 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1667941163
transform 1 0 35512 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1667941163
transform 1 0 1564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1667941163
transform 1 0 1564 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1667941163
transform -1 0 32660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1667941163
transform -1 0 38364 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1667941163
transform 1 0 20700 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1667941163
transform -1 0 2944 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1667941163
transform -1 0 36984 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1667941163
transform 1 0 14904 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1667941163
transform 1 0 1564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1667941163
transform -1 0 38364 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1667941163
transform -1 0 14168 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1667941163
transform 1 0 1564 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1667941163
transform 1 0 2852 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1667941163
transform -1 0 38364 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1667941163
transform 1 0 9752 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1667941163
transform 1 0 1564 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1667941163
transform -1 0 38364 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp 1667941163
transform -1 0 38364 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1667941163
transform -1 0 4968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1667941163
transform 1 0 1564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1667941163
transform 1 0 1564 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1667941163
transform -1 0 28796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1667941163
transform 1 0 1564 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input29
timestamp 1667941163
transform 1 0 9108 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1667941163
transform -1 0 4232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1667941163
transform 1 0 11684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1667941163
transform -1 0 33948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1667941163
transform -1 0 38364 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1667941163
transform -1 0 38364 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input35
timestamp 1667941163
transform 1 0 1564 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input36
timestamp 1667941163
transform -1 0 2484 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input37 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 36248 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1667941163
transform 1 0 1564 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1667941163
transform -1 0 38364 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1667941163
transform 1 0 30452 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1667941163
transform 1 0 37996 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1667941163
transform 1 0 37996 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1667941163
transform -1 0 17204 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1667941163
transform 1 0 37996 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1667941163
transform -1 0 1932 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1667941163
transform 1 0 24564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1667941163
transform 1 0 37996 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1667941163
transform -1 0 2668 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1667941163
transform -1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1667941163
transform -1 0 1932 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1667941163
transform -1 0 8648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1667941163
transform 1 0 19412 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1667941163
transform -1 0 17204 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1667941163
transform 1 0 37996 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1667941163
transform 1 0 25300 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1667941163
transform 1 0 27140 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1667941163
transform 1 0 34868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1667941163
transform -1 0 1932 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1667941163
transform 1 0 37996 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1667941163
transform 1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1667941163
transform -1 0 1932 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1667941163
transform 1 0 29716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1667941163
transform 1 0 37996 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1667941163
transform -1 0 10764 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1667941163
transform 1 0 4600 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1667941163
transform 1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1667941163
transform -1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1667941163
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1667941163
transform -1 0 13340 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1667941163
transform 1 0 21988 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1667941163
transform -1 0 33948 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1667941163
transform -1 0 1932 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1667941163
transform -1 0 1932 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1667941163
transform -1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1667941163
transform 1 0 37444 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1667941163
transform 1 0 29716 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1667941163
transform 1 0 16836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1667941163
transform -1 0 37628 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1667941163
transform 1 0 37996 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1667941163
transform -1 0 1932 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1667941163
transform 1 0 37996 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1667941163
transform -1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1667941163
transform 1 0 12972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1667941163
transform 1 0 20056 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1667941163
transform 1 0 37996 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1667941163
transform 1 0 21988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1667941163
transform 1 0 32292 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1667941163
transform -1 0 7176 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1667941163
transform 1 0 27140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1667941163
transform -1 0 1932 0 -1 13056
box -38 -48 406 592
<< labels >>
flabel metal3 s 39200 26528 39800 26648 0 FreeSans 480 0 0 0 ccff_head
port 0 nsew signal input
flabel metal3 s 39200 37408 39800 37528 0 FreeSans 480 0 0 0 ccff_tail
port 1 nsew signal tristate
flabel metal2 s 38658 39200 38714 39800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 2 nsew signal input
flabel metal2 s 38014 200 38070 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 3 nsew signal input
flabel metal3 s 39200 19728 39800 19848 0 FreeSans 480 0 0 0 chany_bottom_in[11]
port 4 nsew signal input
flabel metal2 s 35438 39200 35494 39800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 5 nsew signal input
flabel metal3 s 200 3408 800 3528 0 FreeSans 480 0 0 0 chany_bottom_in[13]
port 6 nsew signal input
flabel metal3 s 200 19048 800 19168 0 FreeSans 480 0 0 0 chany_bottom_in[14]
port 7 nsew signal input
flabel metal2 s 31574 200 31630 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 8 nsew signal input
flabel metal3 s 39200 12248 39800 12368 0 FreeSans 480 0 0 0 chany_bottom_in[16]
port 9 nsew signal input
flabel metal2 s 20626 39200 20682 39800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 10 nsew signal input
flabel metal2 s 1950 39200 2006 39800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 11 nsew signal input
flabel metal2 s 36726 200 36782 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 12 nsew signal input
flabel metal2 s 14830 200 14886 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 13 nsew signal input
flabel metal3 s 200 4768 800 4888 0 FreeSans 480 0 0 0 chany_bottom_in[3]
port 14 nsew signal input
flabel metal3 s 39200 33328 39800 33448 0 FreeSans 480 0 0 0 chany_bottom_in[4]
port 15 nsew signal input
flabel metal2 s 13542 39200 13598 39800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 16 nsew signal input
flabel metal3 s 200 38768 800 38888 0 FreeSans 480 0 0 0 chany_bottom_in[6]
port 17 nsew signal input
flabel metal3 s 200 33328 800 33448 0 FreeSans 480 0 0 0 chany_bottom_in[7]
port 18 nsew signal input
flabel metal3 s 39200 5448 39800 5568 0 FreeSans 480 0 0 0 chany_bottom_in[8]
port 19 nsew signal input
flabel metal2 s 9678 200 9734 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 20 nsew signal input
flabel metal3 s 39200 28568 39800 28688 0 FreeSans 480 0 0 0 chany_bottom_out[0]
port 21 nsew signal tristate
flabel metal2 s 16762 39200 16818 39800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 22 nsew signal tristate
flabel metal3 s 39200 31968 39800 32088 0 FreeSans 480 0 0 0 chany_bottom_out[11]
port 23 nsew signal tristate
flabel metal3 s 200 27888 800 28008 0 FreeSans 480 0 0 0 chany_bottom_out[12]
port 24 nsew signal tristate
flabel metal2 s 23846 39200 23902 39800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 25 nsew signal tristate
flabel metal3 s 39200 29928 39800 30048 0 FreeSans 480 0 0 0 chany_bottom_out[14]
port 26 nsew signal tristate
flabel metal2 s 18 39200 74 39800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 27 nsew signal tristate
flabel metal3 s 200 1368 800 1488 0 FreeSans 480 0 0 0 chany_bottom_out[16]
port 28 nsew signal tristate
flabel metal3 s 200 15648 800 15768 0 FreeSans 480 0 0 0 chany_bottom_out[17]
port 29 nsew signal tristate
flabel metal2 s 8390 200 8446 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 30 nsew signal tristate
flabel metal2 s 18694 39200 18750 39800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 31 nsew signal tristate
flabel metal2 s 15474 39200 15530 39800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 32 nsew signal tristate
flabel metal3 s 39200 8848 39800 8968 0 FreeSans 480 0 0 0 chany_bottom_out[3]
port 33 nsew signal tristate
flabel metal2 s 25134 39200 25190 39800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 34 nsew signal tristate
flabel metal2 s 27066 39200 27122 39800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 35 nsew signal tristate
flabel metal2 s 34794 200 34850 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 36 nsew signal tristate
flabel metal3 s 200 17688 800 17808 0 FreeSans 480 0 0 0 chany_bottom_out[7]
port 37 nsew signal tristate
flabel metal3 s 39200 35368 39800 35488 0 FreeSans 480 0 0 0 chany_bottom_out[8]
port 38 nsew signal tristate
flabel metal2 s 25134 200 25190 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 39 nsew signal tristate
flabel metal3 s 200 21088 800 21208 0 FreeSans 480 0 0 0 chany_top_in[0]
port 40 nsew signal input
flabel metal3 s 39200 2048 39800 2168 0 FreeSans 480 0 0 0 chany_top_in[10]
port 41 nsew signal input
flabel metal3 s 39200 15648 39800 15768 0 FreeSans 480 0 0 0 chany_top_in[11]
port 42 nsew signal input
flabel metal2 s 4526 200 4582 800 0 FreeSans 224 90 0 0 chany_top_in[12]
port 43 nsew signal input
flabel metal3 s 200 13608 800 13728 0 FreeSans 480 0 0 0 chany_top_in[13]
port 44 nsew signal input
flabel metal3 s 200 31288 800 31408 0 FreeSans 480 0 0 0 chany_top_in[14]
port 45 nsew signal input
flabel metal2 s 28354 200 28410 800 0 FreeSans 224 90 0 0 chany_top_in[15]
port 46 nsew signal input
flabel metal3 s 200 29928 800 30048 0 FreeSans 480 0 0 0 chany_top_in[16]
port 47 nsew signal input
flabel metal2 s 7102 39200 7158 39800 0 FreeSans 224 90 0 0 chany_top_in[17]
port 48 nsew signal input
flabel metal2 s 3238 200 3294 800 0 FreeSans 224 90 0 0 chany_top_in[18]
port 49 nsew signal input
flabel metal2 s 11610 200 11666 800 0 FreeSans 224 90 0 0 chany_top_in[1]
port 50 nsew signal input
flabel metal2 s 33506 200 33562 800 0 FreeSans 224 90 0 0 chany_top_in[2]
port 51 nsew signal input
flabel metal3 s 39200 14288 39800 14408 0 FreeSans 480 0 0 0 chany_top_in[3]
port 52 nsew signal input
flabel metal3 s 39200 6808 39800 6928 0 FreeSans 480 0 0 0 chany_top_in[4]
port 53 nsew signal input
flabel metal3 s 200 6808 800 6928 0 FreeSans 480 0 0 0 chany_top_in[5]
port 54 nsew signal input
flabel metal3 s 200 36728 800 36848 0 FreeSans 480 0 0 0 chany_top_in[6]
port 55 nsew signal input
flabel metal3 s 39200 8 39800 128 0 FreeSans 480 0 0 0 chany_top_in[7]
port 56 nsew signal input
flabel metal3 s 200 8848 800 8968 0 FreeSans 480 0 0 0 chany_top_in[8]
port 57 nsew signal input
flabel metal3 s 39200 10888 39800 11008 0 FreeSans 480 0 0 0 chany_top_in[9]
port 58 nsew signal input
flabel metal3 s 200 24488 800 24608 0 FreeSans 480 0 0 0 chany_top_out[0]
port 59 nsew signal tristate
flabel metal2 s 29642 200 29698 800 0 FreeSans 224 90 0 0 chany_top_out[10]
port 60 nsew signal tristate
flabel metal3 s 39200 24488 39800 24608 0 FreeSans 480 0 0 0 chany_top_out[11]
port 61 nsew signal tristate
flabel metal2 s 10322 39200 10378 39800 0 FreeSans 224 90 0 0 chany_top_out[12]
port 62 nsew signal tristate
flabel metal2 s 5170 39200 5226 39800 0 FreeSans 224 90 0 0 chany_top_out[13]
port 63 nsew signal tristate
flabel metal2 s 18050 200 18106 800 0 FreeSans 224 90 0 0 chany_top_out[14]
port 64 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 chany_top_out[15]
port 65 nsew signal tristate
flabel metal2 s 23202 200 23258 800 0 FreeSans 224 90 0 0 chany_top_out[16]
port 66 nsew signal tristate
flabel metal2 s 12254 39200 12310 39800 0 FreeSans 224 90 0 0 chany_top_out[17]
port 67 nsew signal tristate
flabel metal2 s 21914 39200 21970 39800 0 FreeSans 224 90 0 0 chany_top_out[18]
port 68 nsew signal tristate
flabel metal2 s 33506 39200 33562 39800 0 FreeSans 224 90 0 0 chany_top_out[1]
port 69 nsew signal tristate
flabel metal3 s 200 26528 800 26648 0 FreeSans 480 0 0 0 chany_top_out[2]
port 70 nsew signal tristate
flabel metal3 s 200 22448 800 22568 0 FreeSans 480 0 0 0 chany_top_out[3]
port 71 nsew signal tristate
flabel metal2 s 1306 200 1362 800 0 FreeSans 224 90 0 0 chany_top_out[4]
port 72 nsew signal tristate
flabel metal2 s 37370 39200 37426 39800 0 FreeSans 224 90 0 0 chany_top_out[5]
port 73 nsew signal tristate
flabel metal2 s 28998 39200 29054 39800 0 FreeSans 224 90 0 0 chany_top_out[6]
port 74 nsew signal tristate
flabel metal2 s 16762 200 16818 800 0 FreeSans 224 90 0 0 chany_top_out[7]
port 75 nsew signal tristate
flabel metal3 s 39200 38768 39800 38888 0 FreeSans 480 0 0 0 chany_top_out[8]
port 76 nsew signal tristate
flabel metal3 s 39200 3408 39800 3528 0 FreeSans 480 0 0 0 chany_top_out[9]
port 77 nsew signal tristate
flabel metal3 s 200 10208 800 10328 0 FreeSans 480 0 0 0 left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
port 78 nsew signal tristate
flabel metal3 s 39200 21088 39800 21208 0 FreeSans 480 0 0 0 left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_
port 79 nsew signal tristate
flabel metal2 s 6458 200 6514 800 0 FreeSans 224 90 0 0 left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_
port 80 nsew signal tristate
flabel metal2 s 12898 200 12954 800 0 FreeSans 224 90 0 0 left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_
port 81 nsew signal tristate
flabel metal2 s 19982 200 20038 800 0 FreeSans 224 90 0 0 left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_
port 82 nsew signal tristate
flabel metal3 s 39200 23128 39800 23248 0 FreeSans 480 0 0 0 left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_
port 83 nsew signal tristate
flabel metal2 s 21270 200 21326 800 0 FreeSans 224 90 0 0 left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_
port 84 nsew signal tristate
flabel metal2 s 32218 39200 32274 39800 0 FreeSans 224 90 0 0 left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_
port 85 nsew signal tristate
flabel metal2 s 30286 39200 30342 39800 0 FreeSans 224 90 0 0 pReset
port 86 nsew signal input
flabel metal2 s 3882 39200 3938 39800 0 FreeSans 224 90 0 0 prog_clk
port 87 nsew signal input
flabel metal2 s 8390 39200 8446 39800 0 FreeSans 224 90 0 0 right_grid_left_width_0_height_0_subtile_0__pin_I_11_
port 88 nsew signal tristate
flabel metal2 s 26422 200 26478 800 0 FreeSans 224 90 0 0 right_grid_left_width_0_height_0_subtile_0__pin_I_3_
port 89 nsew signal tristate
flabel metal3 s 200 12248 800 12368 0 FreeSans 480 0 0 0 right_grid_left_width_0_height_0_subtile_0__pin_I_7_
port 90 nsew signal tristate
flabel metal3 s 200 35368 800 35488 0 FreeSans 480 0 0 0 vccd1
port 91 nsew signal bidirectional
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 91 nsew signal bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 91 nsew signal bidirectional
flabel metal3 s 39200 17688 39800 17808 0 FreeSans 480 0 0 0 vssd1
port 92 nsew signal bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 92 nsew signal bidirectional
rlabel metal1 19964 37536 19964 37536 0 vccd1
rlabel metal1 19964 36992 19964 36992 0 vssd1
rlabel metal1 1472 23834 1472 23834 0 _000_
rlabel metal1 16107 37230 16107 37230 0 _001_
rlabel metal1 4048 25466 4048 25466 0 _002_
rlabel metal1 4876 33830 4876 33830 0 _003_
rlabel metal2 7958 33694 7958 33694 0 _004_
rlabel metal1 19504 33626 19504 33626 0 _005_
rlabel metal1 1932 25466 1932 25466 0 _006_
rlabel metal1 2668 24378 2668 24378 0 _007_
rlabel metal1 2484 27098 2484 27098 0 _008_
rlabel metal2 6026 32266 6026 32266 0 _009_
rlabel via3 4669 34612 4669 34612 0 _010_
rlabel metal1 4876 34918 4876 34918 0 _011_
rlabel metal2 3082 28152 3082 28152 0 _012_
rlabel metal1 2070 26554 2070 26554 0 _013_
rlabel metal1 4186 25432 4186 25432 0 _014_
rlabel metal2 8510 32062 8510 32062 0 _015_
rlabel metal1 9469 30294 9469 30294 0 _016_
rlabel metal1 9660 34714 9660 34714 0 _017_
rlabel metal1 10902 34714 10902 34714 0 _018_
rlabel metal1 4370 36346 4370 36346 0 _019_
rlabel metal1 8786 34170 8786 34170 0 _020_
rlabel metal1 8257 31110 8257 31110 0 _021_
rlabel metal2 8326 30872 8326 30872 0 _022_
rlabel metal1 4232 31654 4232 31654 0 _023_
rlabel metal1 1978 26486 1978 26486 0 _024_
rlabel metal1 2024 26010 2024 26010 0 _025_
rlabel metal1 4002 25942 4002 25942 0 _026_
rlabel metal1 5980 31994 5980 31994 0 _027_
rlabel metal2 7774 32606 7774 32606 0 _028_
rlabel metal1 9752 34646 9752 34646 0 _029_
rlabel metal1 2116 24582 2116 24582 0 _030_
rlabel metal2 1978 24531 1978 24531 0 _031_
rlabel metal1 2024 27574 2024 27574 0 _032_
rlabel metal1 3765 32470 3765 32470 0 _033_
rlabel metal1 4094 26282 4094 26282 0 _034_
rlabel metal2 5198 28186 5198 28186 0 _035_
rlabel metal2 2990 36023 2990 36023 0 _036_
rlabel metal2 17342 35564 17342 35564 0 _037_
rlabel metal2 14950 35649 14950 35649 0 _038_
rlabel metal1 6808 34510 6808 34510 0 _039_
rlabel metal1 17572 31994 17572 31994 0 _040_
rlabel metal1 19412 33082 19412 33082 0 _041_
rlabel metal1 17894 36210 17894 36210 0 _042_
rlabel metal1 18308 36278 18308 36278 0 _043_
rlabel via2 13754 36363 13754 36363 0 _044_
rlabel metal1 17112 31178 17112 31178 0 _045_
rlabel metal2 20930 31552 20930 31552 0 _046_
rlabel metal1 16974 34714 16974 34714 0 _047_
rlabel metal1 17986 33422 17986 33422 0 _048_
rlabel metal1 17572 34510 17572 34510 0 _049_
rlabel metal1 11277 36074 11277 36074 0 _050_
rlabel metal1 22172 32538 22172 32538 0 _051_
rlabel metal2 21758 33626 21758 33626 0 _052_
rlabel via2 20746 36805 20746 36805 0 _053_
rlabel metal1 20976 36754 20976 36754 0 _054_
rlabel metal2 10718 37315 10718 37315 0 _055_
rlabel metal2 8234 37332 8234 37332 0 _056_
rlabel metal2 21850 30464 21850 30464 0 _057_
rlabel metal1 20700 30838 20700 30838 0 _058_
rlabel metal1 19596 31858 19596 31858 0 _059_
rlabel metal2 20286 34901 20286 34901 0 _060_
rlabel metal1 19550 35734 19550 35734 0 _061_
rlabel metal2 7866 35122 7866 35122 0 _062_
rlabel metal3 15778 30396 15778 30396 0 _063_
rlabel metal1 19550 31110 19550 31110 0 _064_
rlabel metal2 17986 32453 17986 32453 0 _065_
rlabel metal1 19113 35054 19113 35054 0 _066_
rlabel metal1 2668 23494 2668 23494 0 _067_
rlabel metal1 1886 25296 1886 25296 0 _068_
rlabel metal1 4830 20502 4830 20502 0 _069_
rlabel metal1 2944 21862 2944 21862 0 _070_
rlabel metal1 19504 32878 19504 32878 0 _071_
rlabel metal1 22356 30702 22356 30702 0 _072_
rlabel metal1 15686 33898 15686 33898 0 _073_
rlabel metal1 13478 33830 13478 33830 0 _074_
rlabel metal1 5750 26758 5750 26758 0 _075_
rlabel metal2 13110 30056 13110 30056 0 _076_
rlabel metal1 10120 27030 10120 27030 0 _077_
rlabel metal1 9883 25976 9883 25976 0 _078_
rlabel metal2 12650 28526 12650 28526 0 _079_
rlabel metal1 14720 29546 14720 29546 0 _080_
rlabel metal1 20148 31790 20148 31790 0 _081_
rlabel metal1 8648 28118 8648 28118 0 _082_
rlabel metal2 9522 28866 9522 28866 0 _083_
rlabel metal1 16698 32776 16698 32776 0 _084_
rlabel metal1 6992 25398 6992 25398 0 _085_
rlabel metal1 9246 23732 9246 23732 0 _086_
rlabel via2 7222 23579 7222 23579 0 _087_
rlabel metal2 8050 26588 8050 26588 0 _088_
rlabel metal1 9614 27642 9614 27642 0 _089_
rlabel metal2 9706 27710 9706 27710 0 _090_
rlabel metal1 12144 24854 12144 24854 0 _091_
rlabel metal1 8510 24208 8510 24208 0 _092_
rlabel metal1 7958 27030 7958 27030 0 _093_
rlabel metal1 5980 24786 5980 24786 0 _094_
rlabel metal2 13110 26214 13110 26214 0 _095_
rlabel metal1 14858 28424 14858 28424 0 _096_
rlabel metal2 10626 21760 10626 21760 0 _097_
rlabel metal1 9292 20502 9292 20502 0 _098_
rlabel metal2 11638 21284 11638 21284 0 _099_
rlabel metal2 11086 21012 11086 21012 0 _100_
rlabel metal1 14030 20570 14030 20570 0 _101_
rlabel metal1 14950 20502 14950 20502 0 _102_
rlabel metal1 12788 20026 12788 20026 0 _103_
rlabel metal1 11592 20026 11592 20026 0 _104_
rlabel metal1 9246 22066 9246 22066 0 _105_
rlabel metal1 11362 22542 11362 22542 0 _106_
rlabel metal1 15962 19720 15962 19720 0 _107_
rlabel metal1 10396 23290 10396 23290 0 _108_
rlabel metal1 18354 33286 18354 33286 0 _109_
rlabel metal2 18722 29240 18722 29240 0 _110_
rlabel metal2 17986 26078 17986 26078 0 _111_
rlabel metal1 18860 27030 18860 27030 0 _112_
rlabel metal1 17802 26010 17802 26010 0 _113_
rlabel metal1 18078 27506 18078 27506 0 _114_
rlabel metal2 18170 24174 18170 24174 0 _115_
rlabel metal1 16330 28186 16330 28186 0 _116_
rlabel metal1 18676 29206 18676 29206 0 _117_
rlabel metal2 21114 25636 21114 25636 0 _118_
rlabel metal1 18814 26010 18814 26010 0 _119_
rlabel metal1 15824 24854 15824 24854 0 _120_
rlabel metal1 6670 26418 6670 26418 0 _121_
rlabel metal1 3680 27574 3680 27574 0 _122_
rlabel metal1 3542 28492 3542 28492 0 _123_
rlabel metal1 15594 34510 15594 34510 0 _124_
rlabel metal2 16238 28696 16238 28696 0 _125_
rlabel metal2 16928 31790 16928 31790 0 _126_
rlabel metal2 18262 29784 18262 29784 0 _127_
rlabel metal1 17618 32504 17618 32504 0 _128_
rlabel metal1 10718 32810 10718 32810 0 _129_
rlabel metal2 17434 35326 17434 35326 0 _130_
rlabel metal1 10534 23800 10534 23800 0 _131_
rlabel metal1 16422 27098 16422 27098 0 _132_
rlabel metal1 4324 27506 4324 27506 0 _133_
rlabel metal1 4508 27982 4508 27982 0 _134_
rlabel metal1 8878 22678 8878 22678 0 _135_
rlabel metal2 6210 25704 6210 25704 0 _136_
rlabel metal2 9982 26877 9982 26877 0 _137_
rlabel metal1 5382 27370 5382 27370 0 _138_
rlabel metal1 9752 22746 9752 22746 0 _139_
rlabel metal1 14858 31416 14858 31416 0 _140_
rlabel metal1 5382 29240 5382 29240 0 _141_
rlabel metal1 8924 31790 8924 31790 0 _142_
rlabel metal2 9338 27489 9338 27489 0 _143_
rlabel metal2 16054 34238 16054 34238 0 _144_
rlabel metal1 11822 27370 11822 27370 0 _145_
rlabel metal2 11914 27166 11914 27166 0 _146_
rlabel metal1 8188 24582 8188 24582 0 _147_
rlabel metal1 10166 22678 10166 22678 0 _148_
rlabel metal2 14214 25364 14214 25364 0 _149_
rlabel metal1 8832 23698 8832 23698 0 _150_
rlabel metal1 10396 29206 10396 29206 0 _151_
rlabel metal1 14398 30634 14398 30634 0 _152_
rlabel metal1 16330 27370 16330 27370 0 _153_
rlabel metal2 9246 27081 9246 27081 0 _154_
rlabel metal2 10810 27166 10810 27166 0 _155_
rlabel metal2 14950 32096 14950 32096 0 _156_
rlabel metal1 17526 27030 17526 27030 0 _157_
rlabel metal2 17526 29342 17526 29342 0 _158_
rlabel metal1 17434 33286 17434 33286 0 _159_
rlabel metal1 14628 23766 14628 23766 0 _160_
rlabel metal1 15364 26418 15364 26418 0 _161_
rlabel metal2 14582 25534 14582 25534 0 _162_
rlabel metal2 14398 27438 14398 27438 0 _163_
rlabel metal2 14490 25466 14490 25466 0 _164_
rlabel metal1 17296 29546 17296 29546 0 _165_
rlabel metal1 14214 22712 14214 22712 0 _166_
rlabel metal1 8234 24378 8234 24378 0 _167_
rlabel metal1 12834 26316 12834 26316 0 _168_
rlabel metal1 14214 31858 14214 31858 0 _169_
rlabel metal1 10718 22576 10718 22576 0 _170_
rlabel metal1 13386 20026 13386 20026 0 _171_
rlabel metal2 15502 20706 15502 20706 0 _172_
rlabel metal2 15686 21692 15686 21692 0 _173_
rlabel metal2 16698 21284 16698 21284 0 _174_
rlabel metal1 15410 22066 15410 22066 0 _175_
rlabel metal2 17526 24854 17526 24854 0 _176_
rlabel metal2 11638 27438 11638 27438 0 _177_
rlabel metal1 13110 22066 13110 22066 0 _178_
rlabel metal2 15410 23052 15410 23052 0 _179_
rlabel metal2 12558 24956 12558 24956 0 _180_
rlabel metal2 17342 33218 17342 33218 0 _181_
rlabel metal1 18492 32742 18492 32742 0 _182_
rlabel metal1 18538 24378 18538 24378 0 _183_
rlabel metal2 20378 27234 20378 27234 0 _184_
rlabel metal1 19550 24854 19550 24854 0 _185_
rlabel metal1 20838 26010 20838 26010 0 _186_
rlabel metal2 17158 22814 17158 22814 0 _187_
rlabel metal1 16330 23018 16330 23018 0 _188_
rlabel metal1 17526 33830 17526 33830 0 _189_
rlabel metal1 19826 24378 19826 24378 0 _190_
rlabel metal1 18814 22678 18814 22678 0 _191_
rlabel metal1 16376 23834 16376 23834 0 _192_
rlabel metal2 18262 34680 18262 34680 0 _193_
rlabel metal2 22678 36584 22678 36584 0 _194_
rlabel metal2 20838 30226 20838 30226 0 _195_
rlabel metal1 15732 30294 15732 30294 0 _196_
rlabel metal2 14214 29886 14214 29886 0 _197_
rlabel metal2 14306 29342 14306 29342 0 _198_
rlabel metal1 18584 32470 18584 32470 0 _199_
rlabel metal2 15410 30158 15410 30158 0 _200_
rlabel via1 15134 27387 15134 27387 0 _201_
rlabel metal2 38226 26775 38226 26775 0 ccff_head
rlabel metal1 38272 36346 38272 36346 0 ccff_tail
rlabel metal1 38502 37434 38502 37434 0 chany_bottom_in[0]
rlabel metal1 38226 2414 38226 2414 0 chany_bottom_in[10]
rlabel via2 38318 19805 38318 19805 0 chany_bottom_in[11]
rlabel metal1 35512 37298 35512 37298 0 chany_bottom_in[12]
rlabel via2 1702 3485 1702 3485 0 chany_bottom_in[13]
rlabel metal2 1610 19023 1610 19023 0 chany_bottom_in[14]
rlabel metal2 31786 1989 31786 1989 0 chany_bottom_in[15]
rlabel metal2 38226 12563 38226 12563 0 chany_bottom_in[16]
rlabel metal1 20838 37230 20838 37230 0 chany_bottom_in[17]
rlabel metal2 1978 36866 1978 36866 0 chany_bottom_in[18]
rlabel metal1 36800 2346 36800 2346 0 chany_bottom_in[1]
rlabel metal1 14950 2346 14950 2346 0 chany_bottom_in[2]
rlabel via2 1610 4811 1610 4811 0 chany_bottom_in[3]
rlabel metal2 38226 33439 38226 33439 0 chany_bottom_in[4]
rlabel metal1 14306 34578 14306 34578 0 chany_bottom_in[5]
rlabel via2 2254 18955 2254 18955 0 chany_bottom_in[6]
rlabel metal3 1717 33388 1717 33388 0 chany_bottom_in[7]
rlabel metal2 38226 5559 38226 5559 0 chany_bottom_in[8]
rlabel metal1 9752 2414 9752 2414 0 chany_bottom_in[9]
rlabel metal2 38226 28815 38226 28815 0 chany_bottom_out[0]
rlabel metal1 16882 37094 16882 37094 0 chany_bottom_out[10]
rlabel metal2 38226 32113 38226 32113 0 chany_bottom_out[11]
rlabel metal3 1188 27948 1188 27948 0 chany_bottom_out[12]
rlabel metal2 24794 36992 24794 36992 0 chany_bottom_out[13]
rlabel via2 38226 30005 38226 30005 0 chany_bottom_out[14]
rlabel metal1 1196 37298 1196 37298 0 chany_bottom_out[15]
rlabel metal3 1188 1428 1188 1428 0 chany_bottom_out[16]
rlabel metal3 1188 15708 1188 15708 0 chany_bottom_out[17]
rlabel metal2 8418 1520 8418 1520 0 chany_bottom_out[18]
rlabel metal1 19182 37094 19182 37094 0 chany_bottom_out[1]
rlabel metal1 16376 36890 16376 36890 0 chany_bottom_out[2]
rlabel metal2 38226 8857 38226 8857 0 chany_bottom_out[3]
rlabel metal1 25346 37094 25346 37094 0 chany_bottom_out[4]
rlabel metal1 27232 37094 27232 37094 0 chany_bottom_out[5]
rlabel metal2 34822 1520 34822 1520 0 chany_bottom_out[6]
rlabel metal3 1188 17748 1188 17748 0 chany_bottom_out[7]
rlabel via2 38226 35445 38226 35445 0 chany_bottom_out[8]
rlabel metal2 25162 1520 25162 1520 0 chany_bottom_out[9]
rlabel via2 1610 21131 1610 21131 0 chany_top_in[0]
rlabel metal2 38226 2567 38226 2567 0 chany_top_in[10]
rlabel via2 38318 15691 38318 15691 0 chany_top_in[11]
rlabel metal1 4692 2346 4692 2346 0 chany_top_in[12]
rlabel metal2 1610 13583 1610 13583 0 chany_top_in[13]
rlabel metal2 2346 22749 2346 22749 0 chany_top_in[14]
rlabel metal1 28520 2346 28520 2346 0 chany_top_in[15]
rlabel metal2 1656 22372 1656 22372 0 chany_top_in[16]
rlabel metal2 9154 35105 9154 35105 0 chany_top_in[17]
rlabel metal1 3312 2278 3312 2278 0 chany_top_in[18]
rlabel metal1 11730 2346 11730 2346 0 chany_top_in[1]
rlabel metal1 33672 2346 33672 2346 0 chany_top_in[2]
rlabel via2 38318 14365 38318 14365 0 chany_top_in[3]
rlabel metal3 38740 6868 38740 6868 0 chany_top_in[4]
rlabel metal3 1142 6868 1142 6868 0 chany_top_in[5]
rlabel metal1 1978 19142 1978 19142 0 chany_top_in[6]
rlabel metal1 36708 2414 36708 2414 0 chany_top_in[7]
rlabel via2 1702 8891 1702 8891 0 chany_top_in[8]
rlabel metal2 38226 10999 38226 10999 0 chany_top_in[9]
rlabel metal3 1188 24548 1188 24548 0 chany_top_out[0]
rlabel metal2 29670 1520 29670 1520 0 chany_top_out[10]
rlabel via2 38226 24565 38226 24565 0 chany_top_out[11]
rlabel metal1 10442 35802 10442 35802 0 chany_top_out[12]
rlabel metal1 4968 34170 4968 34170 0 chany_top_out[13]
rlabel metal2 18078 1520 18078 1520 0 chany_top_out[14]
rlabel metal2 46 1656 46 1656 0 chany_top_out[15]
rlabel metal2 23230 1520 23230 1520 0 chany_top_out[16]
rlabel metal1 12926 34918 12926 34918 0 chany_top_out[17]
rlabel metal2 21942 38158 21942 38158 0 chany_top_out[18]
rlabel metal1 33626 37094 33626 37094 0 chany_top_out[1]
rlabel metal3 1188 26588 1188 26588 0 chany_top_out[2]
rlabel metal3 1188 22508 1188 22508 0 chany_top_out[3]
rlabel metal2 1334 1520 1334 1520 0 chany_top_out[4]
rlabel metal1 37536 37094 37536 37094 0 chany_top_out[5]
rlabel metal1 29486 37094 29486 37094 0 chany_top_out[6]
rlabel metal2 16790 1520 16790 1520 0 chany_top_out[7]
rlabel metal1 37306 36346 37306 36346 0 chany_top_out[8]
rlabel metal2 38226 3417 38226 3417 0 chany_top_out[9]
rlabel metal3 1188 10268 1188 10268 0 left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal2 38226 21233 38226 21233 0 left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal2 6486 1520 6486 1520 0 left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal2 12926 1520 12926 1520 0 left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal2 20010 1520 20010 1520 0 left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_
rlabel metal2 38226 23341 38226 23341 0 left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_
rlabel metal2 21298 1520 21298 1520 0 left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_
rlabel metal1 32384 37094 32384 37094 0 left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_
rlabel metal2 20746 32640 20746 32640 0 mem_left_ipin_0.DFFR_0_.Q
rlabel metal1 9062 33286 9062 33286 0 mem_left_ipin_0.DFFR_1_.Q
rlabel metal1 5198 32946 5198 32946 0 mem_left_ipin_0.DFFR_2_.Q
rlabel metal2 16330 36941 16330 36941 0 mem_left_ipin_0.DFFR_3_.Q
rlabel metal2 20746 31127 20746 31127 0 mem_left_ipin_0.DFFR_4_.Q
rlabel metal1 7084 33898 7084 33898 0 mem_left_ipin_0.DFFR_5_.Q
rlabel metal1 5382 34102 5382 34102 0 mem_left_ipin_1.DFFR_0_.Q
rlabel metal1 6486 34646 6486 34646 0 mem_left_ipin_1.DFFR_1_.Q
rlabel metal1 5520 31722 5520 31722 0 mem_left_ipin_1.DFFR_2_.Q
rlabel metal1 1932 37162 1932 37162 0 mem_left_ipin_1.DFFR_3_.Q
rlabel metal2 3358 35088 3358 35088 0 mem_left_ipin_1.DFFR_4_.Q
rlabel metal1 5244 33082 5244 33082 0 mem_left_ipin_1.DFFR_5_.Q
rlabel metal1 15778 28050 15778 28050 0 mem_left_ipin_2.DFFR_0_.Q
rlabel metal1 13938 28934 13938 28934 0 mem_left_ipin_2.DFFR_1_.Q
rlabel metal1 14214 31348 14214 31348 0 mem_left_ipin_2.DFFR_2_.Q
rlabel metal1 7176 36074 7176 36074 0 mem_left_ipin_2.DFFR_3_.Q
rlabel metal2 11638 36006 11638 36006 0 mem_left_ipin_2.DFFR_4_.Q
rlabel metal2 22770 37060 22770 37060 0 mem_left_ipin_2.DFFR_5_.Q
rlabel metal1 13386 21522 13386 21522 0 mem_right_ipin_0.DFFR_0_.Q
rlabel metal2 11546 21369 11546 21369 0 mem_right_ipin_0.DFFR_1_.Q
rlabel metal1 6026 21658 6026 21658 0 mem_right_ipin_0.DFFR_2_.Q
rlabel metal1 3404 31858 3404 31858 0 mem_right_ipin_0.DFFR_3_.Q
rlabel metal2 2852 31994 2852 31994 0 mem_right_ipin_0.DFFR_4_.Q
rlabel metal1 4094 29070 4094 29070 0 mem_right_ipin_0.DFFR_5_.Q
rlabel metal1 7268 22066 7268 22066 0 mem_right_ipin_1.DFFR_0_.Q
rlabel metal2 12834 32249 12834 32249 0 mem_right_ipin_1.DFFR_1_.Q
rlabel metal1 22402 28118 22402 28118 0 mem_right_ipin_1.DFFR_2_.Q
rlabel metal4 12604 31348 12604 31348 0 mem_right_ipin_1.DFFR_3_.Q
rlabel metal1 4968 36074 4968 36074 0 mem_right_ipin_1.DFFR_4_.Q
rlabel metal1 24725 29682 24725 29682 0 mem_right_ipin_1.DFFR_5_.Q
rlabel metal1 22448 27030 22448 27030 0 mem_right_ipin_2.DFFR_0_.Q
rlabel metal1 2208 20026 2208 20026 0 mem_right_ipin_2.DFFR_1_.Q
rlabel metal1 20838 33082 20838 33082 0 mem_right_ipin_2.DFFR_2_.Q
rlabel metal3 5612 31892 5612 31892 0 mem_right_ipin_2.DFFR_3_.Q
rlabel metal1 2392 35598 2392 35598 0 mem_right_ipin_2.DFFR_4_.Q
rlabel metal1 4278 35530 4278 35530 0 mem_right_ipin_2.DFFR_5_.Q
rlabel metal1 4876 22066 4876 22066 0 mem_right_ipin_3.DFFR_0_.Q
rlabel metal1 4554 32334 4554 32334 0 mem_right_ipin_3.DFFR_1_.Q
rlabel metal1 10626 32912 10626 32912 0 mem_right_ipin_3.DFFR_2_.Q
rlabel via2 1610 20587 1610 20587 0 mem_right_ipin_3.DFFR_3_.Q
rlabel metal1 3358 21658 3358 21658 0 mem_right_ipin_3.DFFR_4_.Q
rlabel metal2 3450 33660 3450 33660 0 mem_right_ipin_3.DFFR_5_.Q
rlabel metal1 14812 33966 14812 33966 0 mem_right_ipin_4.DFFR_0_.Q
rlabel metal1 8970 30634 8970 30634 0 mem_right_ipin_4.DFFR_1_.Q
rlabel metal1 15272 35734 15272 35734 0 mem_right_ipin_4.DFFR_2_.Q
rlabel metal2 21482 35360 21482 35360 0 mem_right_ipin_4.DFFR_3_.Q
rlabel metal1 5382 35462 5382 35462 0 mem_right_ipin_4.DFFR_4_.Q
rlabel metal1 10258 34986 10258 34986 0 mem_right_ipin_4.DFFR_5_.Q
rlabel metal2 12650 33286 12650 33286 0 mem_right_ipin_5.DFFR_0_.Q
rlabel metal1 14214 32776 14214 32776 0 mem_right_ipin_5.DFFR_1_.Q
rlabel metal1 20102 26384 20102 26384 0 mem_right_ipin_5.DFFR_2_.Q
rlabel via1 14299 36550 14299 36550 0 mem_right_ipin_5.DFFR_3_.Q
rlabel metal1 15962 36550 15962 36550 0 mem_right_ipin_5.DFFR_4_.Q
rlabel metal2 15962 30141 15962 30141 0 mem_right_ipin_5.DFFR_5_.Q
rlabel metal1 13754 23086 13754 23086 0 mem_right_ipin_6.DFFR_0_.Q
rlabel metal1 17710 21930 17710 21930 0 mem_right_ipin_6.DFFR_1_.Q
rlabel metal1 18032 21114 18032 21114 0 mem_right_ipin_6.DFFR_2_.Q
rlabel metal1 11454 35734 11454 35734 0 mem_right_ipin_6.DFFR_3_.Q
rlabel metal1 13432 34510 13432 34510 0 mem_right_ipin_6.DFFR_4_.Q
rlabel metal2 12006 33898 12006 33898 0 mem_right_ipin_6.DFFR_5_.Q
rlabel metal1 13478 33422 13478 33422 0 mem_right_ipin_7.DFFR_0_.Q
rlabel metal1 12788 30634 12788 30634 0 mem_right_ipin_7.DFFR_1_.Q
rlabel metal1 14858 24174 14858 24174 0 mem_right_ipin_7.DFFR_2_.Q
rlabel metal2 9614 35632 9614 35632 0 mem_right_ipin_7.DFFR_3_.Q
rlabel metal2 14582 37094 14582 37094 0 mem_right_ipin_7.DFFR_4_.Q
rlabel metal1 14904 28594 14904 28594 0 mux_left_ipin_0.INVTX1_0_.out
rlabel metal1 13938 29172 13938 29172 0 mux_left_ipin_0.INVTX1_1_.out
rlabel metal1 15226 33898 15226 33898 0 mux_left_ipin_0.INVTX1_2_.out
rlabel metal1 9108 27438 9108 27438 0 mux_left_ipin_0.INVTX1_3_.out
rlabel metal2 10350 26588 10350 26588 0 mux_left_ipin_0.INVTX1_4_.out
rlabel metal1 4830 28730 4830 28730 0 mux_left_ipin_0.INVTX1_5_.out
rlabel metal1 14674 34510 14674 34510 0 mux_left_ipin_0.INVTX1_6_.out
rlabel metal1 9108 24106 9108 24106 0 mux_left_ipin_0.INVTX1_7_.out
rlabel metal2 16606 33014 16606 33014 0 mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 14122 29682 14122 29682 0 mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 10856 28662 10856 28662 0 mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 21022 3026 21022 3026 0 mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 23391 27506 23391 27506 0 mux_left_ipin_1.INVTX1_2_.out
rlabel metal1 14214 26894 14214 26894 0 mux_left_ipin_1.INVTX1_3_.out
rlabel metal1 14030 25874 14030 25874 0 mux_left_ipin_1.INVTX1_4_.out
rlabel metal1 12696 24718 12696 24718 0 mux_left_ipin_1.INVTX1_5_.out
rlabel metal1 7360 25262 7360 25262 0 mux_left_ipin_1.INVTX1_6_.out
rlabel metal2 9154 24956 9154 24956 0 mux_left_ipin_1.INVTX1_7_.out
rlabel metal1 13570 28118 13570 28118 0 mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 9154 25738 9154 25738 0 mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 7958 25874 7958 25874 0 mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 7222 17170 7222 17170 0 mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 15594 24990 15594 24990 0 mux_left_ipin_2.INVTX1_2_.out
rlabel metal1 15088 21998 15088 21998 0 mux_left_ipin_2.INVTX1_3_.out
rlabel metal1 25967 26350 25967 26350 0 mux_left_ipin_2.INVTX1_4_.out
rlabel metal2 29486 29886 29486 29886 0 mux_left_ipin_2.INVTX1_5_.out
rlabel metal2 14674 27778 14674 27778 0 mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 16238 30974 16238 30974 0 mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 18814 33184 18814 33184 0 mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 15088 24242 15088 24242 0 mux_right_ipin_0.INVTX1_2_.out
rlabel metal2 17802 18598 17802 18598 0 mux_right_ipin_0.INVTX1_3_.out
rlabel metal1 15180 20842 15180 20842 0 mux_right_ipin_0.INVTX1_4_.out
rlabel metal1 18860 17306 18860 17306 0 mux_right_ipin_0.INVTX1_5_.out
rlabel metal1 12236 10778 12236 10778 0 mux_right_ipin_0.INVTX1_6_.out
rlabel metal1 11960 20978 11960 20978 0 mux_right_ipin_0.INVTX1_7_.out
rlabel metal1 11546 22066 11546 22066 0 mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 14122 20978 14122 20978 0 mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 11684 21658 11684 21658 0 mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 11040 20366 11040 20366 0 mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 17986 28594 17986 28594 0 mux_right_ipin_1.INVTX1_2_.out
rlabel metal1 18216 28186 18216 28186 0 mux_right_ipin_1.INVTX1_3_.out
rlabel metal1 22724 10778 22724 10778 0 mux_right_ipin_1.INVTX1_4_.out
rlabel metal1 19688 26894 19688 26894 0 mux_right_ipin_1.INVTX1_5_.out
rlabel metal1 19504 18938 19504 18938 0 mux_right_ipin_1.INVTX1_6_.out
rlabel metal1 16100 25806 16100 25806 0 mux_right_ipin_1.INVTX1_7_.out
rlabel metal1 17480 24650 17480 24650 0 mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 18906 27812 18906 27812 0 mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 19366 25738 19366 25738 0 mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 28014 25330 28014 25330 0 mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 17526 33116 17526 33116 0 mux_right_ipin_2.INVTX1_2_.out
rlabel metal1 10396 20570 10396 20570 0 mux_right_ipin_2.INVTX1_3_.out
rlabel metal1 17618 34646 17618 34646 0 mux_right_ipin_2.INVTX1_6_.out
rlabel metal2 4094 28322 4094 28322 0 mux_right_ipin_2.INVTX1_7_.out
rlabel metal1 17710 32266 17710 32266 0 mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 16100 28594 16100 28594 0 mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 12006 28424 12006 28424 0 mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 8602 15470 8602 15470 0 mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 15226 31025 15226 31025 0 mux_right_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 9798 26928 9798 26928 0 mux_right_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 8326 25738 8326 25738 0 mux_right_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 9614 11118 9614 11118 0 mux_right_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 14260 30158 14260 30158 0 mux_right_ipin_4.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 13754 26282 13754 26282 0 mux_right_ipin_4.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 9936 25330 9936 25330 0 mux_right_ipin_4.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 16882 10132 16882 10132 0 mux_right_ipin_4.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 26289 26418 26289 26418 0 mux_right_ipin_5.INVTX1_4_.out
rlabel metal1 14214 24038 14214 24038 0 mux_right_ipin_5.INVTX1_5_.out
rlabel metal2 14122 22066 14122 22066 0 mux_right_ipin_5.INVTX1_6_.out
rlabel metal1 18262 30634 18262 30634 0 mux_right_ipin_5.INVTX1_7_.out
rlabel metal2 14950 26214 14950 26214 0 mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 15134 26792 15134 26792 0 mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 17618 29920 17618 29920 0 mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 22126 25194 22126 25194 0 mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 14214 22066 14214 22066 0 mux_right_ipin_6.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 16721 21318 16721 21318 0 mux_right_ipin_6.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 13570 20570 13570 20570 0 mux_right_ipin_6.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 19320 10642 19320 10642 0 mux_right_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 17112 31858 17112 31858 0 mux_right_ipin_7.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 19366 25772 19366 25772 0 mux_right_ipin_7.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 20470 29376 20470 29376 0 mux_right_ipin_7.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 18262 31552 18262 31552 0 mux_right_ipin_7.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 37904 27030 37904 27030 0 net1
rlabel metal1 17526 37230 17526 37230 0 net10
rlabel metal1 20056 27506 20056 27506 0 net100
rlabel metal2 22770 36448 22770 36448 0 net101
rlabel metal1 2622 34646 2622 34646 0 net11
rlabel metal1 25070 27438 25070 27438 0 net12
rlabel metal1 15456 2550 15456 2550 0 net13
rlabel metal1 1886 23086 1886 23086 0 net14
rlabel metal2 16698 20434 16698 20434 0 net15
rlabel metal2 17894 35513 17894 35513 0 net16
rlabel metal2 15042 35173 15042 35173 0 net17
rlabel metal2 13432 21420 13432 21420 0 net18
rlabel metal1 38272 5882 38272 5882 0 net19
rlabel metal2 22862 28186 22862 28186 0 net2
rlabel metal1 19044 3026 19044 3026 0 net20
rlabel metal1 3818 21522 3818 21522 0 net21
rlabel metal1 37904 3094 37904 3094 0 net22
rlabel metal1 37858 16082 37858 16082 0 net23
rlabel metal1 3818 2550 3818 2550 0 net24
rlabel metal1 3312 13974 3312 13974 0 net25
rlabel via2 1886 31195 1886 31195 0 net26
rlabel metal2 11270 19550 11270 19550 0 net27
rlabel metal1 3680 14586 3680 14586 0 net28
rlabel metal1 5106 18938 5106 18938 0 net29
rlabel metal2 37306 2788 37306 2788 0 net3
rlabel metal2 8694 2822 8694 2822 0 net30
rlabel metal2 12006 2601 12006 2601 0 net31
rlabel metal2 33718 12886 33718 12886 0 net32
rlabel metal1 37950 12206 37950 12206 0 net33
rlabel metal2 38088 19788 38088 19788 0 net34
rlabel metal1 10488 20774 10488 20774 0 net35
rlabel metal2 13386 24412 13386 24412 0 net36
rlabel metal1 15226 19312 15226 19312 0 net37
rlabel metal2 27278 23562 27278 23562 0 net38
rlabel metal1 24748 6290 24748 6290 0 net39
rlabel metal1 37996 25262 37996 25262 0 net4
rlabel metal2 20470 36958 20470 36958 0 net40
rlabel metal1 37996 36142 37996 36142 0 net41
rlabel metal1 32752 28662 32752 28662 0 net42
rlabel metal2 17158 31892 17158 31892 0 net43
rlabel metal2 38042 31110 38042 31110 0 net44
rlabel metal1 2116 28050 2116 28050 0 net45
rlabel metal1 21298 29274 21298 29274 0 net46
rlabel metal2 37306 30532 37306 30532 0 net47
rlabel via2 3358 20043 3358 20043 0 net48
rlabel metal1 1932 3026 1932 3026 0 net49
rlabel metal1 35834 37196 35834 37196 0 net5
rlabel metal1 3542 18598 3542 18598 0 net50
rlabel metal2 8602 2618 8602 2618 0 net51
rlabel metal1 18446 36346 18446 36346 0 net52
rlabel metal2 17664 34204 17664 34204 0 net53
rlabel metal2 38042 10506 38042 10506 0 net54
rlabel metal1 24564 27098 24564 27098 0 net55
rlabel metal1 19504 21046 19504 21046 0 net56
rlabel via1 20654 3077 20654 3077 0 net57
rlabel metal2 14306 18972 14306 18972 0 net58
rlabel metal1 37766 35666 37766 35666 0 net59
rlabel metal1 2392 3638 2392 3638 0 net6
rlabel metal1 25116 2414 25116 2414 0 net60
rlabel metal1 1886 24718 1886 24718 0 net61
rlabel metal1 29486 2414 29486 2414 0 net62
rlabel metal2 38042 24956 38042 24956 0 net63
rlabel metal2 12558 37145 12558 37145 0 net64
rlabel metal1 4738 33966 4738 33966 0 net65
rlabel metal2 18170 5746 18170 5746 0 net66
rlabel metal2 4738 2686 4738 2686 0 net67
rlabel metal1 22954 2414 22954 2414 0 net68
rlabel metal2 13294 35530 13294 35530 0 net69
rlabel metal1 15042 19210 15042 19210 0 net7
rlabel metal1 19412 35802 19412 35802 0 net70
rlabel metal1 33948 37230 33948 37230 0 net71
rlabel metal1 4140 24310 4140 24310 0 net72
rlabel metal2 1886 22780 1886 22780 0 net73
rlabel metal1 2162 2414 2162 2414 0 net74
rlabel metal2 36846 36958 36846 36958 0 net75
rlabel metal1 27922 36890 27922 36890 0 net76
rlabel metal2 16882 5644 16882 5644 0 net77
rlabel metal1 37720 36142 37720 36142 0 net78
rlabel metal1 37444 3366 37444 3366 0 net79
rlabel metal1 12512 3026 12512 3026 0 net8
rlabel metal1 2162 10642 2162 10642 0 net80
rlabel metal2 36846 23324 36846 23324 0 net81
rlabel metal2 6854 8874 6854 8874 0 net82
rlabel metal1 11960 2414 11960 2414 0 net83
rlabel metal1 19366 2414 19366 2414 0 net84
rlabel metal2 37306 24446 37306 24446 0 net85
rlabel metal1 20562 10506 20562 10506 0 net86
rlabel metal2 32338 36992 32338 36992 0 net87
rlabel metal3 17204 36584 17204 36584 0 net88
rlabel metal2 23414 2584 23414 2584 0 net89
rlabel metal1 21298 18598 21298 18598 0 net9
rlabel metal1 4324 12818 4324 12818 0 net90
rlabel metal2 10350 27234 10350 27234 0 net91
rlabel metal1 8510 23154 8510 23154 0 net92
rlabel metal2 10534 21692 10534 21692 0 net93
rlabel metal2 20010 28220 20010 28220 0 net94
rlabel metal2 15778 33184 15778 33184 0 net95
rlabel metal2 5658 25568 5658 25568 0 net96
rlabel metal1 9982 24718 9982 24718 0 net97
rlabel metal1 16330 23630 16330 23630 0 net98
rlabel metal1 14904 19482 14904 19482 0 net99
rlabel metal1 30544 37230 30544 37230 0 pReset
rlabel metal2 1702 36686 1702 36686 0 prog_clk
rlabel metal1 7682 35802 7682 35802 0 right_grid_left_width_0_height_0_subtile_0__pin_I_11_
rlabel metal2 26450 1520 26450 1520 0 right_grid_left_width_0_height_0_subtile_0__pin_I_3_
rlabel metal3 1188 12308 1188 12308 0 right_grid_left_width_0_height_0_subtile_0__pin_I_7_
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
