magic
tech sky130A
magscale 1 2
timestamp 1674174823
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 14 2128 39638 38344
<< metal2 >>
rect 662 39200 718 39800
rect 1950 39200 2006 39800
rect 2594 39200 2650 39800
rect 3882 39200 3938 39800
rect 5170 39200 5226 39800
rect 5814 39200 5870 39800
rect 7102 39200 7158 39800
rect 8390 39200 8446 39800
rect 9034 39200 9090 39800
rect 10322 39200 10378 39800
rect 11610 39200 11666 39800
rect 12254 39200 12310 39800
rect 13542 39200 13598 39800
rect 14830 39200 14886 39800
rect 16118 39200 16174 39800
rect 16762 39200 16818 39800
rect 18050 39200 18106 39800
rect 19338 39200 19394 39800
rect 19982 39200 20038 39800
rect 21270 39200 21326 39800
rect 22558 39200 22614 39800
rect 23202 39200 23258 39800
rect 24490 39200 24546 39800
rect 25778 39200 25834 39800
rect 26422 39200 26478 39800
rect 27710 39200 27766 39800
rect 28998 39200 29054 39800
rect 29642 39200 29698 39800
rect 30930 39200 30986 39800
rect 32218 39200 32274 39800
rect 32862 39200 32918 39800
rect 34150 39200 34206 39800
rect 35438 39200 35494 39800
rect 36082 39200 36138 39800
rect 37370 39200 37426 39800
rect 38658 39200 38714 39800
rect 39302 39200 39358 39800
rect 18 200 74 800
rect 662 200 718 800
rect 1950 200 2006 800
rect 3238 200 3294 800
rect 3882 200 3938 800
rect 5170 200 5226 800
rect 6458 200 6514 800
rect 7102 200 7158 800
rect 8390 200 8446 800
rect 9678 200 9734 800
rect 10322 200 10378 800
rect 11610 200 11666 800
rect 12898 200 12954 800
rect 13542 200 13598 800
rect 14830 200 14886 800
rect 16118 200 16174 800
rect 16762 200 16818 800
rect 18050 200 18106 800
rect 19338 200 19394 800
rect 19982 200 20038 800
rect 21270 200 21326 800
rect 22558 200 22614 800
rect 23202 200 23258 800
rect 24490 200 24546 800
rect 25778 200 25834 800
rect 27066 200 27122 800
rect 27710 200 27766 800
rect 28998 200 29054 800
rect 30286 200 30342 800
rect 30930 200 30986 800
rect 32218 200 32274 800
rect 33506 200 33562 800
rect 34150 200 34206 800
rect 35438 200 35494 800
rect 36726 200 36782 800
rect 37370 200 37426 800
rect 38658 200 38714 800
<< obsm2 >>
rect 20 39144 606 39545
rect 774 39144 1894 39545
rect 2062 39144 2538 39545
rect 2706 39144 3826 39545
rect 3994 39144 5114 39545
rect 5282 39144 5758 39545
rect 5926 39144 7046 39545
rect 7214 39144 8334 39545
rect 8502 39144 8978 39545
rect 9146 39144 10266 39545
rect 10434 39144 11554 39545
rect 11722 39144 12198 39545
rect 12366 39144 13486 39545
rect 13654 39144 14774 39545
rect 14942 39144 16062 39545
rect 16230 39144 16706 39545
rect 16874 39144 17994 39545
rect 18162 39144 19282 39545
rect 19450 39144 19926 39545
rect 20094 39144 21214 39545
rect 21382 39144 22502 39545
rect 22670 39144 23146 39545
rect 23314 39144 24434 39545
rect 24602 39144 25722 39545
rect 25890 39144 26366 39545
rect 26534 39144 27654 39545
rect 27822 39144 28942 39545
rect 29110 39144 29586 39545
rect 29754 39144 30874 39545
rect 31042 39144 32162 39545
rect 32330 39144 32806 39545
rect 32974 39144 34094 39545
rect 34262 39144 35382 39545
rect 35550 39144 36026 39545
rect 36194 39144 37314 39545
rect 37482 39144 38602 39545
rect 38770 39144 39246 39545
rect 39414 39144 39632 39545
rect 20 856 39632 39144
rect 130 144 606 856
rect 774 144 1894 856
rect 2062 144 3182 856
rect 3350 144 3826 856
rect 3994 144 5114 856
rect 5282 144 6402 856
rect 6570 144 7046 856
rect 7214 144 8334 856
rect 8502 144 9622 856
rect 9790 144 10266 856
rect 10434 144 11554 856
rect 11722 144 12842 856
rect 13010 144 13486 856
rect 13654 144 14774 856
rect 14942 144 16062 856
rect 16230 144 16706 856
rect 16874 144 17994 856
rect 18162 144 19282 856
rect 19450 144 19926 856
rect 20094 144 21214 856
rect 21382 144 22502 856
rect 22670 144 23146 856
rect 23314 144 24434 856
rect 24602 144 25722 856
rect 25890 144 27010 856
rect 27178 144 27654 856
rect 27822 144 28942 856
rect 29110 144 30230 856
rect 30398 144 30874 856
rect 31042 144 32162 856
rect 32330 144 33450 856
rect 33618 144 34094 856
rect 34262 144 35382 856
rect 35550 144 36670 856
rect 36838 144 37314 856
rect 37482 144 38602 856
rect 38770 144 39632 856
rect 20 31 39632 144
<< metal3 >>
rect 200 39448 800 39568
rect 200 38768 800 38888
rect 39200 38768 39800 38888
rect 200 37408 800 37528
rect 39200 37408 39800 37528
rect 200 36048 800 36168
rect 39200 36048 39800 36168
rect 200 35368 800 35488
rect 39200 35368 39800 35488
rect 200 34008 800 34128
rect 39200 34008 39800 34128
rect 200 32648 800 32768
rect 39200 32648 39800 32768
rect 200 31968 800 32088
rect 39200 31968 39800 32088
rect 200 30608 800 30728
rect 39200 30608 39800 30728
rect 200 29248 800 29368
rect 39200 29248 39800 29368
rect 200 28568 800 28688
rect 39200 28568 39800 28688
rect 200 27208 800 27328
rect 39200 27208 39800 27328
rect 200 25848 800 25968
rect 39200 25848 39800 25968
rect 39200 25168 39800 25288
rect 200 24488 800 24608
rect 200 23808 800 23928
rect 39200 23808 39800 23928
rect 200 22448 800 22568
rect 39200 22448 39800 22568
rect 39200 21768 39800 21888
rect 200 21088 800 21208
rect 200 20408 800 20528
rect 39200 20408 39800 20528
rect 200 19048 800 19168
rect 39200 19048 39800 19168
rect 39200 18368 39800 18488
rect 200 17688 800 17808
rect 200 17008 800 17128
rect 39200 17008 39800 17128
rect 200 15648 800 15768
rect 39200 15648 39800 15768
rect 39200 14968 39800 15088
rect 200 14288 800 14408
rect 200 13608 800 13728
rect 39200 13608 39800 13728
rect 200 12248 800 12368
rect 39200 12248 39800 12368
rect 200 10888 800 11008
rect 39200 10888 39800 11008
rect 200 10208 800 10328
rect 39200 10208 39800 10328
rect 200 8848 800 8968
rect 39200 8848 39800 8968
rect 200 7488 800 7608
rect 39200 7488 39800 7608
rect 200 6808 800 6928
rect 39200 6808 39800 6928
rect 200 5448 800 5568
rect 39200 5448 39800 5568
rect 200 4088 800 4208
rect 39200 4088 39800 4208
rect 200 3408 800 3528
rect 39200 3408 39800 3528
rect 200 2048 800 2168
rect 39200 2048 39800 2168
rect 200 688 800 808
rect 39200 688 39800 808
rect 39200 8 39800 128
<< obsm3 >>
rect 880 39368 39200 39541
rect 800 38968 39200 39368
rect 880 38688 39120 38968
rect 800 37608 39200 38688
rect 880 37328 39120 37608
rect 800 36248 39200 37328
rect 880 35968 39120 36248
rect 800 35568 39200 35968
rect 880 35288 39120 35568
rect 800 34208 39200 35288
rect 880 33928 39120 34208
rect 800 32848 39200 33928
rect 880 32568 39120 32848
rect 800 32168 39200 32568
rect 880 31888 39120 32168
rect 800 30808 39200 31888
rect 880 30528 39120 30808
rect 800 29448 39200 30528
rect 880 29168 39120 29448
rect 800 28768 39200 29168
rect 880 28488 39120 28768
rect 800 27408 39200 28488
rect 880 27128 39120 27408
rect 800 26048 39200 27128
rect 880 25768 39120 26048
rect 800 25368 39200 25768
rect 800 25088 39120 25368
rect 800 24688 39200 25088
rect 880 24408 39200 24688
rect 800 24008 39200 24408
rect 880 23728 39120 24008
rect 800 22648 39200 23728
rect 880 22368 39120 22648
rect 800 21968 39200 22368
rect 800 21688 39120 21968
rect 800 21288 39200 21688
rect 880 21008 39200 21288
rect 800 20608 39200 21008
rect 880 20328 39120 20608
rect 800 19248 39200 20328
rect 880 18968 39120 19248
rect 800 18568 39200 18968
rect 800 18288 39120 18568
rect 800 17888 39200 18288
rect 880 17608 39200 17888
rect 800 17208 39200 17608
rect 880 16928 39120 17208
rect 800 15848 39200 16928
rect 880 15568 39120 15848
rect 800 15168 39200 15568
rect 800 14888 39120 15168
rect 800 14488 39200 14888
rect 880 14208 39200 14488
rect 800 13808 39200 14208
rect 880 13528 39120 13808
rect 800 12448 39200 13528
rect 880 12168 39120 12448
rect 800 11088 39200 12168
rect 880 10808 39120 11088
rect 800 10408 39200 10808
rect 880 10128 39120 10408
rect 800 9048 39200 10128
rect 880 8768 39120 9048
rect 800 7688 39200 8768
rect 880 7408 39120 7688
rect 800 7008 39200 7408
rect 880 6728 39120 7008
rect 800 5648 39200 6728
rect 880 5368 39120 5648
rect 800 4288 39200 5368
rect 880 4008 39120 4288
rect 800 3608 39200 4008
rect 880 3328 39120 3608
rect 800 2248 39200 3328
rect 880 1968 39120 2248
rect 800 888 39200 1968
rect 880 608 39120 888
rect 800 208 39200 608
rect 800 35 39120 208
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< obsm4 >>
rect 12939 9827 19488 36821
rect 19968 9827 34848 36821
rect 35328 9827 36925 36821
<< labels >>
rlabel metal3 s 200 19048 800 19168 6 bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 1 nsew signal input
rlabel metal3 s 200 7488 800 7608 6 bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 2 nsew signal input
rlabel metal2 s 5170 39200 5226 39800 6 bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 3 nsew signal input
rlabel metal3 s 200 5448 800 5568 6 bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 4 nsew signal input
rlabel metal2 s 35438 200 35494 800 6 bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_
port 5 nsew signal input
rlabel metal2 s 25778 200 25834 800 6 bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_
port 6 nsew signal input
rlabel metal3 s 200 22448 800 22568 6 bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_
port 7 nsew signal input
rlabel metal3 s 200 6808 800 6928 6 bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_
port 8 nsew signal input
rlabel metal2 s 18050 39200 18106 39800 6 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
port 9 nsew signal input
rlabel metal3 s 200 38768 800 38888 6 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
port 10 nsew signal input
rlabel metal2 s 12898 200 12954 800 6 ccff_head
port 11 nsew signal input
rlabel metal2 s 28998 200 29054 800 6 ccff_tail
port 12 nsew signal output
rlabel metal2 s 25778 39200 25834 39800 6 chanx_right_in[0]
port 13 nsew signal input
rlabel metal2 s 5814 39200 5870 39800 6 chanx_right_in[10]
port 14 nsew signal input
rlabel metal2 s 24490 200 24546 800 6 chanx_right_in[11]
port 15 nsew signal input
rlabel metal2 s 9034 39200 9090 39800 6 chanx_right_in[12]
port 16 nsew signal input
rlabel metal2 s 19982 200 20038 800 6 chanx_right_in[13]
port 17 nsew signal input
rlabel metal3 s 200 17008 800 17128 6 chanx_right_in[14]
port 18 nsew signal input
rlabel metal3 s 200 2048 800 2168 6 chanx_right_in[15]
port 19 nsew signal input
rlabel metal2 s 27710 39200 27766 39800 6 chanx_right_in[16]
port 20 nsew signal input
rlabel metal2 s 11610 200 11666 800 6 chanx_right_in[17]
port 21 nsew signal input
rlabel metal3 s 39200 31968 39800 32088 6 chanx_right_in[18]
port 22 nsew signal input
rlabel metal3 s 39200 27208 39800 27328 6 chanx_right_in[1]
port 23 nsew signal input
rlabel metal2 s 9678 200 9734 800 6 chanx_right_in[2]
port 24 nsew signal input
rlabel metal3 s 200 688 800 808 6 chanx_right_in[3]
port 25 nsew signal input
rlabel metal3 s 39200 8848 39800 8968 6 chanx_right_in[4]
port 26 nsew signal input
rlabel metal2 s 14830 39200 14886 39800 6 chanx_right_in[5]
port 27 nsew signal input
rlabel metal3 s 39200 30608 39800 30728 6 chanx_right_in[6]
port 28 nsew signal input
rlabel metal3 s 39200 28568 39800 28688 6 chanx_right_in[7]
port 29 nsew signal input
rlabel metal2 s 32218 39200 32274 39800 6 chanx_right_in[8]
port 30 nsew signal input
rlabel metal2 s 18050 200 18106 800 6 chanx_right_in[9]
port 31 nsew signal input
rlabel metal2 s 36082 39200 36138 39800 6 chanx_right_out[0]
port 32 nsew signal output
rlabel metal3 s 39200 12248 39800 12368 6 chanx_right_out[10]
port 33 nsew signal output
rlabel metal2 s 33506 200 33562 800 6 chanx_right_out[11]
port 34 nsew signal output
rlabel metal3 s 200 30608 800 30728 6 chanx_right_out[12]
port 35 nsew signal output
rlabel metal3 s 200 15648 800 15768 6 chanx_right_out[13]
port 36 nsew signal output
rlabel metal3 s 39200 2048 39800 2168 6 chanx_right_out[14]
port 37 nsew signal output
rlabel metal2 s 19982 39200 20038 39800 6 chanx_right_out[15]
port 38 nsew signal output
rlabel metal3 s 39200 35368 39800 35488 6 chanx_right_out[16]
port 39 nsew signal output
rlabel metal3 s 39200 8 39800 128 6 chanx_right_out[17]
port 40 nsew signal output
rlabel metal2 s 19338 39200 19394 39800 6 chanx_right_out[18]
port 41 nsew signal output
rlabel metal2 s 34150 200 34206 800 6 chanx_right_out[1]
port 42 nsew signal output
rlabel metal2 s 30930 39200 30986 39800 6 chanx_right_out[2]
port 43 nsew signal output
rlabel metal2 s 34150 39200 34206 39800 6 chanx_right_out[3]
port 44 nsew signal output
rlabel metal3 s 39200 37408 39800 37528 6 chanx_right_out[4]
port 45 nsew signal output
rlabel metal2 s 16118 39200 16174 39800 6 chanx_right_out[5]
port 46 nsew signal output
rlabel metal3 s 39200 10888 39800 11008 6 chanx_right_out[6]
port 47 nsew signal output
rlabel metal3 s 39200 13608 39800 13728 6 chanx_right_out[7]
port 48 nsew signal output
rlabel metal3 s 39200 19048 39800 19168 6 chanx_right_out[8]
port 49 nsew signal output
rlabel metal2 s 27710 200 27766 800 6 chanx_right_out[9]
port 50 nsew signal output
rlabel metal3 s 39200 38768 39800 38888 6 chany_bottom_in[0]
port 51 nsew signal input
rlabel metal3 s 39200 32648 39800 32768 6 chany_bottom_in[10]
port 52 nsew signal input
rlabel metal2 s 24490 39200 24546 39800 6 chany_bottom_in[11]
port 53 nsew signal input
rlabel metal2 s 12254 39200 12310 39800 6 chany_bottom_in[12]
port 54 nsew signal input
rlabel metal3 s 39200 23808 39800 23928 6 chany_bottom_in[13]
port 55 nsew signal input
rlabel metal2 s 8390 39200 8446 39800 6 chany_bottom_in[14]
port 56 nsew signal input
rlabel metal2 s 11610 39200 11666 39800 6 chany_bottom_in[15]
port 57 nsew signal input
rlabel metal2 s 22558 39200 22614 39800 6 chany_bottom_in[16]
port 58 nsew signal input
rlabel metal2 s 10322 200 10378 800 6 chany_bottom_in[17]
port 59 nsew signal input
rlabel metal2 s 2594 39200 2650 39800 6 chany_bottom_in[18]
port 60 nsew signal input
rlabel metal3 s 39200 14968 39800 15088 6 chany_bottom_in[1]
port 61 nsew signal input
rlabel metal2 s 3882 39200 3938 39800 6 chany_bottom_in[2]
port 62 nsew signal input
rlabel metal3 s 39200 688 39800 808 6 chany_bottom_in[3]
port 63 nsew signal input
rlabel metal3 s 200 14288 800 14408 6 chany_bottom_in[4]
port 64 nsew signal input
rlabel metal3 s 39200 7488 39800 7608 6 chany_bottom_in[5]
port 65 nsew signal input
rlabel metal3 s 200 28568 800 28688 6 chany_bottom_in[6]
port 66 nsew signal input
rlabel metal2 s 16762 200 16818 800 6 chany_bottom_in[7]
port 67 nsew signal input
rlabel metal3 s 200 21088 800 21208 6 chany_bottom_in[8]
port 68 nsew signal input
rlabel metal2 s 16118 200 16174 800 6 chany_bottom_in[9]
port 69 nsew signal input
rlabel metal3 s 200 24488 800 24608 6 chany_bottom_out[0]
port 70 nsew signal output
rlabel metal2 s 32862 39200 32918 39800 6 chany_bottom_out[10]
port 71 nsew signal output
rlabel metal3 s 200 32648 800 32768 6 chany_bottom_out[11]
port 72 nsew signal output
rlabel metal2 s 30286 200 30342 800 6 chany_bottom_out[12]
port 73 nsew signal output
rlabel metal3 s 39200 25168 39800 25288 6 chany_bottom_out[13]
port 74 nsew signal output
rlabel metal3 s 39200 5448 39800 5568 6 chany_bottom_out[14]
port 75 nsew signal output
rlabel metal2 s 26422 39200 26478 39800 6 chany_bottom_out[15]
port 76 nsew signal output
rlabel metal2 s 39302 39200 39358 39800 6 chany_bottom_out[16]
port 77 nsew signal output
rlabel metal2 s 37370 39200 37426 39800 6 chany_bottom_out[17]
port 78 nsew signal output
rlabel metal2 s 662 200 718 800 6 chany_bottom_out[18]
port 79 nsew signal output
rlabel metal2 s 5170 200 5226 800 6 chany_bottom_out[1]
port 80 nsew signal output
rlabel metal2 s 38658 200 38714 800 6 chany_bottom_out[2]
port 81 nsew signal output
rlabel metal3 s 200 13608 800 13728 6 chany_bottom_out[3]
port 82 nsew signal output
rlabel metal3 s 39200 21768 39800 21888 6 chany_bottom_out[4]
port 83 nsew signal output
rlabel metal3 s 39200 15648 39800 15768 6 chany_bottom_out[5]
port 84 nsew signal output
rlabel metal2 s 16762 39200 16818 39800 6 chany_bottom_out[6]
port 85 nsew signal output
rlabel metal2 s 3238 200 3294 800 6 chany_bottom_out[7]
port 86 nsew signal output
rlabel metal3 s 39200 3408 39800 3528 6 chany_bottom_out[8]
port 87 nsew signal output
rlabel metal3 s 39200 17008 39800 17128 6 chany_bottom_out[9]
port 88 nsew signal output
rlabel metal3 s 200 27208 800 27328 6 chany_top_in[0]
port 89 nsew signal input
rlabel metal2 s 1950 39200 2006 39800 6 chany_top_in[10]
port 90 nsew signal input
rlabel metal3 s 200 25848 800 25968 6 chany_top_in[11]
port 91 nsew signal input
rlabel metal3 s 200 20408 800 20528 6 chany_top_in[12]
port 92 nsew signal input
rlabel metal3 s 200 39448 800 39568 6 chany_top_in[13]
port 93 nsew signal input
rlabel metal2 s 38658 39200 38714 39800 6 chany_top_in[14]
port 94 nsew signal input
rlabel metal2 s 8390 200 8446 800 6 chany_top_in[15]
port 95 nsew signal input
rlabel metal3 s 200 17688 800 17808 6 chany_top_in[16]
port 96 nsew signal input
rlabel metal2 s 23202 200 23258 800 6 chany_top_in[17]
port 97 nsew signal input
rlabel metal2 s 37370 200 37426 800 6 chany_top_in[18]
port 98 nsew signal input
rlabel metal2 s 13542 39200 13598 39800 6 chany_top_in[1]
port 99 nsew signal input
rlabel metal2 s 30930 200 30986 800 6 chany_top_in[2]
port 100 nsew signal input
rlabel metal2 s 3882 200 3938 800 6 chany_top_in[3]
port 101 nsew signal input
rlabel metal2 s 14830 200 14886 800 6 chany_top_in[4]
port 102 nsew signal input
rlabel metal3 s 39200 4088 39800 4208 6 chany_top_in[5]
port 103 nsew signal input
rlabel metal3 s 39200 29248 39800 29368 6 chany_top_in[6]
port 104 nsew signal input
rlabel metal3 s 39200 20408 39800 20528 6 chany_top_in[7]
port 105 nsew signal input
rlabel metal2 s 32218 200 32274 800 6 chany_top_in[8]
port 106 nsew signal input
rlabel metal3 s 200 23808 800 23928 6 chany_top_in[9]
port 107 nsew signal input
rlabel metal3 s 39200 10208 39800 10328 6 chany_top_out[0]
port 108 nsew signal output
rlabel metal3 s 200 31968 800 32088 6 chany_top_out[10]
port 109 nsew signal output
rlabel metal3 s 39200 22448 39800 22568 6 chany_top_out[11]
port 110 nsew signal output
rlabel metal3 s 39200 34008 39800 34128 6 chany_top_out[12]
port 111 nsew signal output
rlabel metal2 s 36726 200 36782 800 6 chany_top_out[13]
port 112 nsew signal output
rlabel metal3 s 39200 36048 39800 36168 6 chany_top_out[14]
port 113 nsew signal output
rlabel metal3 s 200 12248 800 12368 6 chany_top_out[15]
port 114 nsew signal output
rlabel metal3 s 200 34008 800 34128 6 chany_top_out[16]
port 115 nsew signal output
rlabel metal3 s 200 3408 800 3528 6 chany_top_out[17]
port 116 nsew signal output
rlabel metal2 s 18 200 74 800 6 chany_top_out[18]
port 117 nsew signal output
rlabel metal3 s 200 4088 800 4208 6 chany_top_out[1]
port 118 nsew signal output
rlabel metal3 s 200 37408 800 37528 6 chany_top_out[2]
port 119 nsew signal output
rlabel metal2 s 10322 39200 10378 39800 6 chany_top_out[3]
port 120 nsew signal output
rlabel metal2 s 23202 39200 23258 39800 6 chany_top_out[4]
port 121 nsew signal output
rlabel metal3 s 200 29248 800 29368 6 chany_top_out[5]
port 122 nsew signal output
rlabel metal2 s 6458 200 6514 800 6 chany_top_out[6]
port 123 nsew signal output
rlabel metal2 s 1950 200 2006 800 6 chany_top_out[7]
port 124 nsew signal output
rlabel metal3 s 200 8848 800 8968 6 chany_top_out[8]
port 125 nsew signal output
rlabel metal2 s 21270 39200 21326 39800 6 chany_top_out[9]
port 126 nsew signal output
rlabel metal2 s 19338 200 19394 800 6 pReset
port 127 nsew signal input
rlabel metal2 s 35438 39200 35494 39800 6 prog_clk
port 128 nsew signal input
rlabel metal3 s 39200 6808 39800 6928 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 129 nsew signal input
rlabel metal3 s 200 36048 800 36168 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 130 nsew signal input
rlabel metal3 s 200 10888 800 11008 6 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
port 131 nsew signal input
rlabel metal2 s 7102 200 7158 800 6 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
port 132 nsew signal input
rlabel metal2 s 13542 200 13598 800 6 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 133 nsew signal input
rlabel metal2 s 21270 200 21326 800 6 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 134 nsew signal input
rlabel metal3 s 39200 25848 39800 25968 6 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 135 nsew signal input
rlabel metal2 s 22558 200 22614 800 6 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 136 nsew signal input
rlabel metal2 s 29642 39200 29698 39800 6 top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_
port 137 nsew signal input
rlabel metal2 s 28998 39200 29054 39800 6 top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_
port 138 nsew signal input
rlabel metal2 s 662 39200 718 39800 6 top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_
port 139 nsew signal input
rlabel metal2 s 7102 39200 7158 39800 6 top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_
port 140 nsew signal input
rlabel metal2 s 27066 200 27122 800 6 top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
port 141 nsew signal input
rlabel metal3 s 200 10208 800 10328 6 top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
port 142 nsew signal input
rlabel metal3 s 200 35368 800 35488 6 vccd1
port 143 nsew signal bidirectional
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 143 nsew signal bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 143 nsew signal bidirectional
rlabel metal3 s 39200 18368 39800 18488 6 vssd1
port 144 nsew signal bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 144 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2420526
string GDS_FILE /home/baungarten/Proyectos_caravel/FPGA_3/openlane/sb_0__1_/runs/23_01_19_18_32/results/signoff/sb_0__1_.magic.gds
string GDS_START 174068
<< end >>

