// This is the unpowered netlist.
module sb_0__1_ (bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_,
    bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_,
    bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_,
    bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_,
    bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_,
    bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_,
    bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_,
    bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_,
    bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_,
    bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_,
    ccff_head,
    ccff_tail,
    pReset,
    prog_clk,
    right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_,
    right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_,
    right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_,
    right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_,
    top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_,
    top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_,
    top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_,
    top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_,
    top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_,
    top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_,
    top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_,
    top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_,
    top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_,
    top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_,
    vccd1,
    vssd1,
    chanx_right_in,
    chanx_right_out,
    chany_bottom_in,
    chany_bottom_out,
    chany_top_in,
    chany_top_out);
 input bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
 input bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
 input bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
 input bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
 input bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
 input bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
 input bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
 input bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
 input bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_;
 input bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_;
 input ccff_head;
 output ccff_tail;
 input pReset;
 input prog_clk;
 input right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
 input right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
 input right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_;
 input right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_;
 input top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
 input top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
 input top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
 input top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
 input top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
 input top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
 input top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
 input top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
 input top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_;
 input top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_;
 inout vccd1;
 inout vssd1;
 input [0:18] chanx_right_in;
 output [0:18] chanx_right_out;
 input [0:18] chany_bottom_in;
 output [0:18] chany_bottom_out;
 input [0:18] chany_top_in;
 output [0:18] chany_top_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire clknet_0_prog_clk;
 wire \mem_bottom_track_1.DFFR_0_.D ;
 wire \mem_bottom_track_1.DFFR_0_.Q ;
 wire \mem_bottom_track_1.DFFR_1_.Q ;
 wire \mem_bottom_track_1.DFFR_2_.Q ;
 wire \mem_bottom_track_1.DFFR_3_.Q ;
 wire \mem_bottom_track_1.DFFR_4_.Q ;
 wire \mem_bottom_track_1.DFFR_5_.Q ;
 wire \mem_bottom_track_1.DFFR_6_.Q ;
 wire \mem_bottom_track_1.DFFR_7_.Q ;
 wire \mem_bottom_track_17.DFFR_0_.D ;
 wire \mem_bottom_track_17.DFFR_0_.Q ;
 wire \mem_bottom_track_17.DFFR_1_.Q ;
 wire \mem_bottom_track_17.DFFR_2_.Q ;
 wire \mem_bottom_track_17.DFFR_3_.Q ;
 wire \mem_bottom_track_17.DFFR_4_.Q ;
 wire \mem_bottom_track_17.DFFR_5_.Q ;
 wire \mem_bottom_track_17.DFFR_6_.Q ;
 wire \mem_bottom_track_17.DFFR_7_.Q ;
 wire \mem_bottom_track_25.DFFR_0_.Q ;
 wire \mem_bottom_track_25.DFFR_1_.Q ;
 wire \mem_bottom_track_25.DFFR_2_.Q ;
 wire \mem_bottom_track_25.DFFR_3_.Q ;
 wire \mem_bottom_track_25.DFFR_4_.Q ;
 wire \mem_bottom_track_25.DFFR_5_.Q ;
 wire \mem_bottom_track_25.DFFR_6_.Q ;
 wire \mem_bottom_track_25.DFFR_7_.Q ;
 wire \mem_bottom_track_33.DFFR_0_.Q ;
 wire \mem_bottom_track_33.DFFR_1_.Q ;
 wire \mem_bottom_track_33.DFFR_2_.Q ;
 wire \mem_bottom_track_33.DFFR_3_.Q ;
 wire \mem_bottom_track_33.DFFR_4_.Q ;
 wire \mem_bottom_track_9.DFFR_0_.Q ;
 wire \mem_bottom_track_9.DFFR_1_.Q ;
 wire \mem_bottom_track_9.DFFR_2_.Q ;
 wire \mem_bottom_track_9.DFFR_3_.Q ;
 wire \mem_bottom_track_9.DFFR_4_.Q ;
 wire \mem_bottom_track_9.DFFR_5_.Q ;
 wire \mem_bottom_track_9.DFFR_6_.Q ;
 wire \mem_right_track_0.DFFR_0_.D ;
 wire \mem_right_track_0.DFFR_0_.Q ;
 wire \mem_right_track_0.DFFR_1_.Q ;
 wire \mem_right_track_0.DFFR_2_.Q ;
 wire \mem_right_track_0.DFFR_3_.Q ;
 wire \mem_right_track_0.DFFR_4_.Q ;
 wire \mem_right_track_0.DFFR_5_.Q ;
 wire \mem_right_track_10.DFFR_0_.D ;
 wire \mem_right_track_10.DFFR_0_.Q ;
 wire \mem_right_track_10.DFFR_1_.Q ;
 wire \mem_right_track_12.DFFR_0_.Q ;
 wire \mem_right_track_12.DFFR_1_.Q ;
 wire \mem_right_track_14.DFFR_0_.Q ;
 wire \mem_right_track_14.DFFR_1_.Q ;
 wire \mem_right_track_16.DFFR_0_.Q ;
 wire \mem_right_track_16.DFFR_1_.Q ;
 wire \mem_right_track_18.DFFR_0_.Q ;
 wire \mem_right_track_18.DFFR_1_.Q ;
 wire \mem_right_track_2.DFFR_0_.Q ;
 wire \mem_right_track_2.DFFR_1_.Q ;
 wire \mem_right_track_2.DFFR_2_.Q ;
 wire \mem_right_track_2.DFFR_3_.Q ;
 wire \mem_right_track_2.DFFR_4_.Q ;
 wire \mem_right_track_2.DFFR_5_.Q ;
 wire \mem_right_track_20.DFFR_0_.Q ;
 wire \mem_right_track_20.DFFR_1_.Q ;
 wire \mem_right_track_22.DFFR_0_.Q ;
 wire \mem_right_track_22.DFFR_1_.Q ;
 wire \mem_right_track_24.DFFR_0_.Q ;
 wire \mem_right_track_24.DFFR_1_.Q ;
 wire \mem_right_track_26.DFFR_0_.Q ;
 wire \mem_right_track_4.DFFR_0_.Q ;
 wire \mem_right_track_4.DFFR_1_.Q ;
 wire \mem_right_track_4.DFFR_2_.Q ;
 wire \mem_right_track_4.DFFR_3_.Q ;
 wire \mem_right_track_4.DFFR_4_.Q ;
 wire \mem_right_track_4.DFFR_5_.Q ;
 wire \mem_right_track_6.DFFR_0_.Q ;
 wire \mem_right_track_6.DFFR_1_.Q ;
 wire \mem_right_track_6.DFFR_2_.Q ;
 wire \mem_right_track_6.DFFR_3_.Q ;
 wire \mem_right_track_6.DFFR_4_.Q ;
 wire \mem_right_track_6.DFFR_5_.Q ;
 wire \mem_right_track_8.DFFR_0_.Q ;
 wire \mem_top_track_0.DFFR_0_.Q ;
 wire \mem_top_track_0.DFFR_1_.Q ;
 wire \mem_top_track_0.DFFR_2_.Q ;
 wire \mem_top_track_0.DFFR_3_.Q ;
 wire \mem_top_track_0.DFFR_4_.Q ;
 wire \mem_top_track_0.DFFR_5_.Q ;
 wire \mem_top_track_0.DFFR_6_.Q ;
 wire \mem_top_track_0.DFFR_7_.Q ;
 wire \mem_top_track_16.DFFR_0_.D ;
 wire \mem_top_track_16.DFFR_0_.Q ;
 wire \mem_top_track_16.DFFR_1_.Q ;
 wire \mem_top_track_16.DFFR_2_.Q ;
 wire \mem_top_track_16.DFFR_3_.Q ;
 wire \mem_top_track_16.DFFR_4_.Q ;
 wire \mem_top_track_16.DFFR_5_.Q ;
 wire \mem_top_track_16.DFFR_6_.Q ;
 wire \mem_top_track_16.DFFR_7_.Q ;
 wire \mem_top_track_24.DFFR_0_.Q ;
 wire \mem_top_track_24.DFFR_1_.Q ;
 wire \mem_top_track_24.DFFR_2_.Q ;
 wire \mem_top_track_24.DFFR_3_.Q ;
 wire \mem_top_track_24.DFFR_4_.Q ;
 wire \mem_top_track_24.DFFR_5_.Q ;
 wire \mem_top_track_32.DFFR_0_.Q ;
 wire \mem_top_track_32.DFFR_1_.Q ;
 wire \mem_top_track_32.DFFR_2_.Q ;
 wire \mem_top_track_32.DFFR_3_.Q ;
 wire \mem_top_track_32.DFFR_4_.Q ;
 wire \mem_top_track_8.DFFR_0_.Q ;
 wire \mem_top_track_8.DFFR_1_.Q ;
 wire \mem_top_track_8.DFFR_2_.Q ;
 wire \mem_top_track_8.DFFR_3_.Q ;
 wire \mem_top_track_8.DFFR_4_.Q ;
 wire \mem_top_track_8.DFFR_5_.Q ;
 wire \mem_top_track_8.DFFR_6_.Q ;
 wire \mux_bottom_track_1.INVTX1_0_.out ;
 wire \mux_bottom_track_1.INVTX1_1_.out ;
 wire \mux_bottom_track_1.INVTX1_2_.out ;
 wire \mux_bottom_track_1.INVTX1_3_.out ;
 wire \mux_bottom_track_1.INVTX1_4_.out ;
 wire \mux_bottom_track_1.INVTX1_5_.out ;
 wire \mux_bottom_track_1.INVTX1_6_.out ;
 wire \mux_bottom_track_1.INVTX1_7_.out ;
 wire \mux_bottom_track_1.INVTX1_8_.out ;
 wire \mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out ;
 wire \mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out ;
 wire \mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out ;
 wire \mux_bottom_track_1.out ;
 wire \mux_bottom_track_17.INVTX1_0_.out ;
 wire \mux_bottom_track_17.INVTX1_1_.out ;
 wire \mux_bottom_track_17.INVTX1_2_.out ;
 wire \mux_bottom_track_17.INVTX1_3_.out ;
 wire \mux_bottom_track_17.INVTX1_4_.out ;
 wire \mux_bottom_track_17.INVTX1_5_.out ;
 wire \mux_bottom_track_17.INVTX1_6_.out ;
 wire \mux_bottom_track_17.INVTX1_7_.out ;
 wire \mux_bottom_track_17.INVTX1_8_.out ;
 wire \mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out ;
 wire \mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out ;
 wire \mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out ;
 wire \mux_bottom_track_17.out ;
 wire \mux_bottom_track_25.INVTX1_0_.out ;
 wire \mux_bottom_track_25.INVTX1_1_.out ;
 wire \mux_bottom_track_25.INVTX1_2_.out ;
 wire \mux_bottom_track_25.INVTX1_3_.out ;
 wire \mux_bottom_track_25.INVTX1_4_.out ;
 wire \mux_bottom_track_25.INVTX1_5_.out ;
 wire \mux_bottom_track_25.INVTX1_6_.out ;
 wire \mux_bottom_track_25.INVTX1_7_.out ;
 wire \mux_bottom_track_25.INVTX1_8_.out ;
 wire \mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out ;
 wire \mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out ;
 wire \mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out ;
 wire \mux_bottom_track_25.out ;
 wire \mux_bottom_track_33.INVTX1_0_.out ;
 wire \mux_bottom_track_33.INVTX1_1_.out ;
 wire \mux_bottom_track_33.INVTX1_2_.out ;
 wire \mux_bottom_track_33.INVTX1_3_.out ;
 wire \mux_bottom_track_33.INVTX1_4_.out ;
 wire \mux_bottom_track_33.INVTX1_5_.out ;
 wire \mux_bottom_track_33.INVTX1_6_.out ;
 wire \mux_bottom_track_33.mux_2level_tapbuf_basis_input2_mem2_0_out ;
 wire \mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_bottom_track_33.out ;
 wire \mux_bottom_track_9.INVTX1_0_.out ;
 wire \mux_bottom_track_9.INVTX1_1_.out ;
 wire \mux_bottom_track_9.INVTX1_2_.out ;
 wire \mux_bottom_track_9.INVTX1_3_.out ;
 wire \mux_bottom_track_9.INVTX1_4_.out ;
 wire \mux_bottom_track_9.INVTX1_5_.out ;
 wire \mux_bottom_track_9.INVTX1_6_.out ;
 wire \mux_bottom_track_9.INVTX1_7_.out ;
 wire \mux_bottom_track_9.INVTX1_8_.out ;
 wire \mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out ;
 wire \mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out ;
 wire \mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out ;
 wire \mux_bottom_track_9.out ;
 wire \mux_right_track_0.INVTX1_1_.out ;
 wire \mux_right_track_0.INVTX1_2_.out ;
 wire \mux_right_track_0.INVTX1_3_.out ;
 wire \mux_right_track_0.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_right_track_0.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_right_track_0.out ;
 wire \mux_right_track_10.INVTX1_1_.out ;
 wire \mux_right_track_10.INVTX1_2_.out ;
 wire \mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_right_track_10.out ;
 wire \mux_right_track_12.INVTX1_1_.out ;
 wire \mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_right_track_12.out ;
 wire \mux_right_track_14.INVTX1_1_.out ;
 wire \mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_right_track_14.out ;
 wire \mux_right_track_16.INVTX1_1_.out ;
 wire \mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_right_track_16.out ;
 wire \mux_right_track_18.INVTX1_2_.out ;
 wire \mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_right_track_18.out ;
 wire \mux_right_track_2.INVTX1_1_.out ;
 wire \mux_right_track_2.INVTX1_3_.out ;
 wire \mux_right_track_2.INVTX1_4_.out ;
 wire \mux_right_track_2.mux_2level_tapbuf_basis_input2_mem2_0_out ;
 wire \mux_right_track_2.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_right_track_2.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_right_track_2.out ;
 wire \mux_right_track_20.INVTX1_2_.out ;
 wire \mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_right_track_20.out ;
 wire \mux_right_track_22.INVTX1_2_.out ;
 wire \mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_right_track_22.out ;
 wire \mux_right_track_24.INVTX1_1_.out ;
 wire \mux_right_track_24.INVTX1_2_.out ;
 wire \mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_right_track_24.out ;
 wire \mux_right_track_26.INVTX1_1_.out ;
 wire \mux_right_track_26.INVTX1_2_.out ;
 wire \mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_right_track_26.out ;
 wire \mux_right_track_4.INVTX1_1_.out ;
 wire \mux_right_track_4.INVTX1_4_.out ;
 wire \mux_right_track_4.mux_2level_tapbuf_basis_input2_mem2_0_out ;
 wire \mux_right_track_4.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_right_track_4.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_right_track_4.out ;
 wire \mux_right_track_6.INVTX1_1_.out ;
 wire \mux_right_track_6.INVTX1_3_.out ;
 wire \mux_right_track_6.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_right_track_6.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_right_track_6.out ;
 wire \mux_right_track_8.INVTX1_1_.out ;
 wire \mux_right_track_8.INVTX1_2_.out ;
 wire \mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_right_track_8.out ;
 wire \mux_top_track_0.INVTX1_0_.out ;
 wire \mux_top_track_0.INVTX1_1_.out ;
 wire \mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out ;
 wire \mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out ;
 wire \mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out ;
 wire \mux_top_track_0.out ;
 wire \mux_top_track_16.INVTX1_0_.out ;
 wire \mux_top_track_16.INVTX1_1_.out ;
 wire \mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out ;
 wire \mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out ;
 wire \mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out ;
 wire \mux_top_track_16.out ;
 wire \mux_top_track_24.INVTX1_0_.out ;
 wire \mux_top_track_24.INVTX1_1_.out ;
 wire \mux_top_track_24.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_top_track_24.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_top_track_24.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_top_track_24.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_top_track_24.out ;
 wire \mux_top_track_32.INVTX1_0_.out ;
 wire \mux_top_track_32.INVTX1_1_.out ;
 wire \mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_top_track_32.out ;
 wire \mux_top_track_8.INVTX1_0_.out ;
 wire \mux_top_track_8.INVTX1_1_.out ;
 wire \mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out ;
 wire \mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out ;
 wire \mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out ;
 wire \mux_top_track_8.out ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire clknet_4_0_0_prog_clk;
 wire clknet_4_1_0_prog_clk;
 wire clknet_4_2_0_prog_clk;
 wire clknet_4_3_0_prog_clk;
 wire clknet_4_4_0_prog_clk;
 wire clknet_4_5_0_prog_clk;
 wire clknet_4_6_0_prog_clk;
 wire clknet_4_7_0_prog_clk;
 wire clknet_4_8_0_prog_clk;
 wire clknet_4_9_0_prog_clk;
 wire clknet_4_10_0_prog_clk;
 wire clknet_4_11_0_prog_clk;
 wire clknet_4_12_0_prog_clk;
 wire clknet_4_13_0_prog_clk;
 wire clknet_4_14_0_prog_clk;
 wire clknet_4_15_0_prog_clk;

 sky130_fd_sc_hd__inv_2 _0383_ (.A(\mem_top_track_0.DFFR_5_.Q ),
    .Y(_0158_));
 sky130_fd_sc_hd__inv_2 _0384_ (.A(\mem_bottom_track_33.DFFR_3_.Q ),
    .Y(_0356_));
 sky130_fd_sc_hd__inv_2 _0385_ (.A(\mem_bottom_track_33.DFFR_0_.Q ),
    .Y(_0358_));
 sky130_fd_sc_hd__inv_2 _0386_ (.A(\mem_bottom_track_33.DFFR_2_.Q ),
    .Y(_0354_));
 sky130_fd_sc_hd__inv_2 _0387_ (.A(\mem_bottom_track_33.DFFR_1_.Q ),
    .Y(_0353_));
 sky130_fd_sc_hd__inv_2 _0388_ (.A(net84),
    .Y(_0350_));
 sky130_fd_sc_hd__inv_2 _0389_ (.A(\mem_bottom_track_33.DFFR_0_.Q ),
    .Y(_0355_));
 sky130_fd_sc_hd__inv_2 _0390_ (.A(\mem_bottom_track_33.DFFR_4_.Q ),
    .Y(_0349_));
 sky130_fd_sc_hd__inv_2 _0391_ (.A(\mem_bottom_track_33.DFFR_0_.Q ),
    .Y(_0357_));
 sky130_fd_sc_hd__inv_2 _0392_ (.A(\mem_bottom_track_33.DFFR_2_.Q ),
    .Y(_0352_));
 sky130_fd_sc_hd__inv_2 _0393_ (.A(\mem_bottom_track_33.DFFR_1_.Q ),
    .Y(_0351_));
 sky130_fd_sc_hd__inv_2 _0394_ (.A(\mem_bottom_track_33.DFFR_1_.Q ),
    .Y(_0348_));
 sky130_fd_sc_hd__inv_2 _0395_ (.A(\mem_right_track_16.DFFR_1_.Q ),
    .Y(_0346_));
 sky130_fd_sc_hd__inv_2 _0396_ (.A(\mem_right_track_16.DFFR_0_.Q ),
    .Y(_0347_));
 sky130_fd_sc_hd__clkbuf_1 _0397_ (.A(\mem_right_track_16.DFFR_0_.Q ),
    .X(_0126_));
 sky130_fd_sc_hd__clkbuf_1 _0398_ (.A(_0126_),
    .X(_0345_));
 sky130_fd_sc_hd__clkbuf_1 _0399_ (.A(\mem_right_track_16.DFFR_1_.Q ),
    .X(_0127_));
 sky130_fd_sc_hd__clkbuf_1 _0400_ (.A(_0127_),
    .X(_0344_));
 sky130_fd_sc_hd__inv_2 _0401_ (.A(\mem_right_track_14.DFFR_1_.Q ),
    .Y(_0342_));
 sky130_fd_sc_hd__inv_2 _0402_ (.A(\mem_right_track_14.DFFR_0_.Q ),
    .Y(_0343_));
 sky130_fd_sc_hd__clkbuf_1 _0403_ (.A(\mem_right_track_14.DFFR_0_.Q ),
    .X(_0128_));
 sky130_fd_sc_hd__clkbuf_1 _0404_ (.A(_0128_),
    .X(_0341_));
 sky130_fd_sc_hd__clkbuf_1 _0405_ (.A(\mem_right_track_14.DFFR_1_.Q ),
    .X(_0129_));
 sky130_fd_sc_hd__clkbuf_1 _0406_ (.A(_0129_),
    .X(_0340_));
 sky130_fd_sc_hd__inv_2 _0407_ (.A(\mem_right_track_12.DFFR_1_.Q ),
    .Y(_0338_));
 sky130_fd_sc_hd__inv_2 _0408_ (.A(\mem_right_track_12.DFFR_0_.Q ),
    .Y(_0339_));
 sky130_fd_sc_hd__clkbuf_1 _0409_ (.A(\mem_right_track_12.DFFR_0_.Q ),
    .X(_0130_));
 sky130_fd_sc_hd__clkbuf_1 _0410_ (.A(_0130_),
    .X(_0337_));
 sky130_fd_sc_hd__clkbuf_1 _0411_ (.A(\mem_right_track_12.DFFR_1_.Q ),
    .X(_0131_));
 sky130_fd_sc_hd__clkbuf_1 _0412_ (.A(_0131_),
    .X(_0336_));
 sky130_fd_sc_hd__inv_2 _0413_ (.A(\mem_bottom_track_1.DFFR_0_.D ),
    .Y(_0333_));
 sky130_fd_sc_hd__inv_2 _0414_ (.A(\mem_right_track_26.DFFR_0_.Q ),
    .Y(_0335_));
 sky130_fd_sc_hd__clkbuf_1 _0415_ (.A(\mem_right_track_26.DFFR_0_.Q ),
    .X(_0132_));
 sky130_fd_sc_hd__clkbuf_1 _0416_ (.A(_0132_),
    .X(_0332_));
 sky130_fd_sc_hd__clkbuf_1 _0417_ (.A(\mem_bottom_track_1.DFFR_0_.D ),
    .X(_0133_));
 sky130_fd_sc_hd__clkbuf_1 _0418_ (.A(_0133_),
    .X(_0330_));
 sky130_fd_sc_hd__inv_2 _0419_ (.A(\mem_right_track_26.DFFR_0_.Q ),
    .Y(_0334_));
 sky130_fd_sc_hd__clkbuf_1 _0420_ (.A(\mem_right_track_26.DFFR_0_.Q ),
    .X(_0134_));
 sky130_fd_sc_hd__clkbuf_1 _0421_ (.A(_0134_),
    .X(_0331_));
 sky130_fd_sc_hd__inv_2 _0422_ (.A(\mem_right_track_24.DFFR_1_.Q ),
    .Y(_0327_));
 sky130_fd_sc_hd__inv_2 _0423_ (.A(\mem_right_track_24.DFFR_0_.Q ),
    .Y(_0329_));
 sky130_fd_sc_hd__clkbuf_1 _0424_ (.A(\mem_right_track_24.DFFR_0_.Q ),
    .X(_0135_));
 sky130_fd_sc_hd__clkbuf_1 _0425_ (.A(_0135_),
    .X(_0326_));
 sky130_fd_sc_hd__clkbuf_1 _0426_ (.A(\mem_right_track_24.DFFR_1_.Q ),
    .X(_0136_));
 sky130_fd_sc_hd__clkbuf_1 _0427_ (.A(_0136_),
    .X(_0324_));
 sky130_fd_sc_hd__inv_2 _0428_ (.A(\mem_right_track_24.DFFR_0_.Q ),
    .Y(_0328_));
 sky130_fd_sc_hd__clkbuf_1 _0429_ (.A(\mem_right_track_24.DFFR_0_.Q ),
    .X(_0137_));
 sky130_fd_sc_hd__clkbuf_1 _0430_ (.A(_0137_),
    .X(_0325_));
 sky130_fd_sc_hd__inv_2 _0431_ (.A(\mem_right_track_22.DFFR_1_.Q ),
    .Y(_0321_));
 sky130_fd_sc_hd__inv_2 _0432_ (.A(\mem_right_track_22.DFFR_0_.Q ),
    .Y(_0323_));
 sky130_fd_sc_hd__clkbuf_1 _0433_ (.A(\mem_right_track_22.DFFR_0_.Q ),
    .X(_0138_));
 sky130_fd_sc_hd__clkbuf_1 _0434_ (.A(_0138_),
    .X(_0320_));
 sky130_fd_sc_hd__clkbuf_1 _0435_ (.A(\mem_right_track_22.DFFR_1_.Q ),
    .X(_0139_));
 sky130_fd_sc_hd__clkbuf_1 _0436_ (.A(_0139_),
    .X(_0318_));
 sky130_fd_sc_hd__inv_2 _0437_ (.A(\mem_right_track_22.DFFR_0_.Q ),
    .Y(_0322_));
 sky130_fd_sc_hd__clkbuf_1 _0438_ (.A(\mem_right_track_22.DFFR_0_.Q ),
    .X(_0140_));
 sky130_fd_sc_hd__clkbuf_1 _0439_ (.A(_0140_),
    .X(_0319_));
 sky130_fd_sc_hd__inv_2 _0440_ (.A(\mem_right_track_20.DFFR_1_.Q ),
    .Y(_0315_));
 sky130_fd_sc_hd__inv_2 _0441_ (.A(\mem_right_track_20.DFFR_0_.Q ),
    .Y(_0317_));
 sky130_fd_sc_hd__clkbuf_1 _0442_ (.A(\mem_right_track_20.DFFR_0_.Q ),
    .X(_0141_));
 sky130_fd_sc_hd__clkbuf_1 _0443_ (.A(_0141_),
    .X(_0314_));
 sky130_fd_sc_hd__clkbuf_1 _0444_ (.A(\mem_right_track_20.DFFR_1_.Q ),
    .X(_0142_));
 sky130_fd_sc_hd__clkbuf_1 _0445_ (.A(_0142_),
    .X(_0312_));
 sky130_fd_sc_hd__inv_2 _0446_ (.A(\mem_right_track_20.DFFR_0_.Q ),
    .Y(_0316_));
 sky130_fd_sc_hd__clkbuf_1 _0447_ (.A(\mem_right_track_20.DFFR_0_.Q ),
    .X(_0143_));
 sky130_fd_sc_hd__clkbuf_1 _0448_ (.A(_0143_),
    .X(_0313_));
 sky130_fd_sc_hd__inv_2 _0449_ (.A(\mem_right_track_18.DFFR_1_.Q ),
    .Y(_0309_));
 sky130_fd_sc_hd__inv_2 _0450_ (.A(\mem_right_track_18.DFFR_0_.Q ),
    .Y(_0311_));
 sky130_fd_sc_hd__clkbuf_1 _0451_ (.A(\mem_right_track_18.DFFR_0_.Q ),
    .X(_0144_));
 sky130_fd_sc_hd__clkbuf_1 _0452_ (.A(_0144_),
    .X(_0308_));
 sky130_fd_sc_hd__clkbuf_1 _0453_ (.A(\mem_right_track_18.DFFR_1_.Q ),
    .X(_0145_));
 sky130_fd_sc_hd__clkbuf_1 _0454_ (.A(_0145_),
    .X(_0306_));
 sky130_fd_sc_hd__inv_2 _0455_ (.A(\mem_right_track_18.DFFR_0_.Q ),
    .Y(_0310_));
 sky130_fd_sc_hd__clkbuf_1 _0456_ (.A(\mem_right_track_18.DFFR_0_.Q ),
    .X(_0146_));
 sky130_fd_sc_hd__clkbuf_1 _0457_ (.A(_0146_),
    .X(_0307_));
 sky130_fd_sc_hd__inv_2 _0458_ (.A(\mem_right_track_10.DFFR_1_.Q ),
    .Y(_0303_));
 sky130_fd_sc_hd__inv_2 _0459_ (.A(\mem_right_track_10.DFFR_0_.Q ),
    .Y(_0305_));
 sky130_fd_sc_hd__clkbuf_1 _0460_ (.A(\mem_right_track_10.DFFR_0_.Q ),
    .X(_0147_));
 sky130_fd_sc_hd__clkbuf_1 _0461_ (.A(_0147_),
    .X(_0302_));
 sky130_fd_sc_hd__clkbuf_1 _0462_ (.A(\mem_right_track_10.DFFR_1_.Q ),
    .X(_0148_));
 sky130_fd_sc_hd__clkbuf_1 _0463_ (.A(_0148_),
    .X(_0300_));
 sky130_fd_sc_hd__inv_2 _0464_ (.A(\mem_right_track_10.DFFR_0_.Q ),
    .Y(_0304_));
 sky130_fd_sc_hd__clkbuf_1 _0465_ (.A(\mem_right_track_10.DFFR_0_.Q ),
    .X(_0149_));
 sky130_fd_sc_hd__clkbuf_1 _0466_ (.A(_0149_),
    .X(_0301_));
 sky130_fd_sc_hd__inv_2 _0467_ (.A(\mem_right_track_10.DFFR_0_.D ),
    .Y(_0297_));
 sky130_fd_sc_hd__inv_2 _0468_ (.A(\mem_right_track_8.DFFR_0_.Q ),
    .Y(_0299_));
 sky130_fd_sc_hd__clkbuf_1 _0469_ (.A(\mem_right_track_8.DFFR_0_.Q ),
    .X(_0150_));
 sky130_fd_sc_hd__clkbuf_1 _0470_ (.A(_0150_),
    .X(_0296_));
 sky130_fd_sc_hd__clkbuf_1 _0471_ (.A(\mem_right_track_10.DFFR_0_.D ),
    .X(_0151_));
 sky130_fd_sc_hd__clkbuf_1 _0472_ (.A(_0151_),
    .X(_0294_));
 sky130_fd_sc_hd__inv_2 _0473_ (.A(\mem_right_track_8.DFFR_0_.Q ),
    .Y(_0298_));
 sky130_fd_sc_hd__clkbuf_1 _0474_ (.A(\mem_right_track_8.DFFR_0_.Q ),
    .X(_0152_));
 sky130_fd_sc_hd__clkbuf_1 _0475_ (.A(_0152_),
    .X(_0295_));
 sky130_fd_sc_hd__inv_2 _0476_ (.A(\mem_right_track_4.DFFR_3_.Q ),
    .Y(_0292_));
 sky130_fd_sc_hd__inv_2 _0477_ (.A(\mem_right_track_4.DFFR_0_.Q ),
    .Y(_0293_));
 sky130_fd_sc_hd__inv_2 _0478_ (.A(\mem_right_track_4.DFFR_2_.Q ),
    .Y(_0290_));
 sky130_fd_sc_hd__inv_2 _0479_ (.A(\mem_right_track_4.DFFR_1_.Q ),
    .Y(_0289_));
 sky130_fd_sc_hd__inv_2 _0480_ (.A(\mem_right_track_4.DFFR_5_.Q ),
    .Y(_0288_));
 sky130_fd_sc_hd__inv_2 _0481_ (.A(\mem_right_track_4.DFFR_4_.Q ),
    .Y(_0287_));
 sky130_fd_sc_hd__inv_2 _0482_ (.A(\mem_right_track_4.DFFR_0_.Q ),
    .Y(_0291_));
 sky130_fd_sc_hd__inv_2 _0483_ (.A(\mem_right_track_4.DFFR_1_.Q ),
    .Y(_0286_));
 sky130_fd_sc_hd__inv_2 _0484_ (.A(\mem_right_track_2.DFFR_3_.Q ),
    .Y(_0284_));
 sky130_fd_sc_hd__inv_2 _0485_ (.A(\mem_right_track_2.DFFR_0_.Q ),
    .Y(_0285_));
 sky130_fd_sc_hd__inv_2 _0486_ (.A(\mem_right_track_2.DFFR_2_.Q ),
    .Y(_0282_));
 sky130_fd_sc_hd__inv_2 _0487_ (.A(\mem_right_track_2.DFFR_1_.Q ),
    .Y(_0281_));
 sky130_fd_sc_hd__inv_2 _0488_ (.A(\mem_right_track_2.DFFR_5_.Q ),
    .Y(_0280_));
 sky130_fd_sc_hd__inv_2 _0489_ (.A(\mem_right_track_2.DFFR_4_.Q ),
    .Y(_0279_));
 sky130_fd_sc_hd__inv_2 _0490_ (.A(\mem_right_track_2.DFFR_0_.Q ),
    .Y(_0283_));
 sky130_fd_sc_hd__inv_2 _0491_ (.A(\mem_right_track_2.DFFR_1_.Q ),
    .Y(_0278_));
 sky130_fd_sc_hd__inv_2 _0492_ (.A(\mem_right_track_6.DFFR_3_.Q ),
    .Y(_0276_));
 sky130_fd_sc_hd__inv_2 _0493_ (.A(\mem_right_track_6.DFFR_0_.Q ),
    .Y(_0277_));
 sky130_fd_sc_hd__inv_2 _0494_ (.A(\mem_right_track_6.DFFR_2_.Q ),
    .Y(_0275_));
 sky130_fd_sc_hd__inv_2 _0495_ (.A(\mem_right_track_6.DFFR_1_.Q ),
    .Y(_0274_));
 sky130_fd_sc_hd__inv_2 _0496_ (.A(\mem_right_track_6.DFFR_5_.Q ),
    .Y(_0273_));
 sky130_fd_sc_hd__inv_2 _0497_ (.A(\mem_right_track_6.DFFR_4_.Q ),
    .Y(_0272_));
 sky130_fd_sc_hd__inv_2 _0498_ (.A(\mem_right_track_0.DFFR_3_.Q ),
    .Y(_0270_));
 sky130_fd_sc_hd__inv_2 _0499_ (.A(\mem_right_track_0.DFFR_0_.Q ),
    .Y(_0271_));
 sky130_fd_sc_hd__inv_2 _0500_ (.A(\mem_right_track_0.DFFR_2_.Q ),
    .Y(_0269_));
 sky130_fd_sc_hd__inv_2 _0501_ (.A(\mem_right_track_0.DFFR_1_.Q ),
    .Y(_0268_));
 sky130_fd_sc_hd__inv_2 _0502_ (.A(\mem_right_track_0.DFFR_5_.Q ),
    .Y(_0267_));
 sky130_fd_sc_hd__inv_2 _0503_ (.A(\mem_right_track_0.DFFR_4_.Q ),
    .Y(_0266_));
 sky130_fd_sc_hd__inv_2 _0504_ (.A(\mem_top_track_32.DFFR_3_.Q ),
    .Y(_0262_));
 sky130_fd_sc_hd__inv_2 _0505_ (.A(\mem_top_track_32.DFFR_0_.Q ),
    .Y(_0265_));
 sky130_fd_sc_hd__inv_2 _0506_ (.A(\mem_top_track_32.DFFR_2_.Q ),
    .Y(_0261_));
 sky130_fd_sc_hd__inv_2 _0507_ (.A(\mem_top_track_32.DFFR_1_.Q ),
    .Y(_0260_));
 sky130_fd_sc_hd__inv_2 _0508_ (.A(\mem_right_track_0.DFFR_0_.D ),
    .Y(_0255_));
 sky130_fd_sc_hd__inv_2 _0509_ (.A(\mem_top_track_32.DFFR_0_.Q ),
    .Y(_0263_));
 sky130_fd_sc_hd__inv_2 _0510_ (.A(\mem_top_track_32.DFFR_2_.Q ),
    .Y(_0257_));
 sky130_fd_sc_hd__inv_2 _0511_ (.A(\mem_top_track_32.DFFR_1_.Q ),
    .Y(_0256_));
 sky130_fd_sc_hd__inv_2 _0512_ (.A(\mem_top_track_32.DFFR_4_.Q ),
    .Y(_0254_));
 sky130_fd_sc_hd__inv_2 _0513_ (.A(\mem_top_track_32.DFFR_0_.Q ),
    .Y(_0264_));
 sky130_fd_sc_hd__inv_2 _0514_ (.A(\mem_top_track_32.DFFR_2_.Q ),
    .Y(_0259_));
 sky130_fd_sc_hd__inv_2 _0515_ (.A(\mem_top_track_32.DFFR_1_.Q ),
    .Y(_0258_));
 sky130_fd_sc_hd__inv_2 _0516_ (.A(\mem_top_track_24.DFFR_3_.Q ),
    .Y(_0250_));
 sky130_fd_sc_hd__inv_2 _0517_ (.A(\mem_top_track_24.DFFR_0_.Q ),
    .Y(_0253_));
 sky130_fd_sc_hd__inv_2 _0518_ (.A(\mem_top_track_24.DFFR_2_.Q ),
    .Y(_0249_));
 sky130_fd_sc_hd__inv_2 _0519_ (.A(\mem_top_track_24.DFFR_1_.Q ),
    .Y(_0248_));
 sky130_fd_sc_hd__inv_2 _0520_ (.A(\mem_top_track_24.DFFR_5_.Q ),
    .Y(_0243_));
 sky130_fd_sc_hd__inv_2 _0521_ (.A(\mem_top_track_24.DFFR_0_.Q ),
    .Y(_0251_));
 sky130_fd_sc_hd__inv_2 _0522_ (.A(\mem_top_track_24.DFFR_2_.Q ),
    .Y(_0245_));
 sky130_fd_sc_hd__inv_2 _0523_ (.A(\mem_top_track_24.DFFR_1_.Q ),
    .Y(_0244_));
 sky130_fd_sc_hd__inv_2 _0524_ (.A(\mem_top_track_24.DFFR_4_.Q ),
    .Y(_0242_));
 sky130_fd_sc_hd__inv_2 _0525_ (.A(\mem_top_track_24.DFFR_0_.Q ),
    .Y(_0252_));
 sky130_fd_sc_hd__inv_2 _0526_ (.A(\mem_top_track_24.DFFR_2_.Q ),
    .Y(_0247_));
 sky130_fd_sc_hd__inv_2 _0527_ (.A(\mem_top_track_24.DFFR_1_.Q ),
    .Y(_0246_));
 sky130_fd_sc_hd__inv_2 _0528_ (.A(\mem_bottom_track_25.DFFR_4_.Q ),
    .Y(_0239_));
 sky130_fd_sc_hd__inv_2 _0529_ (.A(\mem_bottom_track_25.DFFR_0_.Q ),
    .Y(_0241_));
 sky130_fd_sc_hd__inv_2 _0530_ (.A(\mem_bottom_track_25.DFFR_3_.Q ),
    .Y(_0238_));
 sky130_fd_sc_hd__inv_2 _0531_ (.A(\mem_bottom_track_25.DFFR_2_.Q ),
    .Y(_0237_));
 sky130_fd_sc_hd__inv_2 _0532_ (.A(\mem_bottom_track_25.DFFR_1_.Q ),
    .Y(_0236_));
 sky130_fd_sc_hd__inv_2 _0533_ (.A(\mem_bottom_track_25.DFFR_7_.Q ),
    .Y(_0232_));
 sky130_fd_sc_hd__inv_2 _0534_ (.A(\mem_bottom_track_25.DFFR_6_.Q ),
    .Y(_0231_));
 sky130_fd_sc_hd__inv_2 _0535_ (.A(\mem_bottom_track_25.DFFR_5_.Q ),
    .Y(_0230_));
 sky130_fd_sc_hd__inv_2 _0536_ (.A(\mem_bottom_track_25.DFFR_0_.Q ),
    .Y(_0240_));
 sky130_fd_sc_hd__inv_2 _0537_ (.A(\mem_bottom_track_25.DFFR_3_.Q ),
    .Y(_0235_));
 sky130_fd_sc_hd__inv_2 _0538_ (.A(\mem_bottom_track_25.DFFR_2_.Q ),
    .Y(_0234_));
 sky130_fd_sc_hd__inv_2 _0539_ (.A(\mem_bottom_track_25.DFFR_1_.Q ),
    .Y(_0233_));
 sky130_fd_sc_hd__inv_2 _0540_ (.A(\mem_bottom_track_17.DFFR_4_.Q ),
    .Y(_0227_));
 sky130_fd_sc_hd__inv_2 _0541_ (.A(\mem_bottom_track_17.DFFR_0_.Q ),
    .Y(_0229_));
 sky130_fd_sc_hd__inv_2 _0542_ (.A(\mem_bottom_track_17.DFFR_3_.Q ),
    .Y(_0226_));
 sky130_fd_sc_hd__inv_2 _0543_ (.A(\mem_bottom_track_17.DFFR_2_.Q ),
    .Y(_0225_));
 sky130_fd_sc_hd__inv_2 _0544_ (.A(\mem_bottom_track_17.DFFR_1_.Q ),
    .Y(_0224_));
 sky130_fd_sc_hd__inv_2 _0545_ (.A(\mem_bottom_track_17.DFFR_7_.Q ),
    .Y(_0220_));
 sky130_fd_sc_hd__inv_2 _0546_ (.A(\mem_bottom_track_17.DFFR_6_.Q ),
    .Y(_0219_));
 sky130_fd_sc_hd__inv_2 _0547_ (.A(\mem_bottom_track_17.DFFR_5_.Q ),
    .Y(_0218_));
 sky130_fd_sc_hd__inv_2 _0548_ (.A(\mem_bottom_track_17.DFFR_0_.Q ),
    .Y(_0228_));
 sky130_fd_sc_hd__inv_2 _0549_ (.A(\mem_bottom_track_17.DFFR_3_.Q ),
    .Y(_0223_));
 sky130_fd_sc_hd__inv_2 _0550_ (.A(\mem_bottom_track_17.DFFR_2_.Q ),
    .Y(_0222_));
 sky130_fd_sc_hd__inv_2 _0551_ (.A(\mem_bottom_track_17.DFFR_1_.Q ),
    .Y(_0221_));
 sky130_fd_sc_hd__inv_2 _0552_ (.A(\mem_bottom_track_9.DFFR_4_.Q ),
    .Y(_0215_));
 sky130_fd_sc_hd__inv_2 _0553_ (.A(\mem_bottom_track_9.DFFR_0_.Q ),
    .Y(_0217_));
 sky130_fd_sc_hd__inv_2 _0554_ (.A(\mem_bottom_track_9.DFFR_3_.Q ),
    .Y(_0214_));
 sky130_fd_sc_hd__inv_2 _0555_ (.A(\mem_bottom_track_9.DFFR_2_.Q ),
    .Y(_0213_));
 sky130_fd_sc_hd__inv_2 _0556_ (.A(\mem_bottom_track_9.DFFR_1_.Q ),
    .Y(_0212_));
 sky130_fd_sc_hd__inv_2 _0557_ (.A(\mem_bottom_track_17.DFFR_0_.D ),
    .Y(_0208_));
 sky130_fd_sc_hd__inv_2 _0558_ (.A(\mem_bottom_track_9.DFFR_6_.Q ),
    .Y(_0207_));
 sky130_fd_sc_hd__inv_2 _0559_ (.A(\mem_bottom_track_9.DFFR_5_.Q ),
    .Y(_0206_));
 sky130_fd_sc_hd__inv_2 _0560_ (.A(\mem_bottom_track_9.DFFR_0_.Q ),
    .Y(_0216_));
 sky130_fd_sc_hd__inv_2 _0561_ (.A(\mem_bottom_track_9.DFFR_3_.Q ),
    .Y(_0211_));
 sky130_fd_sc_hd__inv_2 _0562_ (.A(\mem_bottom_track_9.DFFR_2_.Q ),
    .Y(_0210_));
 sky130_fd_sc_hd__inv_2 _0563_ (.A(\mem_bottom_track_9.DFFR_1_.Q ),
    .Y(_0209_));
 sky130_fd_sc_hd__inv_2 _0564_ (.A(\mem_bottom_track_1.DFFR_4_.Q ),
    .Y(_0203_));
 sky130_fd_sc_hd__inv_2 _0565_ (.A(\mem_bottom_track_1.DFFR_0_.Q ),
    .Y(_0205_));
 sky130_fd_sc_hd__inv_2 _0566_ (.A(\mem_bottom_track_1.DFFR_3_.Q ),
    .Y(_0202_));
 sky130_fd_sc_hd__inv_2 _0567_ (.A(\mem_bottom_track_1.DFFR_2_.Q ),
    .Y(_0201_));
 sky130_fd_sc_hd__inv_2 _0568_ (.A(\mem_bottom_track_1.DFFR_1_.Q ),
    .Y(_0200_));
 sky130_fd_sc_hd__inv_2 _0569_ (.A(\mem_bottom_track_1.DFFR_7_.Q ),
    .Y(_0196_));
 sky130_fd_sc_hd__inv_2 _0570_ (.A(\mem_bottom_track_1.DFFR_6_.Q ),
    .Y(_0195_));
 sky130_fd_sc_hd__inv_2 _0571_ (.A(\mem_bottom_track_1.DFFR_5_.Q ),
    .Y(_0194_));
 sky130_fd_sc_hd__inv_2 _0572_ (.A(\mem_bottom_track_1.DFFR_0_.Q ),
    .Y(_0204_));
 sky130_fd_sc_hd__inv_2 _0573_ (.A(\mem_bottom_track_1.DFFR_3_.Q ),
    .Y(_0199_));
 sky130_fd_sc_hd__inv_2 _0574_ (.A(\mem_bottom_track_1.DFFR_2_.Q ),
    .Y(_0198_));
 sky130_fd_sc_hd__inv_2 _0575_ (.A(\mem_bottom_track_1.DFFR_1_.Q ),
    .Y(_0197_));
 sky130_fd_sc_hd__inv_2 _0576_ (.A(\mem_top_track_16.DFFR_4_.Q ),
    .Y(_0191_));
 sky130_fd_sc_hd__inv_2 _0577_ (.A(\mem_top_track_16.DFFR_0_.Q ),
    .Y(_0193_));
 sky130_fd_sc_hd__inv_2 _0578_ (.A(\mem_top_track_16.DFFR_3_.Q ),
    .Y(_0190_));
 sky130_fd_sc_hd__inv_2 _0579_ (.A(\mem_top_track_16.DFFR_2_.Q ),
    .Y(_0189_));
 sky130_fd_sc_hd__inv_2 _0580_ (.A(\mem_top_track_16.DFFR_1_.Q ),
    .Y(_0188_));
 sky130_fd_sc_hd__inv_2 _0581_ (.A(\mem_top_track_16.DFFR_7_.Q ),
    .Y(_0184_));
 sky130_fd_sc_hd__inv_2 _0582_ (.A(\mem_top_track_16.DFFR_6_.Q ),
    .Y(_0183_));
 sky130_fd_sc_hd__inv_2 _0583_ (.A(\mem_top_track_16.DFFR_5_.Q ),
    .Y(_0182_));
 sky130_fd_sc_hd__inv_2 _0584_ (.A(\mem_top_track_16.DFFR_0_.Q ),
    .Y(_0192_));
 sky130_fd_sc_hd__inv_2 _0585_ (.A(\mem_top_track_16.DFFR_3_.Q ),
    .Y(_0187_));
 sky130_fd_sc_hd__inv_2 _0586_ (.A(\mem_top_track_16.DFFR_2_.Q ),
    .Y(_0186_));
 sky130_fd_sc_hd__inv_2 _0587_ (.A(\mem_top_track_16.DFFR_1_.Q ),
    .Y(_0185_));
 sky130_fd_sc_hd__inv_2 _0588_ (.A(\mem_top_track_8.DFFR_4_.Q ),
    .Y(_0179_));
 sky130_fd_sc_hd__inv_2 _0589_ (.A(\mem_top_track_8.DFFR_0_.Q ),
    .Y(_0181_));
 sky130_fd_sc_hd__inv_2 _0590_ (.A(\mem_top_track_8.DFFR_3_.Q ),
    .Y(_0178_));
 sky130_fd_sc_hd__inv_2 _0591_ (.A(\mem_top_track_8.DFFR_2_.Q ),
    .Y(_0177_));
 sky130_fd_sc_hd__inv_2 _0592_ (.A(\mem_top_track_8.DFFR_1_.Q ),
    .Y(_0176_));
 sky130_fd_sc_hd__inv_2 _0593_ (.A(\mem_top_track_16.DFFR_0_.D ),
    .Y(_0172_));
 sky130_fd_sc_hd__inv_2 _0594_ (.A(\mem_top_track_8.DFFR_6_.Q ),
    .Y(_0171_));
 sky130_fd_sc_hd__inv_2 _0595_ (.A(\mem_top_track_8.DFFR_5_.Q ),
    .Y(_0170_));
 sky130_fd_sc_hd__inv_2 _0596_ (.A(\mem_top_track_8.DFFR_0_.Q ),
    .Y(_0180_));
 sky130_fd_sc_hd__inv_2 _0597_ (.A(\mem_top_track_8.DFFR_3_.Q ),
    .Y(_0175_));
 sky130_fd_sc_hd__inv_2 _0598_ (.A(\mem_top_track_8.DFFR_2_.Q ),
    .Y(_0174_));
 sky130_fd_sc_hd__inv_2 _0599_ (.A(\mem_top_track_8.DFFR_1_.Q ),
    .Y(_0173_));
 sky130_fd_sc_hd__inv_2 _0600_ (.A(\mem_top_track_0.DFFR_0_.Q ),
    .Y(_0168_));
 sky130_fd_sc_hd__inv_2 _0601_ (.A(\mem_top_track_0.DFFR_4_.Q ),
    .Y(_0167_));
 sky130_fd_sc_hd__inv_2 _0602_ (.A(\mem_top_track_0.DFFR_0_.Q ),
    .Y(_0169_));
 sky130_fd_sc_hd__inv_2 _0603_ (.A(\mem_top_track_0.DFFR_3_.Q ),
    .Y(_0166_));
 sky130_fd_sc_hd__inv_2 _0604_ (.A(\mem_top_track_0.DFFR_2_.Q ),
    .Y(_0165_));
 sky130_fd_sc_hd__inv_2 _0605_ (.A(\mem_top_track_0.DFFR_1_.Q ),
    .Y(_0164_));
 sky130_fd_sc_hd__inv_2 _0606_ (.A(\mem_top_track_0.DFFR_3_.Q ),
    .Y(_0163_));
 sky130_fd_sc_hd__inv_2 _0607_ (.A(\mem_top_track_0.DFFR_2_.Q ),
    .Y(_0162_));
 sky130_fd_sc_hd__inv_2 _0608_ (.A(\mem_top_track_0.DFFR_1_.Q ),
    .Y(_0161_));
 sky130_fd_sc_hd__inv_2 _0609_ (.A(\mem_top_track_0.DFFR_7_.Q ),
    .Y(_0160_));
 sky130_fd_sc_hd__inv_2 _0610_ (.A(\mem_top_track_0.DFFR_6_.Q ),
    .Y(_0159_));
 sky130_fd_sc_hd__inv_2 _0611_ (.A(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out ),
    .Y(\mux_top_track_0.out ));
 sky130_fd_sc_hd__inv_2 _0612_ (.A(net79),
    .Y(\mux_top_track_0.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0613_ (.A(net74),
    .Y(\mux_top_track_0.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0614_ (.A(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out ),
    .Y(\mux_top_track_8.out ));
 sky130_fd_sc_hd__inv_2 _0615_ (.A(net80),
    .Y(\mux_top_track_8.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0616_ (.A(net75),
    .Y(\mux_top_track_8.INVTX1_0_.out ));
 sky130_fd_sc_hd__clkinv_2 _0617_ (.A(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out ),
    .Y(\mux_top_track_16.out ));
 sky130_fd_sc_hd__inv_2 _0618_ (.A(net81),
    .Y(\mux_top_track_16.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0619_ (.A(net76),
    .Y(\mux_top_track_16.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0620_ (.A(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out ),
    .Y(\mux_bottom_track_1.out ));
 sky130_fd_sc_hd__inv_2 _0621_ (.A(net9),
    .Y(\mux_bottom_track_1.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _0622_ (.A(net21),
    .Y(\mux_bottom_track_1.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _0623_ (.A(net16),
    .Y(\mux_bottom_track_1.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _0624_ (.A(net29),
    .Y(\mux_bottom_track_1.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _0625_ (.A(net24),
    .Y(\mux_bottom_track_1.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _0626_ (.A(net54),
    .Y(\mux_bottom_track_1.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0627_ (.A(net65),
    .Y(\mux_bottom_track_1.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0628_ (.A(net50),
    .Y(\mux_bottom_track_1.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0629_ (.A(net4),
    .Y(\mux_bottom_track_1.INVTX1_8_.out ));
 sky130_fd_sc_hd__clkinv_2 _0630_ (.A(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out ),
    .Y(\mux_bottom_track_9.out ));
 sky130_fd_sc_hd__inv_2 _0631_ (.A(net10),
    .Y(\mux_bottom_track_9.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _0632_ (.A(net20),
    .Y(\mux_bottom_track_9.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _0633_ (.A(net15),
    .Y(\mux_bottom_track_9.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _0634_ (.A(net28),
    .Y(\mux_bottom_track_9.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _0635_ (.A(net23),
    .Y(\mux_bottom_track_9.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _0636_ (.A(net55),
    .Y(\mux_bottom_track_9.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0637_ (.A(net67),
    .Y(\mux_bottom_track_9.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0638_ (.A(net60),
    .Y(\mux_bottom_track_9.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0639_ (.A(net5),
    .Y(\mux_bottom_track_9.INVTX1_8_.out ));
 sky130_fd_sc_hd__inv_2 _0640_ (.A(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out ),
    .Y(\mux_bottom_track_17.out ));
 sky130_fd_sc_hd__inv_2 _0641_ (.A(net1),
    .Y(\mux_bottom_track_17.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _0642_ (.A(net19),
    .Y(\mux_bottom_track_17.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _0643_ (.A(net14),
    .Y(\mux_bottom_track_17.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _0644_ (.A(net27),
    .Y(\mux_bottom_track_17.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _0645_ (.A(net22),
    .Y(\mux_bottom_track_17.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _0646_ (.A(net57),
    .Y(\mux_bottom_track_17.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0647_ (.A(net68),
    .Y(\mux_bottom_track_17.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0648_ (.A(net61),
    .Y(\mux_bottom_track_17.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0649_ (.A(net6),
    .Y(\mux_bottom_track_17.INVTX1_8_.out ));
 sky130_fd_sc_hd__inv_2 _0650_ (.A(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out ),
    .Y(\mux_bottom_track_25.out ));
 sky130_fd_sc_hd__inv_2 _0651_ (.A(net2),
    .Y(\mux_bottom_track_25.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _0652_ (.A(net18),
    .Y(\mux_bottom_track_25.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _0653_ (.A(net13),
    .Y(\mux_bottom_track_25.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _0654_ (.A(net26),
    .Y(\mux_bottom_track_25.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _0655_ (.A(net12),
    .Y(\mux_bottom_track_25.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _0656_ (.A(net58),
    .Y(\mux_bottom_track_25.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0657_ (.A(net51),
    .Y(\mux_bottom_track_25.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0658_ (.A(net63),
    .Y(\mux_bottom_track_25.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0659_ (.A(net7),
    .Y(\mux_bottom_track_25.INVTX1_8_.out ));
 sky130_fd_sc_hd__inv_2 _0660_ (.A(\mux_top_track_24.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(\mux_top_track_24.out ));
 sky130_fd_sc_hd__clkinv_2 _0661_ (.A(net82),
    .Y(\mux_top_track_24.INVTX1_1_.out ));
 sky130_fd_sc_hd__clkinv_2 _0662_ (.A(net77),
    .Y(\mux_top_track_24.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0663_ (.A(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(\mux_top_track_32.out ));
 sky130_fd_sc_hd__inv_2 _0664_ (.A(net83),
    .Y(\mux_top_track_32.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0665_ (.A(net78),
    .Y(\mux_top_track_32.INVTX1_0_.out ));
 sky130_fd_sc_hd__clkinv_2 _0666_ (.A(\mux_right_track_0.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .Y(\mux_right_track_0.out ));
 sky130_fd_sc_hd__inv_2 _0667_ (.A(net73),
    .Y(\mux_right_track_0.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0668_ (.A(net72),
    .Y(\mux_right_track_0.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0669_ (.A(net31),
    .Y(\mux_right_track_0.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _0670_ (.A(\mux_right_track_6.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .Y(\mux_right_track_6.out ));
 sky130_fd_sc_hd__inv_2 _0671_ (.A(net52),
    .Y(\mux_right_track_6.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0672_ (.A(net44),
    .Y(\mux_right_track_6.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _0673_ (.A(\mux_right_track_2.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .Y(\mux_right_track_2.out ));
 sky130_fd_sc_hd__inv_2 _0674_ (.A(net70),
    .Y(\mux_right_track_2.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _0675_ (.A(net62),
    .Y(\mux_right_track_2.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0676_ (.A(net41),
    .Y(\mux_right_track_2.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _0677_ (.A(\mux_right_track_4.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .Y(\mux_right_track_4.out ));
 sky130_fd_sc_hd__clkinv_2 _0678_ (.A(net66),
    .Y(\mux_right_track_4.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0679_ (.A(net42),
    .Y(\mux_right_track_4.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _0680_ (.A(\mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_right_track_8.out ));
 sky130_fd_sc_hd__inv_2 _0681_ (.A(net56),
    .Y(\mux_right_track_8.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0682_ (.A(net45),
    .Y(\mux_right_track_8.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0683_ (.A(\mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_right_track_10.out ));
 sky130_fd_sc_hd__inv_2 _0684_ (.A(net59),
    .Y(\mux_right_track_10.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0685_ (.A(net46),
    .Y(\mux_right_track_10.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0686_ (.A(\mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_right_track_18.out ));
 sky130_fd_sc_hd__inv_2 _0687_ (.A(net34),
    .Y(\mux_right_track_18.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0688_ (.A(\mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_right_track_20.out ));
 sky130_fd_sc_hd__inv_2 _0689_ (.A(net35),
    .Y(\mux_right_track_20.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0690_ (.A(\mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_right_track_22.out ));
 sky130_fd_sc_hd__inv_2 _0691_ (.A(net36),
    .Y(\mux_right_track_22.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0692_ (.A(\mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_right_track_24.out ));
 sky130_fd_sc_hd__inv_2 _0693_ (.A(net71),
    .Y(\mux_right_track_24.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0694_ (.A(net38),
    .Y(\mux_right_track_24.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0695_ (.A(\mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_right_track_26.out ));
 sky130_fd_sc_hd__inv_2 _0696_ (.A(net39),
    .Y(\mux_right_track_26.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0697_ (.A(net40),
    .Y(\mux_right_track_26.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0698_ (.A(\mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_right_track_12.out ));
 sky130_fd_sc_hd__inv_2 _0699_ (.A(net48),
    .Y(\mux_right_track_12.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0700_ (.A(\mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_right_track_14.out ));
 sky130_fd_sc_hd__inv_2 _0701_ (.A(net49),
    .Y(\mux_right_track_14.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0702_ (.A(\mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_right_track_16.out ));
 sky130_fd_sc_hd__inv_2 _0703_ (.A(net32),
    .Y(\mux_right_track_16.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0704_ (.A(\mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .Y(\mux_bottom_track_33.out ));
 sky130_fd_sc_hd__inv_2 _0705_ (.A(net3),
    .Y(\mux_bottom_track_33.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _0706_ (.A(net17),
    .Y(\mux_bottom_track_33.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _0707_ (.A(net30),
    .Y(\mux_bottom_track_33.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _0708_ (.A(net25),
    .Y(\mux_bottom_track_33.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0709_ (.A(net53),
    .Y(\mux_bottom_track_33.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0710_ (.A(net64),
    .Y(\mux_bottom_track_33.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0711_ (.A(net8),
    .Y(\mux_bottom_track_33.INVTX1_6_.out ));
 sky130_fd_sc_hd__clkbuf_4 _0712_ (.A(net69),
    .X(_0153_));
 sky130_fd_sc_hd__buf_4 _0713_ (.A(_0153_),
    .X(_0154_));
 sky130_fd_sc_hd__buf_4 _0714_ (.A(_0154_),
    .X(_0155_));
 sky130_fd_sc_hd__inv_2 _0715_ (.A(_0155_),
    .Y(_0072_));
 sky130_fd_sc_hd__inv_2 _0716_ (.A(_0155_),
    .Y(_0073_));
 sky130_fd_sc_hd__inv_2 _0717_ (.A(_0155_),
    .Y(_0074_));
 sky130_fd_sc_hd__inv_2 _0718_ (.A(_0155_),
    .Y(_0075_));
 sky130_fd_sc_hd__inv_2 _0719_ (.A(_0155_),
    .Y(_0076_));
 sky130_fd_sc_hd__inv_2 _0720_ (.A(_0155_),
    .Y(_0077_));
 sky130_fd_sc_hd__inv_2 _0721_ (.A(_0155_),
    .Y(_0078_));
 sky130_fd_sc_hd__inv_2 _0722_ (.A(_0155_),
    .Y(_0079_));
 sky130_fd_sc_hd__inv_2 _0723_ (.A(_0155_),
    .Y(_0080_));
 sky130_fd_sc_hd__inv_2 _0724_ (.A(_0155_),
    .Y(_0081_));
 sky130_fd_sc_hd__buf_4 _0725_ (.A(_0154_),
    .X(_0156_));
 sky130_fd_sc_hd__inv_2 _0726_ (.A(_0156_),
    .Y(_0082_));
 sky130_fd_sc_hd__inv_2 _0727_ (.A(_0156_),
    .Y(_0083_));
 sky130_fd_sc_hd__inv_2 _0728_ (.A(_0156_),
    .Y(_0084_));
 sky130_fd_sc_hd__inv_2 _0729_ (.A(_0156_),
    .Y(_0085_));
 sky130_fd_sc_hd__inv_2 _0730_ (.A(_0156_),
    .Y(_0086_));
 sky130_fd_sc_hd__inv_2 _0731_ (.A(_0156_),
    .Y(_0087_));
 sky130_fd_sc_hd__inv_2 _0732_ (.A(_0156_),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_2 _0733_ (.A(_0156_),
    .Y(_0089_));
 sky130_fd_sc_hd__inv_2 _0734_ (.A(_0156_),
    .Y(_0090_));
 sky130_fd_sc_hd__inv_2 _0735_ (.A(_0156_),
    .Y(_0091_));
 sky130_fd_sc_hd__buf_4 _0736_ (.A(_0153_),
    .X(_0157_));
 sky130_fd_sc_hd__inv_2 _0737_ (.A(_0157_),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_2 _0738_ (.A(_0157_),
    .Y(_0093_));
 sky130_fd_sc_hd__inv_2 _0739_ (.A(_0157_),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_2 _0740_ (.A(_0157_),
    .Y(_0095_));
 sky130_fd_sc_hd__inv_2 _0741_ (.A(_0157_),
    .Y(_0096_));
 sky130_fd_sc_hd__inv_2 _0742_ (.A(_0157_),
    .Y(_0097_));
 sky130_fd_sc_hd__inv_2 _0743_ (.A(_0157_),
    .Y(_0098_));
 sky130_fd_sc_hd__inv_2 _0744_ (.A(_0157_),
    .Y(_0099_));
 sky130_fd_sc_hd__inv_2 _0745_ (.A(_0157_),
    .Y(_0100_));
 sky130_fd_sc_hd__inv_2 _0746_ (.A(_0157_),
    .Y(_0101_));
 sky130_fd_sc_hd__buf_4 _0747_ (.A(_0153_),
    .X(_0118_));
 sky130_fd_sc_hd__inv_2 _0748_ (.A(_0118_),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_2 _0749_ (.A(_0118_),
    .Y(_0103_));
 sky130_fd_sc_hd__inv_2 _0750_ (.A(_0118_),
    .Y(_0104_));
 sky130_fd_sc_hd__inv_2 _0751_ (.A(_0118_),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_2 _0752_ (.A(_0118_),
    .Y(_0106_));
 sky130_fd_sc_hd__inv_2 _0753_ (.A(_0118_),
    .Y(_0107_));
 sky130_fd_sc_hd__inv_2 _0754_ (.A(_0118_),
    .Y(_0108_));
 sky130_fd_sc_hd__inv_2 _0755_ (.A(_0118_),
    .Y(_0109_));
 sky130_fd_sc_hd__inv_2 _0756_ (.A(_0118_),
    .Y(_0110_));
 sky130_fd_sc_hd__inv_2 _0757_ (.A(_0118_),
    .Y(_0111_));
 sky130_fd_sc_hd__buf_4 _0758_ (.A(_0153_),
    .X(_0119_));
 sky130_fd_sc_hd__inv_2 _0759_ (.A(_0119_),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_2 _0760_ (.A(_0119_),
    .Y(_0113_));
 sky130_fd_sc_hd__inv_2 _0761_ (.A(_0119_),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_2 _0762_ (.A(_0119_),
    .Y(_0115_));
 sky130_fd_sc_hd__inv_2 _0763_ (.A(_0119_),
    .Y(_0116_));
 sky130_fd_sc_hd__inv_2 _0764_ (.A(_0119_),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_2 _0765_ (.A(_0119_),
    .Y(_0000_));
 sky130_fd_sc_hd__inv_2 _0766_ (.A(_0119_),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _0767_ (.A(_0119_),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _0768_ (.A(_0119_),
    .Y(_0003_));
 sky130_fd_sc_hd__buf_4 _0769_ (.A(_0153_),
    .X(_0120_));
 sky130_fd_sc_hd__inv_2 _0770_ (.A(_0120_),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _0771_ (.A(_0120_),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _0772_ (.A(_0120_),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _0773_ (.A(_0120_),
    .Y(_0007_));
 sky130_fd_sc_hd__inv_2 _0774_ (.A(_0120_),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _0775_ (.A(_0120_),
    .Y(_0009_));
 sky130_fd_sc_hd__inv_2 _0776_ (.A(_0120_),
    .Y(_0010_));
 sky130_fd_sc_hd__inv_2 _0777_ (.A(_0120_),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_2 _0778_ (.A(_0120_),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_2 _0779_ (.A(_0120_),
    .Y(_0013_));
 sky130_fd_sc_hd__clkbuf_8 _0780_ (.A(_0153_),
    .X(_0121_));
 sky130_fd_sc_hd__inv_2 _0781_ (.A(_0121_),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _0782_ (.A(_0121_),
    .Y(_0015_));
 sky130_fd_sc_hd__inv_2 _0783_ (.A(_0121_),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_2 _0784_ (.A(_0121_),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _0785_ (.A(_0121_),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_2 _0786_ (.A(_0121_),
    .Y(_0019_));
 sky130_fd_sc_hd__inv_2 _0787_ (.A(_0121_),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_2 _0788_ (.A(_0121_),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _0789_ (.A(_0121_),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _0790_ (.A(_0121_),
    .Y(_0023_));
 sky130_fd_sc_hd__clkbuf_8 _0791_ (.A(_0153_),
    .X(_0122_));
 sky130_fd_sc_hd__inv_2 _0792_ (.A(_0122_),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _0793_ (.A(_0122_),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _0794_ (.A(_0122_),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _0795_ (.A(_0122_),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _0796_ (.A(_0122_),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _0797_ (.A(_0122_),
    .Y(_0029_));
 sky130_fd_sc_hd__inv_2 _0798_ (.A(_0122_),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_2 _0799_ (.A(_0122_),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _0800_ (.A(_0122_),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _0801_ (.A(_0122_),
    .Y(_0033_));
 sky130_fd_sc_hd__buf_4 _0802_ (.A(_0153_),
    .X(_0123_));
 sky130_fd_sc_hd__inv_2 _0803_ (.A(_0123_),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _0804_ (.A(_0123_),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _0805_ (.A(_0123_),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _0806_ (.A(_0123_),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _0807_ (.A(_0123_),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _0808_ (.A(_0123_),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_2 _0809_ (.A(_0123_),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _0810_ (.A(_0123_),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_2 _0811_ (.A(_0123_),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _0812_ (.A(_0123_),
    .Y(_0043_));
 sky130_fd_sc_hd__buf_4 _0813_ (.A(_0153_),
    .X(_0124_));
 sky130_fd_sc_hd__inv_2 _0814_ (.A(_0124_),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _0815_ (.A(_0124_),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_2 _0816_ (.A(_0124_),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_2 _0817_ (.A(_0124_),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_2 _0818_ (.A(_0124_),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_2 _0819_ (.A(_0124_),
    .Y(_0049_));
 sky130_fd_sc_hd__inv_2 _0820_ (.A(_0124_),
    .Y(_0050_));
 sky130_fd_sc_hd__inv_2 _0821_ (.A(_0124_),
    .Y(_0051_));
 sky130_fd_sc_hd__inv_2 _0822_ (.A(_0124_),
    .Y(_0052_));
 sky130_fd_sc_hd__inv_2 _0823_ (.A(_0124_),
    .Y(_0053_));
 sky130_fd_sc_hd__buf_4 _0824_ (.A(_0153_),
    .X(_0125_));
 sky130_fd_sc_hd__inv_2 _0825_ (.A(_0125_),
    .Y(_0054_));
 sky130_fd_sc_hd__inv_2 _0826_ (.A(_0125_),
    .Y(_0055_));
 sky130_fd_sc_hd__inv_2 _0827_ (.A(_0125_),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_2 _0828_ (.A(_0125_),
    .Y(_0057_));
 sky130_fd_sc_hd__inv_2 _0829_ (.A(_0125_),
    .Y(_0058_));
 sky130_fd_sc_hd__inv_2 _0830_ (.A(_0125_),
    .Y(_0059_));
 sky130_fd_sc_hd__inv_2 _0831_ (.A(_0125_),
    .Y(_0060_));
 sky130_fd_sc_hd__inv_2 _0832_ (.A(_0125_),
    .Y(_0061_));
 sky130_fd_sc_hd__inv_2 _0833_ (.A(_0125_),
    .Y(_0062_));
 sky130_fd_sc_hd__inv_2 _0834_ (.A(_0125_),
    .Y(_0063_));
 sky130_fd_sc_hd__inv_2 _0835_ (.A(_0154_),
    .Y(_0064_));
 sky130_fd_sc_hd__inv_2 _0836_ (.A(_0154_),
    .Y(_0065_));
 sky130_fd_sc_hd__inv_2 _0837_ (.A(_0154_),
    .Y(_0066_));
 sky130_fd_sc_hd__inv_2 _0838_ (.A(_0154_),
    .Y(_0067_));
 sky130_fd_sc_hd__inv_2 _0839_ (.A(_0154_),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_2 _0840_ (.A(_0154_),
    .Y(_0069_));
 sky130_fd_sc_hd__inv_2 _0841_ (.A(_0154_),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_2 _0842_ (.A(_0154_),
    .Y(_0071_));
 sky130_fd_sc_hd__dfrtp_1 _0843_ (.CLK(clknet_4_14_0_prog_clk),
    .D(\mem_top_track_0.DFFR_6_.Q ),
    .RESET_B(_0072_),
    .Q(\mem_top_track_0.DFFR_7_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0844_ (.CLK(clknet_4_14_0_prog_clk),
    .D(\mem_top_track_0.DFFR_5_.Q ),
    .RESET_B(_0073_),
    .Q(\mem_top_track_0.DFFR_6_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0845_ (.CLK(clknet_4_14_0_prog_clk),
    .D(\mem_top_track_0.DFFR_4_.Q ),
    .RESET_B(_0074_),
    .Q(\mem_top_track_0.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0846_ (.CLK(clknet_4_14_0_prog_clk),
    .D(\mem_top_track_0.DFFR_3_.Q ),
    .RESET_B(_0075_),
    .Q(\mem_top_track_0.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0847_ (.CLK(clknet_4_15_0_prog_clk),
    .D(\mem_top_track_0.DFFR_2_.Q ),
    .RESET_B(_0076_),
    .Q(\mem_top_track_0.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0848_ (.CLK(clknet_4_13_0_prog_clk),
    .D(\mem_top_track_0.DFFR_1_.Q ),
    .RESET_B(_0077_),
    .Q(\mem_top_track_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0849_ (.CLK(clknet_4_13_0_prog_clk),
    .D(\mem_top_track_0.DFFR_0_.Q ),
    .RESET_B(_0078_),
    .Q(\mem_top_track_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0850_ (.CLK(clknet_4_3_0_prog_clk),
    .D(net11),
    .RESET_B(_0079_),
    .Q(\mem_top_track_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0851_ (.CLK(clknet_4_7_0_prog_clk),
    .D(\mem_top_track_8.DFFR_6_.Q ),
    .RESET_B(_0080_),
    .Q(\mem_top_track_16.DFFR_0_.D ));
 sky130_fd_sc_hd__dfrtp_1 _0852_ (.CLK(clknet_4_7_0_prog_clk),
    .D(\mem_top_track_8.DFFR_5_.Q ),
    .RESET_B(_0081_),
    .Q(\mem_top_track_8.DFFR_6_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0853_ (.CLK(clknet_4_7_0_prog_clk),
    .D(\mem_top_track_8.DFFR_4_.Q ),
    .RESET_B(_0082_),
    .Q(\mem_top_track_8.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0854_ (.CLK(clknet_4_6_0_prog_clk),
    .D(\mem_top_track_8.DFFR_3_.Q ),
    .RESET_B(_0083_),
    .Q(\mem_top_track_8.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0855_ (.CLK(clknet_4_0_0_prog_clk),
    .D(\mem_top_track_8.DFFR_2_.Q ),
    .RESET_B(_0084_),
    .Q(\mem_top_track_8.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0856_ (.CLK(clknet_4_1_0_prog_clk),
    .D(\mem_top_track_8.DFFR_1_.Q ),
    .RESET_B(_0085_),
    .Q(\mem_top_track_8.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0857_ (.CLK(clknet_4_1_0_prog_clk),
    .D(\mem_top_track_8.DFFR_0_.Q ),
    .RESET_B(_0086_),
    .Q(\mem_top_track_8.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0858_ (.CLK(clknet_4_14_0_prog_clk),
    .D(\mem_top_track_0.DFFR_7_.Q ),
    .RESET_B(_0087_),
    .Q(\mem_top_track_8.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0859_ (.CLK(clknet_4_1_0_prog_clk),
    .D(\mem_top_track_16.DFFR_6_.Q ),
    .RESET_B(_0088_),
    .Q(\mem_top_track_16.DFFR_7_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0860_ (.CLK(clknet_4_1_0_prog_clk),
    .D(\mem_top_track_16.DFFR_5_.Q ),
    .RESET_B(_0089_),
    .Q(\mem_top_track_16.DFFR_6_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0861_ (.CLK(clknet_4_4_0_prog_clk),
    .D(\mem_top_track_16.DFFR_4_.Q ),
    .RESET_B(_0090_),
    .Q(\mem_top_track_16.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0862_ (.CLK(clknet_4_5_0_prog_clk),
    .D(\mem_top_track_16.DFFR_3_.Q ),
    .RESET_B(_0091_),
    .Q(\mem_top_track_16.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0863_ (.CLK(clknet_4_5_0_prog_clk),
    .D(\mem_top_track_16.DFFR_2_.Q ),
    .RESET_B(_0092_),
    .Q(\mem_top_track_16.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0864_ (.CLK(clknet_4_5_0_prog_clk),
    .D(\mem_top_track_16.DFFR_1_.Q ),
    .RESET_B(_0093_),
    .Q(\mem_top_track_16.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0865_ (.CLK(clknet_4_13_0_prog_clk),
    .D(\mem_top_track_16.DFFR_0_.Q ),
    .RESET_B(_0094_),
    .Q(\mem_top_track_16.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0866_ (.CLK(clknet_4_7_0_prog_clk),
    .D(\mem_top_track_16.DFFR_0_.D ),
    .RESET_B(_0095_),
    .Q(\mem_top_track_16.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0867_ (.CLK(clknet_4_3_0_prog_clk),
    .D(\mem_bottom_track_1.DFFR_6_.Q ),
    .RESET_B(_0096_),
    .Q(\mem_bottom_track_1.DFFR_7_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0868_ (.CLK(clknet_4_3_0_prog_clk),
    .D(\mem_bottom_track_1.DFFR_5_.Q ),
    .RESET_B(_0097_),
    .Q(\mem_bottom_track_1.DFFR_6_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0869_ (.CLK(clknet_4_4_0_prog_clk),
    .D(\mem_bottom_track_1.DFFR_4_.Q ),
    .RESET_B(_0098_),
    .Q(\mem_bottom_track_1.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0870_ (.CLK(clknet_4_6_0_prog_clk),
    .D(\mem_bottom_track_1.DFFR_3_.Q ),
    .RESET_B(_0099_),
    .Q(\mem_bottom_track_1.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0871_ (.CLK(clknet_4_5_0_prog_clk),
    .D(\mem_bottom_track_1.DFFR_2_.Q ),
    .RESET_B(_0100_),
    .Q(\mem_bottom_track_1.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0872_ (.CLK(clknet_4_6_0_prog_clk),
    .D(\mem_bottom_track_1.DFFR_1_.Q ),
    .RESET_B(_0101_),
    .Q(\mem_bottom_track_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0873_ (.CLK(clknet_4_6_0_prog_clk),
    .D(\mem_bottom_track_1.DFFR_0_.Q ),
    .RESET_B(_0102_),
    .Q(\mem_bottom_track_1.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0874_ (.CLK(clknet_4_6_0_prog_clk),
    .D(\mem_bottom_track_1.DFFR_0_.D ),
    .RESET_B(_0103_),
    .Q(\mem_bottom_track_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0875_ (.CLK(clknet_4_10_0_prog_clk),
    .D(\mem_bottom_track_9.DFFR_6_.Q ),
    .RESET_B(_0104_),
    .Q(\mem_bottom_track_17.DFFR_0_.D ));
 sky130_fd_sc_hd__dfrtp_1 _0876_ (.CLK(clknet_4_10_0_prog_clk),
    .D(\mem_bottom_track_9.DFFR_5_.Q ),
    .RESET_B(_0105_),
    .Q(\mem_bottom_track_9.DFFR_6_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0877_ (.CLK(clknet_4_10_0_prog_clk),
    .D(\mem_bottom_track_9.DFFR_4_.Q ),
    .RESET_B(_0106_),
    .Q(\mem_bottom_track_9.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0878_ (.CLK(clknet_4_9_0_prog_clk),
    .D(\mem_bottom_track_9.DFFR_3_.Q ),
    .RESET_B(_0107_),
    .Q(\mem_bottom_track_9.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0879_ (.CLK(clknet_4_3_0_prog_clk),
    .D(\mem_bottom_track_9.DFFR_2_.Q ),
    .RESET_B(_0108_),
    .Q(\mem_bottom_track_9.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0880_ (.CLK(clknet_4_12_0_prog_clk),
    .D(\mem_bottom_track_9.DFFR_1_.Q ),
    .RESET_B(_0109_),
    .Q(\mem_bottom_track_9.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0881_ (.CLK(clknet_4_9_0_prog_clk),
    .D(\mem_bottom_track_9.DFFR_0_.Q ),
    .RESET_B(_0110_),
    .Q(\mem_bottom_track_9.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0882_ (.CLK(clknet_4_4_0_prog_clk),
    .D(\mem_bottom_track_1.DFFR_7_.Q ),
    .RESET_B(_0111_),
    .Q(\mem_bottom_track_9.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0883_ (.CLK(clknet_4_10_0_prog_clk),
    .D(\mem_bottom_track_17.DFFR_6_.Q ),
    .RESET_B(_0112_),
    .Q(\mem_bottom_track_17.DFFR_7_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0884_ (.CLK(clknet_4_10_0_prog_clk),
    .D(\mem_bottom_track_17.DFFR_5_.Q ),
    .RESET_B(_0113_),
    .Q(\mem_bottom_track_17.DFFR_6_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0885_ (.CLK(clknet_4_10_0_prog_clk),
    .D(\mem_bottom_track_17.DFFR_4_.Q ),
    .RESET_B(_0114_),
    .Q(\mem_bottom_track_17.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0886_ (.CLK(clknet_4_14_0_prog_clk),
    .D(\mem_bottom_track_17.DFFR_3_.Q ),
    .RESET_B(_0115_),
    .Q(\mem_bottom_track_17.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0887_ (.CLK(clknet_4_6_0_prog_clk),
    .D(\mem_bottom_track_17.DFFR_2_.Q ),
    .RESET_B(_0116_),
    .Q(\mem_bottom_track_17.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0888_ (.CLK(clknet_4_12_0_prog_clk),
    .D(\mem_bottom_track_17.DFFR_1_.Q ),
    .RESET_B(_0117_),
    .Q(\mem_bottom_track_17.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0889_ (.CLK(clknet_4_10_0_prog_clk),
    .D(\mem_bottom_track_17.DFFR_0_.Q ),
    .RESET_B(_0000_),
    .Q(\mem_bottom_track_17.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0890_ (.CLK(clknet_4_10_0_prog_clk),
    .D(\mem_bottom_track_17.DFFR_0_.D ),
    .RESET_B(_0001_),
    .Q(\mem_bottom_track_17.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0891_ (.CLK(clknet_4_0_0_prog_clk),
    .D(\mem_bottom_track_25.DFFR_6_.Q ),
    .RESET_B(_0002_),
    .Q(\mem_bottom_track_25.DFFR_7_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0892_ (.CLK(clknet_4_2_0_prog_clk),
    .D(\mem_bottom_track_25.DFFR_5_.Q ),
    .RESET_B(_0003_),
    .Q(\mem_bottom_track_25.DFFR_6_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0893_ (.CLK(clknet_4_0_0_prog_clk),
    .D(\mem_bottom_track_25.DFFR_4_.Q ),
    .RESET_B(_0004_),
    .Q(\mem_bottom_track_25.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0894_ (.CLK(clknet_4_0_0_prog_clk),
    .D(\mem_bottom_track_25.DFFR_3_.Q ),
    .RESET_B(_0005_),
    .Q(\mem_bottom_track_25.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0895_ (.CLK(clknet_4_0_0_prog_clk),
    .D(\mem_bottom_track_25.DFFR_2_.Q ),
    .RESET_B(_0006_),
    .Q(\mem_bottom_track_25.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0896_ (.CLK(clknet_4_2_0_prog_clk),
    .D(\mem_bottom_track_25.DFFR_1_.Q ),
    .RESET_B(_0007_),
    .Q(\mem_bottom_track_25.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0897_ (.CLK(clknet_4_1_0_prog_clk),
    .D(\mem_bottom_track_25.DFFR_0_.Q ),
    .RESET_B(_0008_),
    .Q(\mem_bottom_track_25.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0898_ (.CLK(clknet_4_9_0_prog_clk),
    .D(\mem_bottom_track_17.DFFR_7_.Q ),
    .RESET_B(_0009_),
    .Q(\mem_bottom_track_25.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0899_ (.CLK(clknet_4_12_0_prog_clk),
    .D(\mem_top_track_24.DFFR_4_.Q ),
    .RESET_B(_0010_),
    .Q(\mem_top_track_24.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0900_ (.CLK(clknet_4_10_0_prog_clk),
    .D(\mem_top_track_24.DFFR_3_.Q ),
    .RESET_B(_0011_),
    .Q(\mem_top_track_24.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0901_ (.CLK(clknet_4_8_0_prog_clk),
    .D(\mem_top_track_24.DFFR_2_.Q ),
    .RESET_B(_0012_),
    .Q(\mem_top_track_24.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0902_ (.CLK(clknet_4_2_0_prog_clk),
    .D(\mem_top_track_24.DFFR_1_.Q ),
    .RESET_B(_0013_),
    .Q(\mem_top_track_24.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0903_ (.CLK(clknet_4_2_0_prog_clk),
    .D(\mem_top_track_24.DFFR_0_.Q ),
    .RESET_B(_0014_),
    .Q(\mem_top_track_24.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0904_ (.CLK(clknet_4_3_0_prog_clk),
    .D(\mem_top_track_16.DFFR_7_.Q ),
    .RESET_B(_0015_),
    .Q(\mem_top_track_24.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0905_ (.CLK(clknet_4_5_0_prog_clk),
    .D(\mem_top_track_32.DFFR_4_.Q ),
    .RESET_B(_0016_),
    .Q(\mem_right_track_0.DFFR_0_.D ));
 sky130_fd_sc_hd__dfrtp_1 _0906_ (.CLK(clknet_4_7_0_prog_clk),
    .D(\mem_top_track_32.DFFR_3_.Q ),
    .RESET_B(_0017_),
    .Q(\mem_top_track_32.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0907_ (.CLK(clknet_4_6_0_prog_clk),
    .D(\mem_top_track_32.DFFR_2_.Q ),
    .RESET_B(_0018_),
    .Q(\mem_top_track_32.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0908_ (.CLK(clknet_4_4_0_prog_clk),
    .D(\mem_top_track_32.DFFR_1_.Q ),
    .RESET_B(_0019_),
    .Q(\mem_top_track_32.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0909_ (.CLK(clknet_4_1_0_prog_clk),
    .D(\mem_top_track_32.DFFR_0_.Q ),
    .RESET_B(_0020_),
    .Q(\mem_top_track_32.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0910_ (.CLK(clknet_4_13_0_prog_clk),
    .D(\mem_top_track_24.DFFR_5_.Q ),
    .RESET_B(_0021_),
    .Q(\mem_top_track_32.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0911_ (.CLK(clknet_4_15_0_prog_clk),
    .D(\mem_right_track_0.DFFR_4_.Q ),
    .RESET_B(_0022_),
    .Q(\mem_right_track_0.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0912_ (.CLK(clknet_4_13_0_prog_clk),
    .D(\mem_right_track_0.DFFR_3_.Q ),
    .RESET_B(_0023_),
    .Q(\mem_right_track_0.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0913_ (.CLK(clknet_4_7_0_prog_clk),
    .D(\mem_right_track_0.DFFR_2_.Q ),
    .RESET_B(_0024_),
    .Q(\mem_right_track_0.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0914_ (.CLK(clknet_4_6_0_prog_clk),
    .D(\mem_right_track_0.DFFR_1_.Q ),
    .RESET_B(_0025_),
    .Q(\mem_right_track_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0915_ (.CLK(clknet_4_4_0_prog_clk),
    .D(\mem_right_track_0.DFFR_0_.Q ),
    .RESET_B(_0026_),
    .Q(\mem_right_track_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0916_ (.CLK(clknet_4_4_0_prog_clk),
    .D(\mem_right_track_0.DFFR_0_.D ),
    .RESET_B(_0027_),
    .Q(\mem_right_track_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0917_ (.CLK(clknet_4_4_0_prog_clk),
    .D(\mem_right_track_6.DFFR_4_.Q ),
    .RESET_B(_0028_),
    .Q(\mem_right_track_6.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0918_ (.CLK(clknet_4_5_0_prog_clk),
    .D(\mem_right_track_6.DFFR_3_.Q ),
    .RESET_B(_0029_),
    .Q(\mem_right_track_6.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0919_ (.CLK(clknet_4_7_0_prog_clk),
    .D(\mem_right_track_6.DFFR_2_.Q ),
    .RESET_B(_0030_),
    .Q(\mem_right_track_6.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0920_ (.CLK(clknet_4_7_0_prog_clk),
    .D(\mem_right_track_6.DFFR_1_.Q ),
    .RESET_B(_0031_),
    .Q(\mem_right_track_6.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0921_ (.CLK(clknet_4_7_0_prog_clk),
    .D(\mem_right_track_6.DFFR_0_.Q ),
    .RESET_B(_0032_),
    .Q(\mem_right_track_6.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0922_ (.CLK(clknet_4_7_0_prog_clk),
    .D(\mem_right_track_4.DFFR_5_.Q ),
    .RESET_B(_0033_),
    .Q(\mem_right_track_6.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0923_ (.CLK(clknet_4_11_0_prog_clk),
    .D(\mem_right_track_2.DFFR_4_.Q ),
    .RESET_B(_0034_),
    .Q(\mem_right_track_2.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0924_ (.CLK(clknet_4_11_0_prog_clk),
    .D(\mem_right_track_2.DFFR_3_.Q ),
    .RESET_B(_0035_),
    .Q(\mem_right_track_2.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0925_ (.CLK(clknet_4_8_0_prog_clk),
    .D(\mem_right_track_2.DFFR_2_.Q ),
    .RESET_B(_0036_),
    .Q(\mem_right_track_2.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0926_ (.CLK(clknet_4_2_0_prog_clk),
    .D(\mem_right_track_2.DFFR_1_.Q ),
    .RESET_B(_0037_),
    .Q(\mem_right_track_2.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0927_ (.CLK(clknet_4_9_0_prog_clk),
    .D(\mem_right_track_2.DFFR_0_.Q ),
    .RESET_B(_0038_),
    .Q(\mem_right_track_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0928_ (.CLK(clknet_4_15_0_prog_clk),
    .D(\mem_right_track_0.DFFR_5_.Q ),
    .RESET_B(_0039_),
    .Q(\mem_right_track_2.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0929_ (.CLK(clknet_4_15_0_prog_clk),
    .D(\mem_right_track_4.DFFR_4_.Q ),
    .RESET_B(_0040_),
    .Q(\mem_right_track_4.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0930_ (.CLK(clknet_4_15_0_prog_clk),
    .D(\mem_right_track_4.DFFR_3_.Q ),
    .RESET_B(_0041_),
    .Q(\mem_right_track_4.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0931_ (.CLK(clknet_4_15_0_prog_clk),
    .D(\mem_right_track_4.DFFR_2_.Q ),
    .RESET_B(_0042_),
    .Q(\mem_right_track_4.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0932_ (.CLK(clknet_4_15_0_prog_clk),
    .D(\mem_right_track_4.DFFR_1_.Q ),
    .RESET_B(_0043_),
    .Q(\mem_right_track_4.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0933_ (.CLK(clknet_4_12_0_prog_clk),
    .D(\mem_right_track_4.DFFR_0_.Q ),
    .RESET_B(_0044_),
    .Q(\mem_right_track_4.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0934_ (.CLK(clknet_4_11_0_prog_clk),
    .D(\mem_right_track_2.DFFR_5_.Q ),
    .RESET_B(_0045_),
    .Q(\mem_right_track_4.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0935_ (.CLK(clknet_4_8_0_prog_clk),
    .D(\mem_right_track_8.DFFR_0_.Q ),
    .RESET_B(_0046_),
    .Q(\mem_right_track_10.DFFR_0_.D ));
 sky130_fd_sc_hd__dfrtp_4 _0936_ (.CLK(clknet_4_13_0_prog_clk),
    .D(\mem_right_track_6.DFFR_5_.Q ),
    .RESET_B(_0047_),
    .Q(\mem_right_track_8.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0937_ (.CLK(clknet_4_1_0_prog_clk),
    .D(\mem_right_track_10.DFFR_0_.Q ),
    .RESET_B(_0048_),
    .Q(\mem_right_track_10.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0938_ (.CLK(clknet_4_11_0_prog_clk),
    .D(\mem_right_track_10.DFFR_0_.D ),
    .RESET_B(_0049_),
    .Q(\mem_right_track_10.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0939_ (.CLK(clknet_4_2_0_prog_clk),
    .D(\mem_right_track_18.DFFR_0_.Q ),
    .RESET_B(_0050_),
    .Q(\mem_right_track_18.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0940_ (.CLK(clknet_4_10_0_prog_clk),
    .D(\mem_right_track_16.DFFR_1_.Q ),
    .RESET_B(_0051_),
    .Q(\mem_right_track_18.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0941_ (.CLK(clknet_4_11_0_prog_clk),
    .D(\mem_right_track_20.DFFR_0_.Q ),
    .RESET_B(_0052_),
    .Q(\mem_right_track_20.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0942_ (.CLK(clknet_4_8_0_prog_clk),
    .D(\mem_right_track_18.DFFR_1_.Q ),
    .RESET_B(_0053_),
    .Q(\mem_right_track_20.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0943_ (.CLK(clknet_4_8_0_prog_clk),
    .D(\mem_right_track_22.DFFR_0_.Q ),
    .RESET_B(_0054_),
    .Q(\mem_right_track_22.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0944_ (.CLK(clknet_4_11_0_prog_clk),
    .D(\mem_right_track_20.DFFR_1_.Q ),
    .RESET_B(_0055_),
    .Q(\mem_right_track_22.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0945_ (.CLK(clknet_4_1_0_prog_clk),
    .D(\mem_right_track_24.DFFR_0_.Q ),
    .RESET_B(_0056_),
    .Q(\mem_right_track_24.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0946_ (.CLK(clknet_4_2_0_prog_clk),
    .D(\mem_right_track_22.DFFR_1_.Q ),
    .RESET_B(_0057_),
    .Q(\mem_right_track_24.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0947_ (.CLK(clknet_4_3_0_prog_clk),
    .D(\mem_right_track_26.DFFR_0_.Q ),
    .RESET_B(_0058_),
    .Q(\mem_bottom_track_1.DFFR_0_.D ));
 sky130_fd_sc_hd__dfrtp_4 _0948_ (.CLK(clknet_4_1_0_prog_clk),
    .D(\mem_right_track_24.DFFR_1_.Q ),
    .RESET_B(_0059_),
    .Q(\mem_right_track_26.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0949_ (.CLK(clknet_4_9_0_prog_clk),
    .D(\mem_right_track_12.DFFR_0_.Q ),
    .RESET_B(_0060_),
    .Q(\mem_right_track_12.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0950_ (.CLK(clknet_4_2_0_prog_clk),
    .D(\mem_right_track_10.DFFR_1_.Q ),
    .RESET_B(_0061_),
    .Q(\mem_right_track_12.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0951_ (.CLK(clknet_4_9_0_prog_clk),
    .D(\mem_right_track_14.DFFR_0_.Q ),
    .RESET_B(_0062_),
    .Q(\mem_right_track_14.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0952_ (.CLK(clknet_4_11_0_prog_clk),
    .D(\mem_right_track_12.DFFR_1_.Q ),
    .RESET_B(_0063_),
    .Q(\mem_right_track_14.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0953_ (.CLK(clknet_4_11_0_prog_clk),
    .D(\mem_right_track_16.DFFR_0_.Q ),
    .RESET_B(_0064_),
    .Q(\mem_right_track_16.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0954_ (.CLK(clknet_4_14_0_prog_clk),
    .D(\mem_right_track_14.DFFR_1_.Q ),
    .RESET_B(_0065_),
    .Q(\mem_right_track_16.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0955_ (.CLK(clknet_4_8_0_prog_clk),
    .D(\mem_bottom_track_33.DFFR_4_.Q ),
    .RESET_B(_0066_),
    .Q(net84));
 sky130_fd_sc_hd__dfrtp_1 _0956_ (.CLK(clknet_4_8_0_prog_clk),
    .D(\mem_bottom_track_33.DFFR_3_.Q ),
    .RESET_B(_0067_),
    .Q(\mem_bottom_track_33.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0957_ (.CLK(clknet_4_9_0_prog_clk),
    .D(\mem_bottom_track_33.DFFR_2_.Q ),
    .RESET_B(_0068_),
    .Q(\mem_bottom_track_33.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0958_ (.CLK(clknet_4_0_0_prog_clk),
    .D(\mem_bottom_track_33.DFFR_1_.Q ),
    .RESET_B(_0069_),
    .Q(\mem_bottom_track_33.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0959_ (.CLK(clknet_4_0_0_prog_clk),
    .D(\mem_bottom_track_33.DFFR_0_.Q ),
    .RESET_B(_0070_),
    .Q(\mem_bottom_track_33.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0960_ (.CLK(clknet_4_0_0_prog_clk),
    .D(\mem_bottom_track_25.DFFR_7_.Q ),
    .RESET_B(_0071_),
    .Q(\mem_bottom_track_33.DFFR_0_.Q ));
 sky130_fd_sc_hd__conb_1 _1056__143 (.HI(net143));
 sky130_fd_sc_hd__conb_1 _1068__144 (.HI(net144));
 sky130_fd_sc_hd__conb_1 _1080__145 (.HI(net145));
 sky130_fd_sc_hd__conb_1 _1092__146 (.HI(net146));
 sky130_fd_sc_hd__conb_1 _1104__147 (.HI(net147));
 sky130_fd_sc_hd__conb_1 _1116__148 (.HI(net148));
 sky130_fd_sc_hd__conb_1 _1129__149 (.HI(net149));
 sky130_fd_sc_hd__conb_1 _1141__150 (.HI(net150));
 sky130_fd_sc_hd__conb_1 _1151__151 (.HI(net151));
 sky130_fd_sc_hd__conb_1 _1157__152 (.HI(net152));
 sky130_fd_sc_hd__conb_1 _1164__153 (.HI(net153));
 sky130_fd_sc_hd__conb_1 _1172__154 (.HI(net154));
 sky130_fd_sc_hd__conb_1 _1179__155 (.HI(net155));
 sky130_fd_sc_hd__conb_1 _1185__156 (.HI(net156));
 sky130_fd_sc_hd__conb_1 _1191__157 (.HI(net157));
 sky130_fd_sc_hd__conb_1 _1197__158 (.HI(net158));
 sky130_fd_sc_hd__conb_1 _1203__159 (.HI(net159));
 sky130_fd_sc_hd__conb_1 _1209__160 (.HI(net160));
 sky130_fd_sc_hd__conb_1 _1215__161 (.HI(net161));
 sky130_fd_sc_hd__conb_1 _1220__162 (.HI(net162));
 sky130_fd_sc_hd__conb_1 _1224__163 (.HI(net163));
 sky130_fd_sc_hd__conb_1 _1228__164 (.HI(net164));
 sky130_fd_sc_hd__conb_1 _1232__165 (.HI(net165));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_prog_clk (.A(prog_clk),
    .X(clknet_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_1 _0985_ (.A(net72),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 _0986_ (.A(net43),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 _0987_ (.A(net47),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 _0988_ (.A(net33),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 _0989_ (.A(net37),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 _0990_ (.A(\mux_right_track_26.out ),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 _0991_ (.A(\mux_right_track_24.out ),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 _0992_ (.A(\mux_right_track_22.out ),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 _0993_ (.A(\mux_right_track_20.out ),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 _0994_ (.A(\mux_right_track_18.out ),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 _0995_ (.A(\mux_right_track_16.out ),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 _0996_ (.A(\mux_right_track_14.out ),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 _0997_ (.A(\mux_right_track_12.out ),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 _0998_ (.A(\mux_right_track_10.out ),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 _0999_ (.A(\mux_right_track_8.out ),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 _1000_ (.A(\mux_right_track_6.out ),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 _1001_ (.A(\mux_right_track_4.out ),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 _1002_ (.A(\mux_right_track_2.out ),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 _1003_ (.A(\mux_right_track_0.out ),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 _1004_ (.A(net58),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_2 _1005_ (.A(net57),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_1 _1006_ (.A(\mux_bottom_track_33.out ),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_1 _1007_ (.A(net55),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_2 _1008_ (.A(net54),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 _1009_ (.A(net53),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_1 _1010_ (.A(\mux_bottom_track_25.out ),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 _1011_ (.A(net51),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_2 _1012_ (.A(net68),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 _1013_ (.A(net67),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 _1014_ (.A(\mux_bottom_track_17.out ),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_2 _1015_ (.A(net65),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 _1016_ (.A(net64),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_2 _1017_ (.A(net63),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_1 _1018_ (.A(\mux_bottom_track_9.out ),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_2 _1019_ (.A(net61),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_2 _1020_ (.A(net60),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_1 _1021_ (.A(net50),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_1 _1022_ (.A(\mux_bottom_track_1.out ),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 _1023_ (.A(net39),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 _1024_ (.A(net38),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 _1025_ (.A(\mux_top_track_32.out ),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_1 _1026_ (.A(net36),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 _1027_ (.A(net35),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 _1028_ (.A(net34),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_1 _1029_ (.A(\mux_top_track_24.out ),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 _1030_ (.A(net32),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_2 _1031_ (.A(net49),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 _1032_ (.A(net48),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 _1033_ (.A(\mux_top_track_16.out ),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 _1034_ (.A(net46),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_1 _1035_ (.A(net45),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_1 _1036_ (.A(net44),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_1 _1037_ (.A(\mux_top_track_8.out ),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_1 _1038_ (.A(net42),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_2 _1039_ (.A(net41),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_2 _1040_ (.A(net31),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 _1041_ (.A(\mux_top_track_0.out ),
    .X(net123));
 sky130_fd_sc_hd__ebufn_2 _1042_ (.A(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out ),
    .TE_B(_0158_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1043_ (.A(\mux_right_track_20.INVTX1_2_.out ),
    .TE_B(_0159_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1044_ (.A(net142),
    .TE_B(_0160_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_8 _1045_ (.A(\mux_bottom_track_17.INVTX1_6_.out ),
    .TE_B(_0161_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_8 _1046_ (.A(\mux_right_track_0.INVTX1_3_.out ),
    .TE_B(_0162_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_8 _1047_ (.A(\mux_right_track_10.INVTX1_2_.out ),
    .TE_B(_0163_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1048_ (.A(\mux_top_track_0.INVTX1_1_.out ),
    .TE_B(_0164_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1049_ (.A(\mux_bottom_track_17.INVTX1_3_.out ),
    .TE_B(_0165_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1050_ (.A(\mux_bottom_track_17.INVTX1_4_.out ),
    .TE_B(_0166_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1051_ (.A(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out ),
    .TE_B(_0167_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_8 _1052_ (.A(\mux_bottom_track_17.INVTX1_5_.out ),
    .TE_B(_0168_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1053_ (.A(\mux_top_track_0.INVTX1_0_.out ),
    .TE_B(_0169_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1054_ (.A(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out ),
    .TE_B(_0170_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1055_ (.A(\mux_right_track_22.INVTX1_2_.out ),
    .TE_B(_0171_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1056_ (.A(net143),
    .TE_B(_0172_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1057_ (.A(\mux_bottom_track_9.INVTX1_6_.out ),
    .TE_B(_0173_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1058_ (.A(\mux_right_track_2.INVTX1_4_.out ),
    .TE_B(_0174_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1059_ (.A(\mux_right_track_12.INVTX1_1_.out ),
    .TE_B(_0175_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1060_ (.A(\mux_top_track_8.INVTX1_1_.out ),
    .TE_B(_0176_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1061_ (.A(\mux_bottom_track_9.INVTX1_3_.out ),
    .TE_B(_0177_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1062_ (.A(\mux_bottom_track_9.INVTX1_4_.out ),
    .TE_B(_0178_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1063_ (.A(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out ),
    .TE_B(_0179_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1064_ (.A(\mux_bottom_track_9.INVTX1_5_.out ),
    .TE_B(_0180_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1065_ (.A(\mux_top_track_8.INVTX1_0_.out ),
    .TE_B(_0181_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1066_ (.A(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out ),
    .TE_B(_0182_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1067_ (.A(\mux_right_track_24.INVTX1_2_.out ),
    .TE_B(_0183_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1068_ (.A(net144),
    .TE_B(_0184_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_8 _1069_ (.A(\mux_bottom_track_1.INVTX1_6_.out ),
    .TE_B(_0185_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_8 _1070_ (.A(\mux_right_track_4.INVTX1_4_.out ),
    .TE_B(_0186_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_8 _1071_ (.A(\mux_right_track_14.INVTX1_1_.out ),
    .TE_B(_0187_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_8 _1072_ (.A(\mux_top_track_16.INVTX1_1_.out ),
    .TE_B(_0188_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_8 _1073_ (.A(\mux_bottom_track_1.INVTX1_3_.out ),
    .TE_B(_0189_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_8 _1074_ (.A(\mux_bottom_track_1.INVTX1_4_.out ),
    .TE_B(_0190_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1075_ (.A(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out ),
    .TE_B(_0191_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_8 _1076_ (.A(\mux_bottom_track_1.INVTX1_5_.out ),
    .TE_B(_0192_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_8 _1077_ (.A(\mux_top_track_16.INVTX1_0_.out ),
    .TE_B(_0193_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1078_ (.A(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out ),
    .TE_B(_0194_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1079_ (.A(\mux_bottom_track_1.INVTX1_8_.out ),
    .TE_B(_0195_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1080_ (.A(net145),
    .TE_B(_0196_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1081_ (.A(\mux_bottom_track_1.INVTX1_5_.out ),
    .TE_B(_0197_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1082_ (.A(\mux_bottom_track_1.INVTX1_6_.out ),
    .TE_B(_0198_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1083_ (.A(\mux_bottom_track_1.INVTX1_7_.out ),
    .TE_B(_0199_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1084_ (.A(\mux_bottom_track_1.INVTX1_1_.out ),
    .TE_B(_0200_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1085_ (.A(\mux_bottom_track_1.INVTX1_2_.out ),
    .TE_B(_0201_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1086_ (.A(\mux_bottom_track_1.INVTX1_3_.out ),
    .TE_B(_0202_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1087_ (.A(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out ),
    .TE_B(_0203_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1088_ (.A(\mux_bottom_track_1.INVTX1_4_.out ),
    .TE_B(_0204_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1089_ (.A(\mux_bottom_track_1.INVTX1_0_.out ),
    .TE_B(_0205_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1090_ (.A(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out ),
    .TE_B(_0206_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1091_ (.A(\mux_bottom_track_9.INVTX1_8_.out ),
    .TE_B(_0207_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1092_ (.A(net146),
    .TE_B(_0208_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1093_ (.A(\mux_bottom_track_9.INVTX1_5_.out ),
    .TE_B(_0209_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1094_ (.A(\mux_bottom_track_9.INVTX1_6_.out ),
    .TE_B(_0210_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1095_ (.A(\mux_bottom_track_9.INVTX1_7_.out ),
    .TE_B(_0211_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1096_ (.A(\mux_bottom_track_9.INVTX1_1_.out ),
    .TE_B(_0212_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1097_ (.A(\mux_bottom_track_9.INVTX1_2_.out ),
    .TE_B(_0213_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1098_ (.A(\mux_bottom_track_9.INVTX1_3_.out ),
    .TE_B(_0214_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1099_ (.A(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out ),
    .TE_B(_0215_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1100_ (.A(\mux_bottom_track_9.INVTX1_4_.out ),
    .TE_B(_0216_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1101_ (.A(\mux_bottom_track_9.INVTX1_0_.out ),
    .TE_B(_0217_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1102_ (.A(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out ),
    .TE_B(_0218_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1103_ (.A(\mux_bottom_track_17.INVTX1_8_.out ),
    .TE_B(_0219_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1104_ (.A(net147),
    .TE_B(_0220_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1105_ (.A(\mux_bottom_track_17.INVTX1_5_.out ),
    .TE_B(_0221_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1106_ (.A(\mux_bottom_track_17.INVTX1_6_.out ),
    .TE_B(_0222_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1107_ (.A(\mux_bottom_track_17.INVTX1_7_.out ),
    .TE_B(_0223_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1108_ (.A(\mux_bottom_track_17.INVTX1_1_.out ),
    .TE_B(_0224_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1109_ (.A(\mux_bottom_track_17.INVTX1_2_.out ),
    .TE_B(_0225_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1110_ (.A(\mux_bottom_track_17.INVTX1_3_.out ),
    .TE_B(_0226_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1111_ (.A(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out ),
    .TE_B(_0227_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1112_ (.A(\mux_bottom_track_17.INVTX1_4_.out ),
    .TE_B(_0228_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1113_ (.A(\mux_bottom_track_17.INVTX1_0_.out ),
    .TE_B(_0229_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1114_ (.A(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out ),
    .TE_B(_0230_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1115_ (.A(\mux_bottom_track_25.INVTX1_8_.out ),
    .TE_B(_0231_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1116_ (.A(net148),
    .TE_B(_0232_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1117_ (.A(\mux_bottom_track_25.INVTX1_5_.out ),
    .TE_B(_0233_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1118_ (.A(\mux_bottom_track_25.INVTX1_6_.out ),
    .TE_B(_0234_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1119_ (.A(\mux_bottom_track_25.INVTX1_7_.out ),
    .TE_B(_0235_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1120_ (.A(\mux_bottom_track_25.INVTX1_1_.out ),
    .TE_B(_0236_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1121_ (.A(\mux_bottom_track_25.INVTX1_2_.out ),
    .TE_B(_0237_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1122_ (.A(\mux_bottom_track_25.INVTX1_3_.out ),
    .TE_B(_0238_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1123_ (.A(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out ),
    .TE_B(_0239_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1124_ (.A(\mux_bottom_track_25.INVTX1_4_.out ),
    .TE_B(_0240_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1125_ (.A(\mux_bottom_track_25.INVTX1_0_.out ),
    .TE_B(_0241_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1126_ (.A(\mux_top_track_24.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_0242_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _1127_ (.A(\mux_top_track_24.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_0243_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _1128_ (.A(\mux_right_track_26.INVTX1_1_.out ),
    .TE_B(_0244_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1129_ (.A(net149),
    .TE_B(_0245_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1130_ (.A(\mux_bottom_track_33.INVTX1_4_.out ),
    .TE_B(_0246_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1131_ (.A(\mux_right_track_6.INVTX1_3_.out ),
    .TE_B(_0247_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1132_ (.A(\mux_top_track_24.INVTX1_1_.out ),
    .TE_B(_0248_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1133_ (.A(\mux_bottom_track_33.INVTX1_2_.out ),
    .TE_B(_0249_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1134_ (.A(\mux_top_track_24.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_0250_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _1135_ (.A(\mux_right_track_16.INVTX1_1_.out ),
    .TE_B(_0251_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1136_ (.A(\mux_bottom_track_33.INVTX1_3_.out ),
    .TE_B(_0252_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1137_ (.A(\mux_top_track_24.INVTX1_0_.out ),
    .TE_B(_0253_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1138_ (.A(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_0254_),
    .Z(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _1139_ (.A(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_0255_),
    .Z(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _1140_ (.A(\mux_right_track_18.INVTX1_2_.out ),
    .TE_B(_0256_),
    .Z(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1141_ (.A(net150),
    .TE_B(_0257_),
    .Z(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1142_ (.A(\mux_bottom_track_25.INVTX1_5_.out ),
    .TE_B(_0258_),
    .Z(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1143_ (.A(\mux_bottom_track_25.INVTX1_6_.out ),
    .TE_B(_0259_),
    .Z(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1144_ (.A(\mux_top_track_32.INVTX1_1_.out ),
    .TE_B(_0260_),
    .Z(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1145_ (.A(\mux_bottom_track_25.INVTX1_3_.out ),
    .TE_B(_0261_),
    .Z(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1146_ (.A(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_0262_),
    .Z(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _1147_ (.A(\mux_right_track_8.INVTX1_2_.out ),
    .TE_B(_0263_),
    .Z(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1148_ (.A(\mux_bottom_track_25.INVTX1_4_.out ),
    .TE_B(_0264_),
    .Z(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1149_ (.A(\mux_top_track_32.INVTX1_0_.out ),
    .TE_B(_0265_),
    .Z(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1150_ (.A(\mux_right_track_0.INVTX1_3_.out ),
    .TE_B(_0266_),
    .Z(\mux_right_track_0.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1151_ (.A(net151),
    .TE_B(_0267_),
    .Z(\mux_right_track_0.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1152_ (.A(\mux_right_track_0.INVTX1_1_.out ),
    .TE_B(_0268_),
    .Z(\mux_right_track_0.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1153_ (.A(\mux_right_track_0.INVTX1_2_.out ),
    .TE_B(_0269_),
    .Z(\mux_right_track_0.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1154_ (.A(\mux_right_track_0.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_0270_),
    .Z(\mux_right_track_0.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1155_ (.A(\mux_bottom_track_1.INVTX1_0_.out ),
    .TE_B(_0271_),
    .Z(\mux_right_track_0.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1156_ (.A(\mux_right_track_6.INVTX1_3_.out ),
    .TE_B(_0272_),
    .Z(\mux_right_track_6.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1157_ (.A(net152),
    .TE_B(_0273_),
    .Z(\mux_right_track_6.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1158_ (.A(\mux_right_track_6.INVTX1_1_.out ),
    .TE_B(_0274_),
    .Z(\mux_right_track_6.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1159_ (.A(\mux_right_track_24.INVTX1_1_.out ),
    .TE_B(_0275_),
    .Z(\mux_right_track_6.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1160_ (.A(\mux_right_track_6.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_0276_),
    .Z(\mux_right_track_6.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1161_ (.A(\mux_bottom_track_25.INVTX1_0_.out ),
    .TE_B(_0277_),
    .Z(\mux_right_track_6.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1162_ (.A(\mux_right_track_2.INVTX1_4_.out ),
    .TE_B(_0278_),
    .Z(\mux_right_track_2.mux_2level_tapbuf_basis_input2_mem2_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1163_ (.A(\mux_right_track_2.mux_2level_tapbuf_basis_input2_mem2_0_out ),
    .TE_B(_0279_),
    .Z(\mux_right_track_2.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1164_ (.A(net153),
    .TE_B(_0280_),
    .Z(\mux_right_track_2.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1165_ (.A(\mux_right_track_2.INVTX1_1_.out ),
    .TE_B(_0281_),
    .Z(\mux_right_track_2.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1166_ (.A(\mux_right_track_0.INVTX1_2_.out ),
    .TE_B(_0282_),
    .Z(\mux_right_track_2.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1167_ (.A(\mux_right_track_2.INVTX1_3_.out ),
    .TE_B(_0283_),
    .Z(\mux_right_track_2.mux_2level_tapbuf_basis_input2_mem2_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1168_ (.A(\mux_right_track_2.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_0284_),
    .Z(\mux_right_track_2.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1169_ (.A(\mux_bottom_track_9.INVTX1_0_.out ),
    .TE_B(_0285_),
    .Z(\mux_right_track_2.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1170_ (.A(\mux_right_track_4.INVTX1_4_.out ),
    .TE_B(_0286_),
    .Z(\mux_right_track_4.mux_2level_tapbuf_basis_input2_mem2_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1171_ (.A(\mux_right_track_4.mux_2level_tapbuf_basis_input2_mem2_0_out ),
    .TE_B(_0287_),
    .Z(\mux_right_track_4.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1172_ (.A(net154),
    .TE_B(_0288_),
    .Z(\mux_right_track_4.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1173_ (.A(\mux_right_track_4.INVTX1_1_.out ),
    .TE_B(_0289_),
    .Z(\mux_right_track_4.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1174_ (.A(\mux_right_track_2.INVTX1_3_.out ),
    .TE_B(_0290_),
    .Z(\mux_right_track_4.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1175_ (.A(\mux_right_track_24.INVTX1_1_.out ),
    .TE_B(_0291_),
    .Z(\mux_right_track_4.mux_2level_tapbuf_basis_input2_mem2_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1176_ (.A(\mux_right_track_4.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_0292_),
    .Z(\mux_right_track_4.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1177_ (.A(\mux_bottom_track_17.INVTX1_0_.out ),
    .TE_B(_0293_),
    .Z(\mux_right_track_4.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1178_ (.A(\mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0294_),
    .Z(\mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1179_ (.A(net155),
    .TE_B(_0295_),
    .Z(\mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1180_ (.A(\mux_right_track_8.INVTX1_1_.out ),
    .TE_B(_0296_),
    .Z(\mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1181_ (.A(\mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0297_),
    .Z(\mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1182_ (.A(\mux_right_track_8.INVTX1_2_.out ),
    .TE_B(_0298_),
    .Z(\mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1183_ (.A(\mux_bottom_track_33.INVTX1_0_.out ),
    .TE_B(_0299_),
    .Z(\mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1184_ (.A(\mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0300_),
    .Z(\mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1185_ (.A(net156),
    .TE_B(_0301_),
    .Z(\mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1186_ (.A(\mux_right_track_10.INVTX1_1_.out ),
    .TE_B(_0302_),
    .Z(\mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1187_ (.A(\mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0303_),
    .Z(\mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1188_ (.A(\mux_right_track_10.INVTX1_2_.out ),
    .TE_B(_0304_),
    .Z(\mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1189_ (.A(\mux_bottom_track_1.INVTX1_1_.out ),
    .TE_B(_0305_),
    .Z(\mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1190_ (.A(\mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0306_),
    .Z(\mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1191_ (.A(net157),
    .TE_B(_0307_),
    .Z(\mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1192_ (.A(\mux_right_track_0.INVTX1_1_.out ),
    .TE_B(_0308_),
    .Z(\mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1193_ (.A(\mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0309_),
    .Z(\mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1194_ (.A(\mux_right_track_18.INVTX1_2_.out ),
    .TE_B(_0310_),
    .Z(\mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1195_ (.A(\mux_bottom_track_33.INVTX1_1_.out ),
    .TE_B(_0311_),
    .Z(\mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1196_ (.A(\mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0312_),
    .Z(\mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1197_ (.A(net158),
    .TE_B(_0313_),
    .Z(\mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1198_ (.A(\mux_right_track_0.INVTX1_2_.out ),
    .TE_B(_0314_),
    .Z(\mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1199_ (.A(\mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0315_),
    .Z(\mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1200_ (.A(\mux_right_track_20.INVTX1_2_.out ),
    .TE_B(_0316_),
    .Z(\mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1201_ (.A(\mux_bottom_track_1.INVTX1_2_.out ),
    .TE_B(_0317_),
    .Z(\mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1202_ (.A(\mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0318_),
    .Z(\mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1203_ (.A(net159),
    .TE_B(_0319_),
    .Z(\mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1204_ (.A(\mux_right_track_2.INVTX1_3_.out ),
    .TE_B(_0320_),
    .Z(\mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1205_ (.A(\mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0321_),
    .Z(\mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1206_ (.A(\mux_right_track_22.INVTX1_2_.out ),
    .TE_B(_0322_),
    .Z(\mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1207_ (.A(\mux_bottom_track_9.INVTX1_2_.out ),
    .TE_B(_0323_),
    .Z(\mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1208_ (.A(\mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0324_),
    .Z(\mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1209_ (.A(net160),
    .TE_B(_0325_),
    .Z(\mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1210_ (.A(\mux_right_track_24.INVTX1_1_.out ),
    .TE_B(_0326_),
    .Z(\mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1211_ (.A(\mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0327_),
    .Z(\mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1212_ (.A(\mux_right_track_24.INVTX1_2_.out ),
    .TE_B(_0328_),
    .Z(\mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1213_ (.A(\mux_bottom_track_17.INVTX1_2_.out ),
    .TE_B(_0329_),
    .Z(\mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1214_ (.A(\mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0330_),
    .Z(\mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1215_ (.A(net161),
    .TE_B(_0331_),
    .Z(\mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1216_ (.A(\mux_right_track_26.INVTX1_1_.out ),
    .TE_B(_0332_),
    .Z(\mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1217_ (.A(\mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0333_),
    .Z(\mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1218_ (.A(\mux_right_track_26.INVTX1_2_.out ),
    .TE_B(_0334_),
    .Z(\mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1219_ (.A(\mux_bottom_track_25.INVTX1_2_.out ),
    .TE_B(_0335_),
    .Z(\mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1220_ (.A(net162),
    .TE_B(_0336_),
    .Z(\mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1221_ (.A(\mux_right_track_12.INVTX1_1_.out ),
    .TE_B(_0337_),
    .Z(\mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1222_ (.A(\mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0338_),
    .Z(\mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1223_ (.A(\mux_bottom_track_9.INVTX1_1_.out ),
    .TE_B(_0339_),
    .Z(\mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1224_ (.A(net163),
    .TE_B(_0340_),
    .Z(\mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1225_ (.A(\mux_right_track_14.INVTX1_1_.out ),
    .TE_B(_0341_),
    .Z(\mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1226_ (.A(\mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0342_),
    .Z(\mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1227_ (.A(\mux_bottom_track_17.INVTX1_1_.out ),
    .TE_B(_0343_),
    .Z(\mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1228_ (.A(net164),
    .TE_B(_0344_),
    .Z(\mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1229_ (.A(\mux_right_track_16.INVTX1_1_.out ),
    .TE_B(_0345_),
    .Z(\mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1230_ (.A(\mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0346_),
    .Z(\mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1231_ (.A(\mux_bottom_track_25.INVTX1_1_.out ),
    .TE_B(_0347_),
    .Z(\mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1232_ (.A(net165),
    .TE_B(_0348_),
    .Z(\mux_bottom_track_33.mux_2level_tapbuf_basis_input2_mem2_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1233_ (.A(\mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_0349_),
    .Z(\mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1234_ (.A(\mux_bottom_track_33.mux_2level_tapbuf_basis_input2_mem2_0_out ),
    .TE_B(_0350_),
    .Z(\mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1235_ (.A(\mux_bottom_track_33.INVTX1_4_.out ),
    .TE_B(_0351_),
    .Z(\mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1236_ (.A(\mux_bottom_track_33.INVTX1_5_.out ),
    .TE_B(_0352_),
    .Z(\mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1237_ (.A(\mux_bottom_track_33.INVTX1_1_.out ),
    .TE_B(_0353_),
    .Z(\mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1238_ (.A(\mux_bottom_track_33.INVTX1_2_.out ),
    .TE_B(_0354_),
    .Z(\mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1239_ (.A(\mux_bottom_track_33.INVTX1_6_.out ),
    .TE_B(_0355_),
    .Z(\mux_bottom_track_33.mux_2level_tapbuf_basis_input2_mem2_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1240_ (.A(\mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_0356_),
    .Z(\mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1241_ (.A(\mux_bottom_track_33.INVTX1_3_.out ),
    .TE_B(_0357_),
    .Z(\mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1242_ (.A(\mux_bottom_track_33.INVTX1_0_.out ),
    .TE_B(_0358_),
    .Z(\mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_),
    .X(net10));
 sky130_fd_sc_hd__dlymetal6s2s_1 input11 (.A(ccff_head),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(chanx_right_in[0]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(chanx_right_in[10]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(chanx_right_in[11]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(chanx_right_in[12]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(chanx_right_in[13]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(chanx_right_in[14]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(chanx_right_in[15]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(chanx_right_in[16]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(chanx_right_in[17]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(chanx_right_in[18]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(chanx_right_in[1]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(chanx_right_in[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(chanx_right_in[3]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(chanx_right_in[4]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(chanx_right_in[5]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(chanx_right_in[6]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(chanx_right_in[7]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(chanx_right_in[8]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(chanx_right_in[9]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(chany_bottom_in[0]),
    .X(net31));
 sky130_fd_sc_hd__dlymetal6s2s_1 input32 (.A(chany_bottom_in[10]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(chany_bottom_in[11]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(chany_bottom_in[12]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(chany_bottom_in[13]),
    .X(net35));
 sky130_fd_sc_hd__dlymetal6s2s_1 input36 (.A(chany_bottom_in[14]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(chany_bottom_in[15]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(chany_bottom_in[16]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(chany_bottom_in[17]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(chany_bottom_in[18]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(chany_bottom_in[1]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(chany_bottom_in[2]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(chany_bottom_in[3]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(chany_bottom_in[4]),
    .X(net44));
 sky130_fd_sc_hd__dlymetal6s2s_1 input45 (.A(chany_bottom_in[5]),
    .X(net45));
 sky130_fd_sc_hd__dlymetal6s2s_1 input46 (.A(chany_bottom_in[6]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(chany_bottom_in[7]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(chany_bottom_in[8]),
    .X(net48));
 sky130_fd_sc_hd__dlymetal6s2s_1 input49 (.A(chany_bottom_in[9]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(chany_top_in[0]),
    .X(net50));
 sky130_fd_sc_hd__dlymetal6s2s_1 input51 (.A(chany_top_in[10]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(chany_top_in[11]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(chany_top_in[12]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(chany_top_in[13]),
    .X(net54));
 sky130_fd_sc_hd__dlymetal6s2s_1 input55 (.A(chany_top_in[14]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(chany_top_in[15]),
    .X(net56));
 sky130_fd_sc_hd__dlymetal6s2s_1 input57 (.A(chany_top_in[16]),
    .X(net57));
 sky130_fd_sc_hd__dlymetal6s2s_1 input58 (.A(chany_top_in[17]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(chany_top_in[18]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(chany_top_in[1]),
    .X(net60));
 sky130_fd_sc_hd__dlymetal6s2s_1 input61 (.A(chany_top_in[2]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(chany_top_in[3]),
    .X(net62));
 sky130_fd_sc_hd__dlymetal6s2s_1 input63 (.A(chany_top_in[4]),
    .X(net63));
 sky130_fd_sc_hd__dlymetal6s2s_1 input64 (.A(chany_top_in[5]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 input65 (.A(chany_top_in[6]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(chany_top_in[7]),
    .X(net66));
 sky130_fd_sc_hd__dlymetal6s2s_1 input67 (.A(chany_top_in[8]),
    .X(net67));
 sky130_fd_sc_hd__dlymetal6s2s_1 input68 (.A(chany_top_in[9]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(pReset),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_2 input72 (.A(right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 input73 (.A(right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 input74 (.A(top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 input75 (.A(top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 input76 (.A(top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 input78 (.A(top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 input79 (.A(top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 input80 (.A(top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 input81 (.A(top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 input82 (.A(top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 input83 (.A(top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_),
    .X(net83));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(ccff_tail));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(chanx_right_out[0]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(chanx_right_out[10]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(chanx_right_out[11]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(chanx_right_out[12]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(chanx_right_out[13]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(chanx_right_out[14]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .X(chanx_right_out[15]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(chanx_right_out[16]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net93),
    .X(chanx_right_out[17]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net94),
    .X(chanx_right_out[18]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(chanx_right_out[1]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(chanx_right_out[2]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net97),
    .X(chanx_right_out[3]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(chanx_right_out[4]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(chanx_right_out[5]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .X(chanx_right_out[6]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(chanx_right_out[7]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(chanx_right_out[8]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(chanx_right_out[9]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(chany_bottom_out[0]));
 sky130_fd_sc_hd__buf_2 output105 (.A(net105),
    .X(chany_bottom_out[10]));
 sky130_fd_sc_hd__buf_2 output106 (.A(net106),
    .X(chany_bottom_out[11]));
 sky130_fd_sc_hd__buf_2 output107 (.A(net107),
    .X(chany_bottom_out[12]));
 sky130_fd_sc_hd__buf_2 output108 (.A(net108),
    .X(chany_bottom_out[13]));
 sky130_fd_sc_hd__buf_2 output109 (.A(net109),
    .X(chany_bottom_out[14]));
 sky130_fd_sc_hd__buf_2 output110 (.A(net110),
    .X(chany_bottom_out[15]));
 sky130_fd_sc_hd__buf_2 output111 (.A(net111),
    .X(chany_bottom_out[16]));
 sky130_fd_sc_hd__buf_2 output112 (.A(net112),
    .X(chany_bottom_out[17]));
 sky130_fd_sc_hd__buf_2 output113 (.A(net113),
    .X(chany_bottom_out[18]));
 sky130_fd_sc_hd__buf_2 output114 (.A(net114),
    .X(chany_bottom_out[1]));
 sky130_fd_sc_hd__buf_2 output115 (.A(net115),
    .X(chany_bottom_out[2]));
 sky130_fd_sc_hd__buf_2 output116 (.A(net116),
    .X(chany_bottom_out[3]));
 sky130_fd_sc_hd__buf_2 output117 (.A(net117),
    .X(chany_bottom_out[4]));
 sky130_fd_sc_hd__buf_2 output118 (.A(net118),
    .X(chany_bottom_out[5]));
 sky130_fd_sc_hd__buf_2 output119 (.A(net119),
    .X(chany_bottom_out[6]));
 sky130_fd_sc_hd__buf_2 output120 (.A(net120),
    .X(chany_bottom_out[7]));
 sky130_fd_sc_hd__buf_2 output121 (.A(net121),
    .X(chany_bottom_out[8]));
 sky130_fd_sc_hd__buf_2 output122 (.A(net122),
    .X(chany_bottom_out[9]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net123),
    .X(chany_top_out[0]));
 sky130_fd_sc_hd__buf_2 output124 (.A(net124),
    .X(chany_top_out[10]));
 sky130_fd_sc_hd__buf_2 output125 (.A(net125),
    .X(chany_top_out[11]));
 sky130_fd_sc_hd__buf_2 output126 (.A(net126),
    .X(chany_top_out[12]));
 sky130_fd_sc_hd__buf_2 output127 (.A(net127),
    .X(chany_top_out[13]));
 sky130_fd_sc_hd__buf_2 output128 (.A(net128),
    .X(chany_top_out[14]));
 sky130_fd_sc_hd__buf_2 output129 (.A(net129),
    .X(chany_top_out[15]));
 sky130_fd_sc_hd__buf_2 output130 (.A(net130),
    .X(chany_top_out[16]));
 sky130_fd_sc_hd__buf_2 output131 (.A(net131),
    .X(chany_top_out[17]));
 sky130_fd_sc_hd__buf_2 output132 (.A(net132),
    .X(chany_top_out[18]));
 sky130_fd_sc_hd__buf_2 output133 (.A(net133),
    .X(chany_top_out[1]));
 sky130_fd_sc_hd__buf_2 output134 (.A(net134),
    .X(chany_top_out[2]));
 sky130_fd_sc_hd__buf_2 output135 (.A(net135),
    .X(chany_top_out[3]));
 sky130_fd_sc_hd__buf_2 output136 (.A(net136),
    .X(chany_top_out[4]));
 sky130_fd_sc_hd__buf_2 output137 (.A(net137),
    .X(chany_top_out[5]));
 sky130_fd_sc_hd__buf_2 output138 (.A(net138),
    .X(chany_top_out[6]));
 sky130_fd_sc_hd__buf_2 output139 (.A(net139),
    .X(chany_top_out[7]));
 sky130_fd_sc_hd__buf_2 output140 (.A(net140),
    .X(chany_top_out[8]));
 sky130_fd_sc_hd__buf_2 output141 (.A(net141),
    .X(chany_top_out[9]));
 sky130_fd_sc_hd__conb_1 _1044__142 (.HI(net142));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_0_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_1_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_2_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_3_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_4_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_5_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_6_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_7_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_8_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_9_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_10_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_11_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_12_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_13_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_14_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_15_0_prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\mem_right_track_10.DFFR_0_.Q ));
 sky130_fd_sc_hd__decap_6 FILLER_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_405 ();
endmodule

