magic
tech sky130A
magscale 1 2
timestamp 1674175246
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 14 1640 39362 37584
<< metal2 >>
rect 18 39200 74 39800
rect 1306 39200 1362 39800
rect 3238 39200 3294 39800
rect 4526 39200 4582 39800
rect 5814 39200 5870 39800
rect 7746 39200 7802 39800
rect 9034 39200 9090 39800
rect 10322 39200 10378 39800
rect 12254 39200 12310 39800
rect 13542 39200 13598 39800
rect 15474 39200 15530 39800
rect 16762 39200 16818 39800
rect 18050 39200 18106 39800
rect 19982 39200 20038 39800
rect 21270 39200 21326 39800
rect 22558 39200 22614 39800
rect 24490 39200 24546 39800
rect 25778 39200 25834 39800
rect 27710 39200 27766 39800
rect 28998 39200 29054 39800
rect 30286 39200 30342 39800
rect 32218 39200 32274 39800
rect 33506 39200 33562 39800
rect 34794 39200 34850 39800
rect 36726 39200 36782 39800
rect 38014 39200 38070 39800
rect 39302 39200 39358 39800
rect 18 200 74 800
rect 1306 200 1362 800
rect 2594 200 2650 800
rect 4526 200 4582 800
rect 5814 200 5870 800
rect 7102 200 7158 800
rect 9034 200 9090 800
rect 10322 200 10378 800
rect 11610 200 11666 800
rect 13542 200 13598 800
rect 14830 200 14886 800
rect 16762 200 16818 800
rect 18050 200 18106 800
rect 19338 200 19394 800
rect 21270 200 21326 800
rect 22558 200 22614 800
rect 23846 200 23902 800
rect 25778 200 25834 800
rect 27066 200 27122 800
rect 28998 200 29054 800
rect 30286 200 30342 800
rect 31574 200 31630 800
rect 33506 200 33562 800
rect 34794 200 34850 800
rect 36082 200 36138 800
rect 38014 200 38070 800
rect 39302 200 39358 800
<< obsm2 >>
rect 130 39144 1250 39200
rect 1418 39144 3182 39200
rect 3350 39144 4470 39200
rect 4638 39144 5758 39200
rect 5926 39144 7690 39200
rect 7858 39144 8978 39200
rect 9146 39144 10266 39200
rect 10434 39144 12198 39200
rect 12366 39144 13486 39200
rect 13654 39144 15418 39200
rect 15586 39144 16706 39200
rect 16874 39144 17994 39200
rect 18162 39144 19926 39200
rect 20094 39144 21214 39200
rect 21382 39144 22502 39200
rect 22670 39144 24434 39200
rect 24602 39144 25722 39200
rect 25890 39144 27654 39200
rect 27822 39144 28942 39200
rect 29110 39144 30230 39200
rect 30398 39144 32162 39200
rect 32330 39144 33450 39200
rect 33618 39144 34738 39200
rect 34906 39144 36670 39200
rect 36838 39144 37958 39200
rect 38126 39144 39246 39200
rect 20 856 39356 39144
rect 130 734 1250 856
rect 1418 734 2538 856
rect 2706 734 4470 856
rect 4638 734 5758 856
rect 5926 734 7046 856
rect 7214 734 8978 856
rect 9146 734 10266 856
rect 10434 734 11554 856
rect 11722 734 13486 856
rect 13654 734 14774 856
rect 14942 734 16706 856
rect 16874 734 17994 856
rect 18162 734 19282 856
rect 19450 734 21214 856
rect 21382 734 22502 856
rect 22670 734 23790 856
rect 23958 734 25722 856
rect 25890 734 27010 856
rect 27178 734 28942 856
rect 29110 734 30230 856
rect 30398 734 31518 856
rect 31686 734 33450 856
rect 33618 734 34738 856
rect 34906 734 36026 856
rect 36194 734 37958 856
rect 38126 734 39246 856
<< metal3 >>
rect 200 38088 800 38208
rect 39200 38088 39800 38208
rect 200 36728 800 36848
rect 39200 36728 39800 36848
rect 200 35368 800 35488
rect 39200 34688 39800 34808
rect 200 33328 800 33448
rect 39200 33328 39800 33448
rect 200 31968 800 32088
rect 39200 31968 39800 32088
rect 200 30608 800 30728
rect 39200 29928 39800 30048
rect 200 28568 800 28688
rect 39200 28568 39800 28688
rect 200 27208 800 27328
rect 39200 27208 39800 27328
rect 200 25168 800 25288
rect 39200 25168 39800 25288
rect 200 23808 800 23928
rect 39200 23808 39800 23928
rect 200 22448 800 22568
rect 39200 21768 39800 21888
rect 200 20408 800 20528
rect 39200 20408 39800 20528
rect 200 19048 800 19168
rect 39200 19048 39800 19168
rect 200 17688 800 17808
rect 39200 17008 39800 17128
rect 200 15648 800 15768
rect 39200 15648 39800 15768
rect 200 14288 800 14408
rect 39200 14288 39800 14408
rect 200 12248 800 12368
rect 39200 12248 39800 12368
rect 200 10888 800 11008
rect 39200 10888 39800 11008
rect 200 9528 800 9648
rect 39200 8848 39800 8968
rect 200 7488 800 7608
rect 39200 7488 39800 7608
rect 200 6128 800 6248
rect 39200 6128 39800 6248
rect 200 4768 800 4888
rect 39200 4088 39800 4208
rect 200 2728 800 2848
rect 39200 2728 39800 2848
rect 200 1368 800 1488
rect 39200 1368 39800 1488
<< obsm3 >>
rect 880 38008 39120 38181
rect 800 36928 39200 38008
rect 880 36648 39120 36928
rect 800 35568 39200 36648
rect 880 35288 39200 35568
rect 800 34888 39200 35288
rect 800 34608 39120 34888
rect 800 33528 39200 34608
rect 880 33248 39120 33528
rect 800 32168 39200 33248
rect 880 31888 39120 32168
rect 800 30808 39200 31888
rect 880 30528 39200 30808
rect 800 30128 39200 30528
rect 800 29848 39120 30128
rect 800 28768 39200 29848
rect 880 28488 39120 28768
rect 800 27408 39200 28488
rect 880 27128 39120 27408
rect 800 25368 39200 27128
rect 880 25088 39120 25368
rect 800 24008 39200 25088
rect 880 23728 39120 24008
rect 800 22648 39200 23728
rect 880 22368 39200 22648
rect 800 21968 39200 22368
rect 800 21688 39120 21968
rect 800 20608 39200 21688
rect 880 20328 39120 20608
rect 800 19248 39200 20328
rect 880 18968 39120 19248
rect 800 17888 39200 18968
rect 880 17608 39200 17888
rect 800 17208 39200 17608
rect 800 16928 39120 17208
rect 800 15848 39200 16928
rect 880 15568 39120 15848
rect 800 14488 39200 15568
rect 880 14208 39120 14488
rect 800 12448 39200 14208
rect 880 12168 39120 12448
rect 800 11088 39200 12168
rect 880 10808 39120 11088
rect 800 9728 39200 10808
rect 880 9448 39200 9728
rect 800 9048 39200 9448
rect 800 8768 39120 9048
rect 800 7688 39200 8768
rect 880 7408 39120 7688
rect 800 6328 39200 7408
rect 880 6048 39120 6328
rect 800 4968 39200 6048
rect 880 4688 39200 4968
rect 800 4288 39200 4688
rect 800 4008 39120 4288
rect 800 2928 39200 4008
rect 880 2648 39120 2928
rect 800 1568 39200 2648
rect 880 1395 39120 1568
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< obsm4 >>
rect 3187 2347 4128 22677
rect 4608 2347 19445 22677
<< labels >>
rlabel metal3 s 39200 6128 39800 6248 6 ccff_head
port 1 nsew signal input
rlabel metal3 s 39200 33328 39800 33448 6 ccff_tail
port 2 nsew signal output
rlabel metal2 s 22558 39200 22614 39800 6 chanx_left_in[0]
port 3 nsew signal input
rlabel metal3 s 39200 38088 39800 38208 6 chanx_left_in[10]
port 4 nsew signal input
rlabel metal3 s 200 12248 800 12368 6 chanx_left_in[11]
port 5 nsew signal input
rlabel metal2 s 34794 200 34850 800 6 chanx_left_in[12]
port 6 nsew signal input
rlabel metal3 s 200 36728 800 36848 6 chanx_left_in[13]
port 7 nsew signal input
rlabel metal2 s 38014 39200 38070 39800 6 chanx_left_in[14]
port 8 nsew signal input
rlabel metal2 s 28998 200 29054 800 6 chanx_left_in[15]
port 9 nsew signal input
rlabel metal3 s 200 7488 800 7608 6 chanx_left_in[16]
port 10 nsew signal input
rlabel metal3 s 200 30608 800 30728 6 chanx_left_in[17]
port 11 nsew signal input
rlabel metal2 s 10322 200 10378 800 6 chanx_left_in[18]
port 12 nsew signal input
rlabel metal3 s 200 38088 800 38208 6 chanx_left_in[1]
port 13 nsew signal input
rlabel metal2 s 4526 200 4582 800 6 chanx_left_in[2]
port 14 nsew signal input
rlabel metal3 s 200 20408 800 20528 6 chanx_left_in[3]
port 15 nsew signal input
rlabel metal3 s 200 17688 800 17808 6 chanx_left_in[4]
port 16 nsew signal input
rlabel metal3 s 39200 28568 39800 28688 6 chanx_left_in[5]
port 17 nsew signal input
rlabel metal2 s 18050 39200 18106 39800 6 chanx_left_in[6]
port 18 nsew signal input
rlabel metal2 s 33506 200 33562 800 6 chanx_left_in[7]
port 19 nsew signal input
rlabel metal3 s 200 25168 800 25288 6 chanx_left_in[8]
port 20 nsew signal input
rlabel metal3 s 200 31968 800 32088 6 chanx_left_in[9]
port 21 nsew signal input
rlabel metal3 s 200 27208 800 27328 6 chanx_left_out[0]
port 22 nsew signal output
rlabel metal2 s 22558 200 22614 800 6 chanx_left_out[10]
port 23 nsew signal output
rlabel metal2 s 14830 200 14886 800 6 chanx_left_out[11]
port 24 nsew signal output
rlabel metal2 s 39302 200 39358 800 6 chanx_left_out[12]
port 25 nsew signal output
rlabel metal3 s 200 1368 800 1488 6 chanx_left_out[13]
port 26 nsew signal output
rlabel metal3 s 39200 20408 39800 20528 6 chanx_left_out[14]
port 27 nsew signal output
rlabel metal2 s 24490 39200 24546 39800 6 chanx_left_out[15]
port 28 nsew signal output
rlabel metal2 s 13542 39200 13598 39800 6 chanx_left_out[16]
port 29 nsew signal output
rlabel metal3 s 39200 36728 39800 36848 6 chanx_left_out[17]
port 30 nsew signal output
rlabel metal2 s 16762 200 16818 800 6 chanx_left_out[18]
port 31 nsew signal output
rlabel metal3 s 200 15648 800 15768 6 chanx_left_out[1]
port 32 nsew signal output
rlabel metal3 s 39200 34688 39800 34808 6 chanx_left_out[2]
port 33 nsew signal output
rlabel metal2 s 15474 39200 15530 39800 6 chanx_left_out[3]
port 34 nsew signal output
rlabel metal3 s 39200 8848 39800 8968 6 chanx_left_out[4]
port 35 nsew signal output
rlabel metal3 s 39200 12248 39800 12368 6 chanx_left_out[5]
port 36 nsew signal output
rlabel metal2 s 16762 39200 16818 39800 6 chanx_left_out[6]
port 37 nsew signal output
rlabel metal2 s 10322 39200 10378 39800 6 chanx_left_out[7]
port 38 nsew signal output
rlabel metal2 s 25778 200 25834 800 6 chanx_left_out[8]
port 39 nsew signal output
rlabel metal2 s 9034 200 9090 800 6 chanx_left_out[9]
port 40 nsew signal output
rlabel metal3 s 39200 29928 39800 30048 6 chany_top_in[0]
port 41 nsew signal input
rlabel metal2 s 38014 200 38070 800 6 chany_top_in[10]
port 42 nsew signal input
rlabel metal3 s 39200 15648 39800 15768 6 chany_top_in[11]
port 43 nsew signal input
rlabel metal2 s 28998 39200 29054 39800 6 chany_top_in[12]
port 44 nsew signal input
rlabel metal2 s 12254 39200 12310 39800 6 chany_top_in[13]
port 45 nsew signal input
rlabel metal3 s 39200 1368 39800 1488 6 chany_top_in[14]
port 46 nsew signal input
rlabel metal3 s 39200 31968 39800 32088 6 chany_top_in[15]
port 47 nsew signal input
rlabel metal2 s 36726 39200 36782 39800 6 chany_top_in[16]
port 48 nsew signal input
rlabel metal2 s 21270 39200 21326 39800 6 chany_top_in[17]
port 49 nsew signal input
rlabel metal3 s 200 19048 800 19168 6 chany_top_in[18]
port 50 nsew signal input
rlabel metal3 s 39200 7488 39800 7608 6 chany_top_in[1]
port 51 nsew signal input
rlabel metal3 s 200 22448 800 22568 6 chany_top_in[2]
port 52 nsew signal input
rlabel metal3 s 200 2728 800 2848 6 chany_top_in[3]
port 53 nsew signal input
rlabel metal2 s 25778 39200 25834 39800 6 chany_top_in[4]
port 54 nsew signal input
rlabel metal3 s 200 28568 800 28688 6 chany_top_in[5]
port 55 nsew signal input
rlabel metal2 s 30286 200 30342 800 6 chany_top_in[6]
port 56 nsew signal input
rlabel metal2 s 33506 39200 33562 39800 6 chany_top_in[7]
port 57 nsew signal input
rlabel metal3 s 200 9528 800 9648 6 chany_top_in[8]
port 58 nsew signal input
rlabel metal2 s 2594 200 2650 800 6 chany_top_in[9]
port 59 nsew signal input
rlabel metal2 s 11610 200 11666 800 6 chany_top_out[0]
port 60 nsew signal output
rlabel metal2 s 36082 200 36138 800 6 chany_top_out[10]
port 61 nsew signal output
rlabel metal3 s 39200 17008 39800 17128 6 chany_top_out[11]
port 62 nsew signal output
rlabel metal3 s 39200 10888 39800 11008 6 chany_top_out[12]
port 63 nsew signal output
rlabel metal3 s 200 6128 800 6248 6 chany_top_out[13]
port 64 nsew signal output
rlabel metal3 s 200 33328 800 33448 6 chany_top_out[14]
port 65 nsew signal output
rlabel metal3 s 39200 2728 39800 2848 6 chany_top_out[15]
port 66 nsew signal output
rlabel metal2 s 4526 39200 4582 39800 6 chany_top_out[16]
port 67 nsew signal output
rlabel metal3 s 39200 14288 39800 14408 6 chany_top_out[17]
port 68 nsew signal output
rlabel metal3 s 39200 25168 39800 25288 6 chany_top_out[18]
port 69 nsew signal output
rlabel metal2 s 31574 200 31630 800 6 chany_top_out[1]
port 70 nsew signal output
rlabel metal3 s 39200 27208 39800 27328 6 chany_top_out[2]
port 71 nsew signal output
rlabel metal2 s 5814 39200 5870 39800 6 chany_top_out[3]
port 72 nsew signal output
rlabel metal3 s 200 23808 800 23928 6 chany_top_out[4]
port 73 nsew signal output
rlabel metal2 s 19338 200 19394 800 6 chany_top_out[5]
port 74 nsew signal output
rlabel metal2 s 18 200 74 800 6 chany_top_out[6]
port 75 nsew signal output
rlabel metal2 s 23846 200 23902 800 6 chany_top_out[7]
port 76 nsew signal output
rlabel metal2 s 7746 39200 7802 39800 6 chany_top_out[8]
port 77 nsew signal output
rlabel metal2 s 19982 39200 20038 39800 6 chany_top_out[9]
port 78 nsew signal output
rlabel metal3 s 200 4768 800 4888 6 left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 79 nsew signal input
rlabel metal2 s 18 39200 74 39800 6 left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 80 nsew signal input
rlabel metal2 s 5814 200 5870 800 6 left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 81 nsew signal input
rlabel metal2 s 1306 200 1362 800 6 left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 82 nsew signal input
rlabel metal2 s 34794 39200 34850 39800 6 left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_
port 83 nsew signal input
rlabel metal2 s 27710 39200 27766 39800 6 left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_
port 84 nsew signal input
rlabel metal2 s 18050 200 18106 800 6 left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_
port 85 nsew signal input
rlabel metal2 s 39302 39200 39358 39800 6 left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_
port 86 nsew signal input
rlabel metal3 s 39200 4088 39800 4208 6 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
port 87 nsew signal input
rlabel metal2 s 1306 39200 1362 39800 6 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
port 88 nsew signal input
rlabel metal3 s 39200 21768 39800 21888 6 pReset
port 89 nsew signal input
rlabel metal2 s 7102 200 7158 800 6 prog_clk
port 90 nsew signal input
rlabel metal2 s 13542 200 13598 800 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
port 91 nsew signal input
rlabel metal3 s 200 14288 800 14408 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
port 92 nsew signal input
rlabel metal3 s 39200 23808 39800 23928 6 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 93 nsew signal input
rlabel metal2 s 21270 200 21326 800 6 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
port 94 nsew signal input
rlabel metal2 s 32218 39200 32274 39800 6 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
port 95 nsew signal input
rlabel metal2 s 30286 39200 30342 39800 6 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
port 96 nsew signal input
rlabel metal2 s 3238 39200 3294 39800 6 top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_
port 97 nsew signal input
rlabel metal2 s 9034 39200 9090 39800 6 top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_
port 98 nsew signal input
rlabel metal2 s 27066 200 27122 800 6 top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_
port 99 nsew signal input
rlabel metal3 s 200 10888 800 11008 6 top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_
port 100 nsew signal input
rlabel metal3 s 200 35368 800 35488 6 vccd1
port 101 nsew signal bidirectional
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 101 nsew signal bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 101 nsew signal bidirectional
rlabel metal3 s 39200 19048 39800 19168 6 vssd1
port 102 nsew signal bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 102 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2203872
string GDS_FILE /home/baungarten/Proyectos_caravel/FPGA_3/openlane/sb_4__0_/runs/23_01_19_18_39/results/signoff/sb_4__0_.magic.gds
string GDS_START 138498
<< end >>

