magic
tech sky130A
magscale 1 2
timestamp 1674174879
<< viali >>
rect 37473 37281 37507 37315
rect 1593 37213 1627 37247
rect 2513 37213 2547 37247
rect 3157 37213 3191 37247
rect 4169 37213 4203 37247
rect 4813 37213 4847 37247
rect 6561 37213 6595 37247
rect 7849 37213 7883 37247
rect 9321 37213 9355 37247
rect 10425 37213 10459 37247
rect 12357 37213 12391 37247
rect 14473 37213 14507 37247
rect 15577 37213 15611 37247
rect 16865 37213 16899 37247
rect 18337 37213 18371 37247
rect 20085 37213 20119 37247
rect 22017 37213 22051 37247
rect 22937 37213 22971 37247
rect 24777 37213 24811 37247
rect 26065 37213 26099 37247
rect 27813 37213 27847 37247
rect 29745 37213 29779 37247
rect 30665 37213 30699 37247
rect 32505 37213 32539 37247
rect 33793 37213 33827 37247
rect 34897 37213 34931 37247
rect 36645 37213 36679 37247
rect 37749 37213 37783 37247
rect 1777 37077 1811 37111
rect 2329 37077 2363 37111
rect 2973 37077 3007 37111
rect 3985 37077 4019 37111
rect 4629 37077 4663 37111
rect 6745 37077 6779 37111
rect 8033 37077 8067 37111
rect 9137 37077 9171 37111
rect 10609 37077 10643 37111
rect 12541 37077 12575 37111
rect 14289 37077 14323 37111
rect 15761 37077 15795 37111
rect 17049 37077 17083 37111
rect 18153 37077 18187 37111
rect 20269 37077 20303 37111
rect 22201 37077 22235 37111
rect 22753 37077 22787 37111
rect 24593 37077 24627 37111
rect 25881 37077 25915 37111
rect 27997 37077 28031 37111
rect 29929 37077 29963 37111
rect 30481 37077 30515 37111
rect 32321 37077 32355 37111
rect 33609 37077 33643 37111
rect 35081 37077 35115 37111
rect 36829 37077 36863 37111
rect 1777 36873 1811 36907
rect 38209 36873 38243 36907
rect 1593 36737 1627 36771
rect 36921 36737 36955 36771
rect 38025 36737 38059 36771
rect 36737 36533 36771 36567
rect 38301 36125 38335 36159
rect 38117 35989 38151 36023
rect 7021 35241 7055 35275
rect 7205 35037 7239 35071
rect 38025 35037 38059 35071
rect 38209 34901 38243 34935
rect 31493 34697 31527 34731
rect 32413 34697 32447 34731
rect 31677 34561 31711 34595
rect 32597 34561 32631 34595
rect 1777 33473 1811 33507
rect 38301 33473 38335 33507
rect 1593 33269 1627 33303
rect 38117 33269 38151 33303
rect 11897 33065 11931 33099
rect 31217 33065 31251 33099
rect 32781 33065 32815 33099
rect 12081 32861 12115 32895
rect 31125 32861 31159 32895
rect 32965 32861 32999 32895
rect 4169 32521 4203 32555
rect 11713 32521 11747 32555
rect 17509 32521 17543 32555
rect 28641 32521 28675 32555
rect 1777 32385 1811 32419
rect 4353 32385 4387 32419
rect 11897 32385 11931 32419
rect 17693 32385 17727 32419
rect 28825 32385 28859 32419
rect 38025 32385 38059 32419
rect 1593 32181 1627 32215
rect 38209 32181 38243 32215
rect 9965 31977 9999 32011
rect 16865 31977 16899 32011
rect 30021 31841 30055 31875
rect 10149 31773 10183 31807
rect 17049 31773 17083 31807
rect 26985 31773 27019 31807
rect 29929 31773 29963 31807
rect 26801 31637 26835 31671
rect 25973 31433 26007 31467
rect 15301 31297 15335 31331
rect 15945 31297 15979 31331
rect 19717 31297 19751 31331
rect 26157 31297 26191 31331
rect 30665 31297 30699 31331
rect 20177 31229 20211 31263
rect 15117 31161 15151 31195
rect 15761 31093 15795 31127
rect 19533 31093 19567 31127
rect 30481 31093 30515 31127
rect 14289 30889 14323 30923
rect 17417 30889 17451 30923
rect 18061 30889 18095 30923
rect 19533 30753 19567 30787
rect 19717 30753 19751 30787
rect 23305 30753 23339 30787
rect 1593 30685 1627 30719
rect 1869 30685 1903 30719
rect 11253 30685 11287 30719
rect 11897 30685 11931 30719
rect 14473 30685 14507 30719
rect 17325 30685 17359 30719
rect 18245 30685 18279 30719
rect 22569 30685 22603 30719
rect 33333 30685 33367 30719
rect 23397 30617 23431 30651
rect 23949 30617 23983 30651
rect 11069 30549 11103 30583
rect 11713 30549 11747 30583
rect 20177 30549 20211 30583
rect 22661 30549 22695 30583
rect 33425 30549 33459 30583
rect 14933 30345 14967 30379
rect 19533 30345 19567 30379
rect 10609 30277 10643 30311
rect 12541 30277 12575 30311
rect 14289 30277 14323 30311
rect 16957 30277 16991 30311
rect 28917 30277 28951 30311
rect 10517 30209 10551 30243
rect 12449 30209 12483 30243
rect 14197 30209 14231 30243
rect 14841 30209 14875 30243
rect 16865 30209 16899 30243
rect 19717 30209 19751 30243
rect 23121 30209 23155 30243
rect 28825 30209 28859 30243
rect 33609 30209 33643 30243
rect 38025 30209 38059 30243
rect 7113 30141 7147 30175
rect 7297 30141 7331 30175
rect 33425 30073 33459 30107
rect 7757 30005 7791 30039
rect 23213 30005 23247 30039
rect 38209 30005 38243 30039
rect 5181 29801 5215 29835
rect 7297 29801 7331 29835
rect 11253 29801 11287 29835
rect 15025 29801 15059 29835
rect 24869 29801 24903 29835
rect 28181 29801 28215 29835
rect 10609 29733 10643 29767
rect 12449 29733 12483 29767
rect 20085 29733 20119 29767
rect 14841 29665 14875 29699
rect 19717 29665 19751 29699
rect 5089 29597 5123 29631
rect 7205 29597 7239 29631
rect 11161 29597 11195 29631
rect 14657 29597 14691 29631
rect 15761 29597 15795 29631
rect 19901 29597 19935 29631
rect 21097 29597 21131 29631
rect 24777 29597 24811 29631
rect 28089 29597 28123 29631
rect 10057 29529 10091 29563
rect 10149 29529 10183 29563
rect 11897 29529 11931 29563
rect 11989 29529 12023 29563
rect 18153 29529 18187 29563
rect 18245 29529 18279 29563
rect 18797 29529 18831 29563
rect 15853 29461 15887 29495
rect 21281 29461 21315 29495
rect 8677 29257 8711 29291
rect 10057 29257 10091 29291
rect 11897 29257 11931 29291
rect 15117 29257 15151 29291
rect 18153 29257 18187 29291
rect 19349 29257 19383 29291
rect 19993 29257 20027 29291
rect 20821 29257 20855 29291
rect 1777 29121 1811 29155
rect 9965 29121 9999 29155
rect 14473 29121 14507 29155
rect 14657 29121 14691 29155
rect 19257 29121 19291 29155
rect 19901 29121 19935 29155
rect 21005 29121 21039 29155
rect 38301 29121 38335 29155
rect 8033 29053 8067 29087
rect 8217 29053 8251 29087
rect 1593 28985 1627 29019
rect 38117 28985 38151 29019
rect 13093 28713 13127 28747
rect 29009 28713 29043 28747
rect 7757 28645 7791 28679
rect 7665 28509 7699 28543
rect 8493 28509 8527 28543
rect 10241 28509 10275 28543
rect 10701 28509 10735 28543
rect 12725 28509 12759 28543
rect 12909 28509 12943 28543
rect 15393 28509 15427 28543
rect 16037 28509 16071 28543
rect 28917 28509 28951 28543
rect 31033 28509 31067 28543
rect 8309 28373 8343 28407
rect 10057 28373 10091 28407
rect 10793 28373 10827 28407
rect 14565 28373 14599 28407
rect 15209 28373 15243 28407
rect 15853 28373 15887 28407
rect 19901 28373 19935 28407
rect 31125 28373 31159 28407
rect 8217 28169 8251 28203
rect 12081 28169 12115 28203
rect 13277 28169 13311 28203
rect 23489 28169 23523 28203
rect 28549 28169 28583 28203
rect 35449 28169 35483 28203
rect 14473 28101 14507 28135
rect 14565 28101 14599 28135
rect 19625 28101 19659 28135
rect 19717 28101 19751 28135
rect 20913 28101 20947 28135
rect 6929 28033 6963 28067
rect 8401 28033 8435 28067
rect 8953 28033 8987 28067
rect 10057 28033 10091 28067
rect 11989 28033 12023 28067
rect 22017 28033 22051 28067
rect 23673 28033 23707 28067
rect 24317 28033 24351 28067
rect 27353 28033 27387 28067
rect 27997 28033 28031 28067
rect 28457 28033 28491 28067
rect 29469 28033 29503 28067
rect 35633 28033 35667 28067
rect 9045 27965 9079 27999
rect 9873 27965 9907 27999
rect 12633 27965 12667 27999
rect 12817 27965 12851 27999
rect 20821 27965 20855 27999
rect 24869 27965 24903 27999
rect 25053 27965 25087 27999
rect 29653 27965 29687 27999
rect 15025 27897 15059 27931
rect 20177 27897 20211 27931
rect 21373 27897 21407 27931
rect 22109 27897 22143 27931
rect 24133 27897 24167 27931
rect 25513 27897 25547 27931
rect 27813 27897 27847 27931
rect 7021 27829 7055 27863
rect 10517 27829 10551 27863
rect 27169 27829 27203 27863
rect 29837 27829 29871 27863
rect 29837 27625 29871 27659
rect 6561 27557 6595 27591
rect 11621 27557 11655 27591
rect 32965 27557 32999 27591
rect 10149 27489 10183 27523
rect 12725 27489 12759 27523
rect 26433 27489 26467 27523
rect 1777 27421 1811 27455
rect 5733 27421 5767 27455
rect 6745 27421 6779 27455
rect 7205 27421 7239 27455
rect 8033 27421 8067 27455
rect 9321 27421 9355 27455
rect 10333 27421 10367 27455
rect 10793 27421 10827 27455
rect 11253 27421 11287 27455
rect 11437 27421 11471 27455
rect 16773 27421 16807 27455
rect 26617 27421 26651 27455
rect 28825 27421 28859 27455
rect 29745 27421 29779 27455
rect 32873 27421 32907 27455
rect 38025 27421 38059 27455
rect 7297 27353 7331 27387
rect 17509 27353 17543 27387
rect 17601 27353 17635 27387
rect 18153 27353 18187 27387
rect 1593 27285 1627 27319
rect 5825 27285 5859 27319
rect 7849 27285 7883 27319
rect 9137 27285 9171 27319
rect 16865 27285 16899 27319
rect 27077 27285 27111 27319
rect 28917 27285 28951 27319
rect 38209 27285 38243 27319
rect 10241 27081 10275 27115
rect 11805 27081 11839 27115
rect 18153 27081 18187 27115
rect 19165 27081 19199 27115
rect 22017 27081 22051 27115
rect 23305 27081 23339 27115
rect 25881 27081 25915 27115
rect 13277 27013 13311 27047
rect 13369 27013 13403 27047
rect 7113 26945 7147 26979
rect 9137 26945 9171 26979
rect 10149 26945 10183 26979
rect 10977 26945 11011 26979
rect 11713 26945 11747 26979
rect 14749 26945 14783 26979
rect 17417 26945 17451 26979
rect 17969 26945 18003 26979
rect 19349 26945 19383 26979
rect 21189 26945 21223 26979
rect 22201 26945 22235 26979
rect 22845 26945 22879 26979
rect 23489 26945 23523 26979
rect 24133 26945 24167 26979
rect 25145 26945 25179 26979
rect 25789 26945 25823 26979
rect 32413 26945 32447 26979
rect 7297 26877 7331 26911
rect 14933 26877 14967 26911
rect 16129 26877 16163 26911
rect 26433 26877 26467 26911
rect 10793 26809 10827 26843
rect 13829 26809 13863 26843
rect 22661 26809 22695 26843
rect 7757 26741 7791 26775
rect 8953 26741 8987 26775
rect 15393 26741 15427 26775
rect 17233 26741 17267 26775
rect 21005 26741 21039 26775
rect 23949 26741 23983 26775
rect 25237 26741 25271 26775
rect 32505 26741 32539 26775
rect 9781 26537 9815 26571
rect 12081 26537 12115 26571
rect 13553 26537 13587 26571
rect 14565 26537 14599 26571
rect 17601 26537 17635 26571
rect 20177 26537 20211 26571
rect 27813 26537 27847 26571
rect 12725 26469 12759 26503
rect 24961 26469 24995 26503
rect 9137 26401 9171 26435
rect 9321 26401 9355 26435
rect 16497 26401 16531 26435
rect 16681 26401 16715 26435
rect 17141 26401 17175 26435
rect 20913 26401 20947 26435
rect 21557 26401 21591 26435
rect 25973 26401 26007 26435
rect 26157 26401 26191 26435
rect 12265 26333 12299 26367
rect 12909 26333 12943 26367
rect 13737 26333 13771 26367
rect 14473 26333 14507 26367
rect 17785 26333 17819 26367
rect 20361 26333 20395 26367
rect 25145 26333 25179 26367
rect 26617 26333 26651 26367
rect 27445 26333 27479 26367
rect 27629 26333 27663 26367
rect 28825 26333 28859 26367
rect 21005 26265 21039 26299
rect 28917 26265 28951 26299
rect 7297 26197 7331 26231
rect 23121 26197 23155 26231
rect 7941 25993 7975 26027
rect 14381 25993 14415 26027
rect 18889 25993 18923 26027
rect 20177 25993 20211 26027
rect 20821 25993 20855 26027
rect 26157 25993 26191 26027
rect 27813 25993 27847 26027
rect 8953 25925 8987 25959
rect 9045 25925 9079 25959
rect 15577 25925 15611 25959
rect 23029 25925 23063 25959
rect 23121 25925 23155 25959
rect 24317 25925 24351 25959
rect 7297 25857 7331 25891
rect 7481 25857 7515 25891
rect 11161 25857 11195 25891
rect 11713 25857 11747 25891
rect 13645 25857 13679 25891
rect 14565 25857 14599 25891
rect 16129 25857 16163 25891
rect 19073 25857 19107 25891
rect 20361 25857 20395 25891
rect 21005 25857 21039 25891
rect 23673 25857 23707 25891
rect 26341 25857 26375 25891
rect 27169 25857 27203 25891
rect 9597 25789 9631 25823
rect 11897 25789 11931 25823
rect 12817 25789 12851 25823
rect 15485 25789 15519 25823
rect 24225 25789 24259 25823
rect 24501 25789 24535 25823
rect 27353 25789 27387 25823
rect 12357 25721 12391 25755
rect 10977 25653 11011 25687
rect 13461 25653 13495 25687
rect 8309 25449 8343 25483
rect 9781 25449 9815 25483
rect 11529 25449 11563 25483
rect 13369 25449 13403 25483
rect 15485 25449 15519 25483
rect 16129 25449 16163 25483
rect 16773 25381 16807 25415
rect 20085 25381 20119 25415
rect 28457 25381 28491 25415
rect 32137 25381 32171 25415
rect 12725 25313 12759 25347
rect 12909 25313 12943 25347
rect 25053 25313 25087 25347
rect 31769 25313 31803 25347
rect 1777 25245 1811 25279
rect 8217 25245 8251 25279
rect 9965 25245 9999 25279
rect 11713 25245 11747 25279
rect 15669 25245 15703 25279
rect 16313 25245 16347 25279
rect 16957 25245 16991 25279
rect 18705 25245 18739 25279
rect 28365 25245 28399 25279
rect 31953 25245 31987 25279
rect 38301 25245 38335 25279
rect 19533 25177 19567 25211
rect 19625 25177 19659 25211
rect 25145 25177 25179 25211
rect 25697 25177 25731 25211
rect 1593 25109 1627 25143
rect 18797 25109 18831 25143
rect 38117 25109 38151 25143
rect 10885 24905 10919 24939
rect 12357 24905 12391 24939
rect 27261 24905 27295 24939
rect 14933 24837 14967 24871
rect 22201 24837 22235 24871
rect 5365 24769 5399 24803
rect 7573 24769 7607 24803
rect 11069 24769 11103 24803
rect 12541 24769 12575 24803
rect 13001 24769 13035 24803
rect 27169 24769 27203 24803
rect 13185 24701 13219 24735
rect 14841 24701 14875 24735
rect 15485 24701 15519 24735
rect 22109 24701 22143 24735
rect 22661 24633 22695 24667
rect 5457 24565 5491 24599
rect 7665 24565 7699 24599
rect 13369 24565 13403 24599
rect 4261 24361 4295 24395
rect 15945 24361 15979 24395
rect 20821 24361 20855 24395
rect 24777 24361 24811 24395
rect 32045 24361 32079 24395
rect 13461 24293 13495 24327
rect 18245 24225 18279 24259
rect 18889 24225 18923 24259
rect 19625 24225 19659 24259
rect 19993 24225 20027 24259
rect 25421 24225 25455 24259
rect 26065 24225 26099 24259
rect 1593 24157 1627 24191
rect 4169 24157 4203 24191
rect 7573 24157 7607 24191
rect 7757 24157 7791 24191
rect 11161 24157 11195 24191
rect 13001 24157 13035 24191
rect 13645 24157 13679 24191
rect 16129 24157 16163 24191
rect 20729 24157 20763 24191
rect 22201 24157 22235 24191
rect 24685 24157 24719 24191
rect 28457 24157 28491 24191
rect 31309 24157 31343 24191
rect 31953 24157 31987 24191
rect 38301 24157 38335 24191
rect 11253 24089 11287 24123
rect 18337 24089 18371 24123
rect 19717 24089 19751 24123
rect 25513 24089 25547 24123
rect 1777 24021 1811 24055
rect 8217 24021 8251 24055
rect 10517 24021 10551 24055
rect 12817 24021 12851 24055
rect 22017 24021 22051 24055
rect 28457 24021 28491 24055
rect 31401 24021 31435 24055
rect 38117 24021 38151 24055
rect 7113 23817 7147 23851
rect 11161 23817 11195 23851
rect 12817 23817 12851 23851
rect 13369 23817 13403 23851
rect 21373 23817 21407 23851
rect 31769 23817 31803 23851
rect 33333 23817 33367 23851
rect 17049 23749 17083 23783
rect 22661 23749 22695 23783
rect 7297 23681 7331 23715
rect 10517 23681 10551 23715
rect 10701 23681 10735 23715
rect 12357 23681 12391 23715
rect 13277 23681 13311 23715
rect 15025 23681 15059 23715
rect 21281 23681 21315 23715
rect 29193 23681 29227 23715
rect 32505 23681 32539 23715
rect 33517 23681 33551 23715
rect 12173 23613 12207 23647
rect 16957 23613 16991 23647
rect 22569 23613 22603 23647
rect 22845 23613 22879 23647
rect 30481 23613 30515 23647
rect 31125 23613 31159 23647
rect 31309 23613 31343 23647
rect 17509 23545 17543 23579
rect 32321 23545 32355 23579
rect 14841 23477 14875 23511
rect 29285 23477 29319 23511
rect 7941 23273 7975 23307
rect 16221 23273 16255 23307
rect 17141 23273 17175 23307
rect 18061 23273 18095 23307
rect 20361 23273 20395 23307
rect 31217 23273 31251 23307
rect 25421 23205 25455 23239
rect 28917 23205 28951 23239
rect 30113 23205 30147 23239
rect 12173 23137 12207 23171
rect 14381 23137 14415 23171
rect 15393 23137 15427 23171
rect 26985 23137 27019 23171
rect 28273 23137 28307 23171
rect 29929 23137 29963 23171
rect 7849 23069 7883 23103
rect 15853 23069 15887 23103
rect 16037 23069 16071 23103
rect 17325 23069 17359 23103
rect 17969 23069 18003 23103
rect 19901 23069 19935 23103
rect 20545 23069 20579 23103
rect 21833 23069 21867 23103
rect 25605 23069 25639 23103
rect 26249 23069 26283 23103
rect 27169 23069 27203 23103
rect 28457 23069 28491 23103
rect 29745 23069 29779 23103
rect 31401 23069 31435 23103
rect 34897 23069 34931 23103
rect 14473 23001 14507 23035
rect 19717 22933 19751 22967
rect 21649 22933 21683 22967
rect 26065 22933 26099 22967
rect 27629 22933 27663 22967
rect 34989 22933 35023 22967
rect 15117 22729 15151 22763
rect 16221 22729 16255 22763
rect 19809 22729 19843 22763
rect 21281 22729 21315 22763
rect 27813 22729 27847 22763
rect 5365 22661 5399 22695
rect 5457 22661 5491 22695
rect 8861 22661 8895 22695
rect 9413 22661 9447 22695
rect 11897 22661 11931 22695
rect 22385 22661 22419 22695
rect 23673 22661 23707 22695
rect 24225 22661 24259 22695
rect 25881 22661 25915 22695
rect 26433 22661 26467 22695
rect 1777 22593 1811 22627
rect 3157 22593 3191 22627
rect 13461 22593 13495 22627
rect 15301 22593 15335 22627
rect 16129 22593 16163 22627
rect 17141 22593 17175 22627
rect 18245 22593 18279 22627
rect 18889 22593 18923 22627
rect 19993 22593 20027 22627
rect 21465 22593 21499 22627
rect 27353 22593 27387 22627
rect 27997 22593 28031 22627
rect 28457 22593 28491 22627
rect 30481 22593 30515 22627
rect 8769 22525 8803 22559
rect 10241 22525 10275 22559
rect 11805 22525 11839 22559
rect 12081 22525 12115 22559
rect 22293 22525 22327 22559
rect 22569 22525 22603 22559
rect 23581 22525 23615 22559
rect 25789 22525 25823 22559
rect 28641 22525 28675 22559
rect 30665 22525 30699 22559
rect 1593 22457 1627 22491
rect 5917 22457 5951 22491
rect 16957 22457 16991 22491
rect 18705 22457 18739 22491
rect 27169 22457 27203 22491
rect 3249 22389 3283 22423
rect 13277 22389 13311 22423
rect 18061 22389 18095 22423
rect 29009 22389 29043 22423
rect 30849 22389 30883 22423
rect 9229 22185 9263 22219
rect 16221 22185 16255 22219
rect 26617 22185 26651 22219
rect 28825 22185 28859 22219
rect 30389 22185 30423 22219
rect 30849 22185 30883 22219
rect 6377 22049 6411 22083
rect 7021 22049 7055 22083
rect 10149 22049 10183 22083
rect 11529 22049 11563 22083
rect 17417 22049 17451 22083
rect 22293 22049 22327 22083
rect 23213 22049 23247 22083
rect 24685 22049 24719 22083
rect 25881 22049 25915 22083
rect 29745 22049 29779 22083
rect 6285 21981 6319 22015
rect 8493 21981 8527 22015
rect 9137 21981 9171 22015
rect 10333 21981 10367 22015
rect 13277 21981 13311 22015
rect 16129 21981 16163 22015
rect 16773 21981 16807 22015
rect 16957 21981 16991 22015
rect 20453 21981 20487 22015
rect 20913 21981 20947 22015
rect 23121 21981 23155 22015
rect 24593 21981 24627 22015
rect 26525 21981 26559 22015
rect 28733 21981 28767 22015
rect 29929 21981 29963 22015
rect 31033 21981 31067 22015
rect 37473 21981 37507 22015
rect 37749 21981 37783 22015
rect 7113 21913 7147 21947
rect 7665 21913 7699 21947
rect 22017 21913 22051 21947
rect 22109 21913 22143 21947
rect 8309 21845 8343 21879
rect 10793 21845 10827 21879
rect 13093 21845 13127 21879
rect 20269 21845 20303 21879
rect 21005 21845 21039 21879
rect 28089 21845 28123 21879
rect 7113 21641 7147 21675
rect 8677 21641 8711 21675
rect 10885 21641 10919 21675
rect 12081 21641 12115 21675
rect 13921 21641 13955 21675
rect 28733 21641 28767 21675
rect 29285 21641 29319 21675
rect 29837 21641 29871 21675
rect 9873 21573 9907 21607
rect 17969 21573 18003 21607
rect 19901 21573 19935 21607
rect 20453 21573 20487 21607
rect 22201 21573 22235 21607
rect 7297 21505 7331 21539
rect 8861 21505 8895 21539
rect 11069 21505 11103 21539
rect 12265 21505 12299 21539
rect 28089 21505 28123 21539
rect 29193 21505 29227 21539
rect 30021 21505 30055 21539
rect 7941 21437 7975 21471
rect 9781 21437 9815 21471
rect 13277 21437 13311 21471
rect 13461 21437 13495 21471
rect 17877 21437 17911 21471
rect 18153 21437 18187 21471
rect 19809 21437 19843 21471
rect 22109 21437 22143 21471
rect 22385 21437 22419 21471
rect 28273 21437 28307 21471
rect 10333 21369 10367 21403
rect 4997 21097 5031 21131
rect 7021 21097 7055 21131
rect 9229 21097 9263 21131
rect 9873 21097 9907 21131
rect 13093 21097 13127 21131
rect 28273 21097 28307 21131
rect 15669 21029 15703 21063
rect 17969 21029 18003 21063
rect 27629 21029 27663 21063
rect 7941 20961 7975 20995
rect 15117 20961 15151 20995
rect 1777 20893 1811 20927
rect 4905 20893 4939 20927
rect 7205 20893 7239 20927
rect 8585 20893 8619 20927
rect 9137 20893 9171 20927
rect 10057 20893 10091 20927
rect 13001 20893 13035 20927
rect 14565 20893 14599 20927
rect 19441 20893 19475 20927
rect 20821 20893 20855 20927
rect 25605 20893 25639 20927
rect 27813 20893 27847 20927
rect 28457 20893 28491 20927
rect 29745 20893 29779 20927
rect 30389 20893 30423 20927
rect 38301 20893 38335 20927
rect 8033 20825 8067 20859
rect 15209 20825 15243 20859
rect 17417 20825 17451 20859
rect 17509 20825 17543 20859
rect 1593 20757 1627 20791
rect 14381 20757 14415 20791
rect 19533 20757 19567 20791
rect 20637 20757 20671 20791
rect 25421 20757 25455 20791
rect 29837 20757 29871 20791
rect 30481 20757 30515 20791
rect 38117 20757 38151 20791
rect 5917 20553 5951 20587
rect 10977 20553 11011 20587
rect 24961 20553 24995 20587
rect 8125 20485 8159 20519
rect 8217 20485 8251 20519
rect 23581 20485 23615 20519
rect 29377 20485 29411 20519
rect 2789 20417 2823 20451
rect 5825 20417 5859 20451
rect 6561 20417 6595 20451
rect 11161 20417 11195 20451
rect 12725 20417 12759 20451
rect 14657 20417 14691 20451
rect 15669 20417 15703 20451
rect 25145 20417 25179 20451
rect 25881 20417 25915 20451
rect 26525 20417 26559 20451
rect 27353 20417 27387 20451
rect 28273 20417 28307 20451
rect 2973 20349 3007 20383
rect 11897 20349 11931 20383
rect 12541 20349 12575 20383
rect 15853 20349 15887 20383
rect 20821 20349 20855 20383
rect 21005 20349 21039 20383
rect 23489 20349 23523 20383
rect 28089 20349 28123 20383
rect 29285 20349 29319 20383
rect 8677 20281 8711 20315
rect 13185 20281 13219 20315
rect 16037 20281 16071 20315
rect 24041 20281 24075 20315
rect 25697 20281 25731 20315
rect 29837 20281 29871 20315
rect 3433 20213 3467 20247
rect 6653 20213 6687 20247
rect 14473 20213 14507 20247
rect 21189 20213 21223 20247
rect 26341 20213 26375 20247
rect 27169 20213 27203 20247
rect 28733 20213 28767 20247
rect 9781 20009 9815 20043
rect 12081 20009 12115 20043
rect 12817 20009 12851 20043
rect 15761 20009 15795 20043
rect 21373 20009 21407 20043
rect 28549 20009 28583 20043
rect 30757 20009 30791 20043
rect 14933 19941 14967 19975
rect 27445 19941 27479 19975
rect 5089 19873 5123 19907
rect 5733 19873 5767 19907
rect 11161 19873 11195 19907
rect 17141 19873 17175 19907
rect 22845 19873 22879 19907
rect 26341 19873 26375 19907
rect 26893 19873 26927 19907
rect 6193 19805 6227 19839
rect 9965 19805 9999 19839
rect 12265 19805 12299 19839
rect 12725 19805 12759 19839
rect 14289 19805 14323 19839
rect 15117 19805 15151 19839
rect 15669 19805 15703 19839
rect 16497 19805 16531 19839
rect 21281 19805 21315 19839
rect 28457 19805 28491 19839
rect 30205 19805 30239 19839
rect 30665 19805 30699 19839
rect 31493 19805 31527 19839
rect 5181 19737 5215 19771
rect 10517 19737 10551 19771
rect 10609 19737 10643 19771
rect 14381 19737 14415 19771
rect 17233 19737 17267 19771
rect 17785 19737 17819 19771
rect 22569 19737 22603 19771
rect 22661 19737 22695 19771
rect 25697 19737 25731 19771
rect 25789 19737 25823 19771
rect 26985 19737 27019 19771
rect 6285 19669 6319 19703
rect 16313 19669 16347 19703
rect 30021 19669 30055 19703
rect 31309 19669 31343 19703
rect 4905 19465 4939 19499
rect 9781 19465 9815 19499
rect 10977 19465 11011 19499
rect 11805 19465 11839 19499
rect 17141 19465 17175 19499
rect 19257 19465 19291 19499
rect 20821 19465 20855 19499
rect 22109 19465 22143 19499
rect 27169 19465 27203 19499
rect 14197 19397 14231 19431
rect 17969 19397 18003 19431
rect 18521 19397 18555 19431
rect 1593 19329 1627 19363
rect 4261 19329 4295 19363
rect 5549 19329 5583 19363
rect 9689 19329 9723 19363
rect 11161 19329 11195 19363
rect 11989 19329 12023 19363
rect 15209 19329 15243 19363
rect 15853 19329 15887 19363
rect 17325 19329 17359 19363
rect 19441 19329 19475 19363
rect 22017 19329 22051 19363
rect 27353 19329 27387 19363
rect 30481 19329 30515 19363
rect 4445 19261 4479 19295
rect 14105 19261 14139 19295
rect 15393 19261 15427 19295
rect 17877 19261 17911 19295
rect 20177 19261 20211 19295
rect 20361 19261 20395 19295
rect 29837 19261 29871 19295
rect 30021 19261 30055 19295
rect 5365 19193 5399 19227
rect 14657 19193 14691 19227
rect 1777 19125 1811 19159
rect 4537 18921 4571 18955
rect 5181 18921 5215 18955
rect 14289 18921 14323 18955
rect 16129 18921 16163 18955
rect 22385 18921 22419 18955
rect 5825 18785 5859 18819
rect 6101 18785 6135 18819
rect 17233 18785 17267 18819
rect 18245 18785 18279 18819
rect 24593 18785 24627 18819
rect 29929 18785 29963 18819
rect 4445 18717 4479 18751
rect 5089 18717 5123 18751
rect 6929 18717 6963 18751
rect 7113 18717 7147 18751
rect 8033 18717 8067 18751
rect 11069 18717 11103 18751
rect 14473 18717 14507 18751
rect 16037 18717 16071 18751
rect 20637 18717 20671 18751
rect 21557 18717 21591 18751
rect 22293 18717 22327 18751
rect 24777 18717 24811 18751
rect 28273 18717 28307 18751
rect 5917 18649 5951 18683
rect 8125 18649 8159 18683
rect 11990 18649 12024 18683
rect 12081 18649 12115 18683
rect 12633 18649 12667 18683
rect 17325 18649 17359 18683
rect 7573 18581 7607 18615
rect 9229 18581 9263 18615
rect 11161 18581 11195 18615
rect 20729 18581 20763 18615
rect 21373 18581 21407 18615
rect 25237 18581 25271 18615
rect 28089 18581 28123 18615
rect 1593 18377 1627 18411
rect 5549 18377 5583 18411
rect 12173 18377 12207 18411
rect 17233 18377 17267 18411
rect 23949 18377 23983 18411
rect 28457 18377 28491 18411
rect 8493 18309 8527 18343
rect 9413 18309 9447 18343
rect 12817 18309 12851 18343
rect 12909 18309 12943 18343
rect 14197 18309 14231 18343
rect 17969 18309 18003 18343
rect 18705 18309 18739 18343
rect 21189 18309 21223 18343
rect 24593 18309 24627 18343
rect 24685 18309 24719 18343
rect 25789 18309 25823 18343
rect 1777 18241 1811 18275
rect 5365 18241 5399 18275
rect 7297 18241 7331 18275
rect 10057 18241 10091 18275
rect 12081 18241 12115 18275
rect 17417 18241 17451 18275
rect 17877 18241 17911 18275
rect 20545 18241 20579 18275
rect 20729 18241 20763 18275
rect 22017 18241 22051 18275
rect 23857 18241 23891 18275
rect 25697 18241 25731 18275
rect 27353 18241 27387 18275
rect 28641 18241 28675 18275
rect 31217 18241 31251 18275
rect 8401 18173 8435 18207
rect 13093 18173 13127 18207
rect 14105 18173 14139 18207
rect 14749 18173 14783 18207
rect 18613 18173 18647 18207
rect 18889 18173 18923 18207
rect 22201 18173 22235 18207
rect 25237 18173 25271 18207
rect 27537 18173 27571 18207
rect 29101 18173 29135 18207
rect 7113 18105 7147 18139
rect 9873 18037 9907 18071
rect 22385 18037 22419 18071
rect 27997 18037 28031 18071
rect 31033 18037 31067 18071
rect 5457 17833 5491 17867
rect 8401 17833 8435 17867
rect 11069 17833 11103 17867
rect 13645 17833 13679 17867
rect 14381 17833 14415 17867
rect 17049 17833 17083 17867
rect 21833 17833 21867 17867
rect 22569 17833 22603 17867
rect 26893 17833 26927 17867
rect 2145 17765 2179 17799
rect 6929 17765 6963 17799
rect 7665 17765 7699 17799
rect 28365 17765 28399 17799
rect 4169 17697 4203 17731
rect 9229 17697 9263 17731
rect 10701 17697 10735 17731
rect 11897 17697 11931 17731
rect 16405 17697 16439 17731
rect 16589 17697 16623 17731
rect 18705 17697 18739 17731
rect 20085 17697 20119 17731
rect 28181 17697 28215 17731
rect 2329 17629 2363 17663
rect 3249 17629 3283 17663
rect 3985 17629 4019 17663
rect 5641 17629 5675 17663
rect 6285 17629 6319 17663
rect 7113 17629 7147 17663
rect 7849 17629 7883 17663
rect 8585 17629 8619 17663
rect 10885 17629 10919 17663
rect 13553 17629 13587 17663
rect 14289 17629 14323 17663
rect 22017 17629 22051 17663
rect 22477 17629 22511 17663
rect 26801 17629 26835 17663
rect 27997 17629 28031 17663
rect 31033 17629 31067 17663
rect 9321 17561 9355 17595
rect 9873 17561 9907 17595
rect 11989 17561 12023 17595
rect 12541 17561 12575 17595
rect 19809 17561 19843 17595
rect 19901 17561 19935 17595
rect 4629 17493 4663 17527
rect 6101 17493 6135 17527
rect 30849 17493 30883 17527
rect 31953 17493 31987 17527
rect 5917 17289 5951 17323
rect 7665 17289 7699 17323
rect 17509 17289 17543 17323
rect 18521 17289 18555 17323
rect 25697 17289 25731 17323
rect 3065 17221 3099 17255
rect 8769 17221 8803 17255
rect 20821 17221 20855 17255
rect 23305 17221 23339 17255
rect 23397 17221 23431 17255
rect 27261 17221 27295 17255
rect 27353 17221 27387 17255
rect 32413 17221 32447 17255
rect 32505 17221 32539 17255
rect 3893 17153 3927 17187
rect 4721 17153 4755 17187
rect 5365 17153 5399 17187
rect 5825 17153 5859 17187
rect 7205 17153 7239 17187
rect 7849 17153 7883 17187
rect 10333 17153 10367 17187
rect 12357 17153 12391 17187
rect 13001 17153 13035 17187
rect 16129 17153 16163 17187
rect 16221 17153 16255 17187
rect 17049 17153 17083 17187
rect 18705 17153 18739 17187
rect 25605 17153 25639 17187
rect 38301 17153 38335 17187
rect 2421 17085 2455 17119
rect 2605 17085 2639 17119
rect 3985 17085 4019 17119
rect 8677 17085 8711 17119
rect 16865 17085 16899 17119
rect 20729 17085 20763 17119
rect 30205 17085 30239 17119
rect 32689 17085 32723 17119
rect 4537 17017 4571 17051
rect 7021 17017 7055 17051
rect 9229 17017 9263 17051
rect 21281 17017 21315 17051
rect 23857 17017 23891 17051
rect 27813 17017 27847 17051
rect 5181 16949 5215 16983
rect 10425 16949 10459 16983
rect 12173 16949 12207 16983
rect 12817 16949 12851 16983
rect 38117 16949 38151 16983
rect 2329 16745 2363 16779
rect 4721 16745 4755 16779
rect 5365 16745 5399 16779
rect 9229 16745 9263 16779
rect 12081 16745 12115 16779
rect 18521 16745 18555 16779
rect 23673 16745 23707 16779
rect 30573 16745 30607 16779
rect 32413 16745 32447 16779
rect 30205 16609 30239 16643
rect 30389 16609 30423 16643
rect 2513 16541 2547 16575
rect 3249 16541 3283 16575
rect 3341 16541 3375 16575
rect 4077 16541 4111 16575
rect 4905 16541 4939 16575
rect 5549 16541 5583 16575
rect 6561 16541 6595 16575
rect 7205 16541 7239 16575
rect 7297 16541 7331 16575
rect 9137 16541 9171 16575
rect 12265 16541 12299 16575
rect 17877 16541 17911 16575
rect 17969 16541 18003 16575
rect 18705 16541 18739 16575
rect 23857 16541 23891 16575
rect 25973 16541 26007 16575
rect 32597 16541 32631 16575
rect 33241 16541 33275 16575
rect 4169 16405 4203 16439
rect 6653 16405 6687 16439
rect 25789 16405 25823 16439
rect 33057 16405 33091 16439
rect 4813 16201 4847 16235
rect 5549 16201 5583 16235
rect 20177 16201 20211 16235
rect 23305 16201 23339 16235
rect 27169 16201 27203 16235
rect 30849 16201 30883 16235
rect 10517 16133 10551 16167
rect 10609 16133 10643 16167
rect 25605 16133 25639 16167
rect 28549 16133 28583 16167
rect 1593 16065 1627 16099
rect 2789 16065 2823 16099
rect 4721 16065 4755 16099
rect 5733 16065 5767 16099
rect 20913 16065 20947 16099
rect 22477 16065 22511 16099
rect 23489 16065 23523 16099
rect 24133 16065 24167 16099
rect 27353 16065 27387 16099
rect 29745 16065 29779 16099
rect 31493 16065 31527 16099
rect 38025 16065 38059 16099
rect 10793 15997 10827 16031
rect 18429 15997 18463 16031
rect 18705 15997 18739 16031
rect 25513 15997 25547 16031
rect 25973 15997 26007 16031
rect 28457 15997 28491 16031
rect 29101 15997 29135 16031
rect 30205 15997 30239 16031
rect 30389 15997 30423 16031
rect 31309 15929 31343 15963
rect 1777 15861 1811 15895
rect 2881 15861 2915 15895
rect 21005 15861 21039 15895
rect 22569 15861 22603 15895
rect 23949 15861 23983 15895
rect 29561 15861 29595 15895
rect 38209 15861 38243 15895
rect 8493 15657 8527 15691
rect 18521 15657 18555 15691
rect 22661 15657 22695 15691
rect 31493 15657 31527 15691
rect 33517 15657 33551 15691
rect 6285 15589 6319 15623
rect 10885 15589 10919 15623
rect 25513 15589 25547 15623
rect 28825 15589 28859 15623
rect 30481 15589 30515 15623
rect 4537 15521 4571 15555
rect 6734 15521 6768 15555
rect 9137 15521 9171 15555
rect 11345 15521 11379 15555
rect 13369 15521 13403 15555
rect 15301 15521 15335 15555
rect 21281 15521 21315 15555
rect 23857 15521 23891 15555
rect 29929 15521 29963 15555
rect 18705 15453 18739 15487
rect 20361 15453 20395 15487
rect 21189 15453 21223 15487
rect 21833 15453 21867 15487
rect 22569 15453 22603 15487
rect 25053 15453 25087 15487
rect 25697 15453 25731 15487
rect 27537 15453 27571 15487
rect 28365 15453 28399 15487
rect 29009 15453 29043 15487
rect 31401 15453 31435 15487
rect 32781 15453 32815 15487
rect 33425 15453 33459 15487
rect 4813 15385 4847 15419
rect 7021 15385 7055 15419
rect 9413 15385 9447 15419
rect 11621 15385 11655 15419
rect 15577 15385 15611 15419
rect 17325 15385 17359 15419
rect 23397 15385 23431 15419
rect 23489 15385 23523 15419
rect 30021 15385 30055 15419
rect 20453 15317 20487 15351
rect 21925 15317 21959 15351
rect 24869 15317 24903 15351
rect 27353 15317 27387 15351
rect 28181 15317 28215 15351
rect 32873 15317 32907 15351
rect 13921 15113 13955 15147
rect 23029 15113 23063 15147
rect 23673 15113 23707 15147
rect 26065 15113 26099 15147
rect 29285 15113 29319 15147
rect 3893 15045 3927 15079
rect 9045 15045 9079 15079
rect 28181 15045 28215 15079
rect 28273 15045 28307 15079
rect 1777 14977 1811 15011
rect 8769 14977 8803 15011
rect 12173 14977 12207 15011
rect 14473 14977 14507 15011
rect 18153 14977 18187 15011
rect 22293 14977 22327 15011
rect 22937 14977 22971 15011
rect 23581 14977 23615 15011
rect 26249 14977 26283 15011
rect 27353 14977 27387 15011
rect 29469 14977 29503 15011
rect 3617 14909 3651 14943
rect 5365 14909 5399 14943
rect 12449 14909 12483 14943
rect 14749 14909 14783 14943
rect 20177 14909 20211 14943
rect 28825 14909 28859 14943
rect 16221 14841 16255 14875
rect 1593 14773 1627 14807
rect 10517 14773 10551 14807
rect 18410 14773 18444 14807
rect 22385 14773 22419 14807
rect 27169 14773 27203 14807
rect 11069 14569 11103 14603
rect 22293 14569 22327 14603
rect 23489 14569 23523 14603
rect 26801 14569 26835 14603
rect 28273 14569 28307 14603
rect 38117 14569 38151 14603
rect 15853 14433 15887 14467
rect 22845 14433 22879 14467
rect 23029 14433 23063 14467
rect 31309 14433 31343 14467
rect 1961 14365 1995 14399
rect 10977 14365 11011 14399
rect 21097 14365 21131 14399
rect 22201 14365 22235 14399
rect 25237 14365 25271 14399
rect 26985 14365 27019 14399
rect 28457 14365 28491 14399
rect 38301 14365 38335 14399
rect 16129 14297 16163 14331
rect 31401 14297 31435 14331
rect 31953 14297 31987 14331
rect 1777 14229 1811 14263
rect 17601 14229 17635 14263
rect 21189 14229 21223 14263
rect 25329 14229 25363 14263
rect 1777 14025 1811 14059
rect 2513 14025 2547 14059
rect 22109 14025 22143 14059
rect 24501 14025 24535 14059
rect 25697 14025 25731 14059
rect 31033 14025 31067 14059
rect 5549 13957 5583 13991
rect 28457 13957 28491 13991
rect 1961 13889 1995 13923
rect 2421 13889 2455 13923
rect 7665 13889 7699 13923
rect 13553 13889 13587 13923
rect 18337 13889 18371 13923
rect 20361 13889 20395 13923
rect 21189 13889 21223 13923
rect 22017 13889 22051 13923
rect 22661 13889 22695 13923
rect 23857 13889 23891 13923
rect 24041 13889 24075 13923
rect 25237 13889 25271 13923
rect 27169 13889 27203 13923
rect 27353 13889 27387 13923
rect 30941 13889 30975 13923
rect 3525 13821 3559 13855
rect 3801 13821 3835 13855
rect 9689 13821 9723 13855
rect 15301 13821 15335 13855
rect 18613 13821 18647 13855
rect 25053 13821 25087 13855
rect 27813 13821 27847 13855
rect 28365 13821 28399 13855
rect 28825 13821 28859 13855
rect 21281 13753 21315 13787
rect 7928 13685 7962 13719
rect 13816 13685 13850 13719
rect 22753 13685 22787 13719
rect 5733 13481 5767 13515
rect 14546 13481 14580 13515
rect 28733 13481 28767 13515
rect 31953 13481 31987 13515
rect 26525 13413 26559 13447
rect 31125 13413 31159 13447
rect 1961 13345 1995 13379
rect 4261 13345 4295 13379
rect 11069 13345 11103 13379
rect 14289 13345 14323 13379
rect 21833 13345 21867 13379
rect 25145 13345 25179 13379
rect 26157 13345 26191 13379
rect 30573 13345 30607 13379
rect 1869 13277 1903 13311
rect 3985 13277 4019 13311
rect 9137 13277 9171 13311
rect 21097 13277 21131 13311
rect 21741 13277 21775 13311
rect 22385 13277 22419 13311
rect 26341 13277 26375 13311
rect 28917 13277 28951 13311
rect 29929 13277 29963 13311
rect 32137 13277 32171 13311
rect 11345 13209 11379 13243
rect 30665 13209 30699 13243
rect 9229 13141 9263 13175
rect 12817 13141 12851 13175
rect 16037 13141 16071 13175
rect 21189 13141 21223 13175
rect 22477 13141 22511 13175
rect 29745 13141 29779 13175
rect 1593 12937 1627 12971
rect 19165 12937 19199 12971
rect 25237 12937 25271 12971
rect 27905 12937 27939 12971
rect 6837 12869 6871 12903
rect 7389 12869 7423 12903
rect 14289 12869 14323 12903
rect 22109 12869 22143 12903
rect 24133 12869 24167 12903
rect 30941 12869 30975 12903
rect 1777 12801 1811 12835
rect 8677 12801 8711 12835
rect 10701 12801 10735 12835
rect 12265 12801 12299 12835
rect 17417 12801 17451 12835
rect 21097 12801 21131 12835
rect 22017 12801 22051 12835
rect 23489 12801 23523 12835
rect 24593 12801 24627 12835
rect 27813 12801 27847 12835
rect 28641 12801 28675 12835
rect 38025 12801 38059 12835
rect 6745 12733 6779 12767
rect 8953 12733 8987 12767
rect 12541 12733 12575 12767
rect 23673 12733 23707 12767
rect 24777 12733 24811 12767
rect 30849 12733 30883 12767
rect 31125 12733 31159 12767
rect 28457 12665 28491 12699
rect 11897 12597 11931 12631
rect 17674 12597 17708 12631
rect 21189 12597 21223 12631
rect 38209 12597 38243 12631
rect 1961 12393 1995 12427
rect 24961 12393 24995 12427
rect 30389 12393 30423 12427
rect 31677 12393 31711 12427
rect 35817 12393 35851 12427
rect 14381 12325 14415 12359
rect 26341 12325 26375 12359
rect 28273 12325 28307 12359
rect 11805 12257 11839 12291
rect 12265 12257 12299 12291
rect 30941 12257 30975 12291
rect 1869 12189 1903 12223
rect 3985 12189 4019 12223
rect 6009 12189 6043 12223
rect 14289 12189 14323 12223
rect 21925 12189 21959 12223
rect 22569 12189 22603 12223
rect 24869 12189 24903 12223
rect 25973 12189 26007 12223
rect 26157 12189 26191 12223
rect 28825 12189 28859 12223
rect 30297 12189 30331 12223
rect 31861 12189 31895 12223
rect 33333 12189 33367 12223
rect 33425 12189 33459 12223
rect 36001 12189 36035 12223
rect 4261 12121 4295 12155
rect 11897 12121 11931 12155
rect 22845 12121 22879 12155
rect 27721 12121 27755 12155
rect 27813 12121 27847 12155
rect 22017 12053 22051 12087
rect 28917 12053 28951 12087
rect 32321 12053 32355 12087
rect 6009 11849 6043 11883
rect 16221 11849 16255 11883
rect 21373 11849 21407 11883
rect 14749 11781 14783 11815
rect 29193 11781 29227 11815
rect 29745 11781 29779 11815
rect 32413 11781 32447 11815
rect 32505 11781 32539 11815
rect 11713 11713 11747 11747
rect 14473 11713 14507 11747
rect 21281 11713 21315 11747
rect 22385 11713 22419 11747
rect 25329 11713 25363 11747
rect 4261 11645 4295 11679
rect 4537 11645 4571 11679
rect 7389 11645 7423 11679
rect 7665 11645 7699 11679
rect 9137 11645 9171 11679
rect 11989 11645 12023 11679
rect 18245 11645 18279 11679
rect 18521 11645 18555 11679
rect 20269 11645 20303 11679
rect 22569 11645 22603 11679
rect 29101 11645 29135 11679
rect 32689 11645 32723 11679
rect 13461 11509 13495 11543
rect 25145 11509 25179 11543
rect 9854 11305 9888 11339
rect 11345 11305 11379 11339
rect 25237 11305 25271 11339
rect 26709 11305 26743 11339
rect 28089 11305 28123 11339
rect 28917 11305 28951 11339
rect 38117 11305 38151 11339
rect 1593 11237 1627 11271
rect 23121 11237 23155 11271
rect 4353 11169 4387 11203
rect 17417 11169 17451 11203
rect 18889 11169 18923 11203
rect 1777 11101 1811 11135
rect 4077 11101 4111 11135
rect 6101 11101 6135 11135
rect 6469 11101 6503 11135
rect 9597 11101 9631 11135
rect 17141 11101 17175 11135
rect 21557 11101 21591 11135
rect 23305 11101 23339 11135
rect 23949 11101 23983 11135
rect 24593 11101 24627 11135
rect 24777 11101 24811 11135
rect 26617 11101 26651 11135
rect 27997 11101 28031 11135
rect 29101 11101 29135 11135
rect 31401 11101 31435 11135
rect 38301 11101 38335 11135
rect 21833 11033 21867 11067
rect 31493 11033 31527 11067
rect 6837 10965 6871 10999
rect 23765 10965 23799 10999
rect 10609 10761 10643 10795
rect 18613 10761 18647 10795
rect 25053 10761 25087 10795
rect 5457 10693 5491 10727
rect 6009 10693 6043 10727
rect 6745 10693 6779 10727
rect 6837 10693 6871 10727
rect 12909 10693 12943 10727
rect 22293 10693 22327 10727
rect 23673 10693 23707 10727
rect 1869 10625 1903 10659
rect 10517 10625 10551 10659
rect 12633 10625 12667 10659
rect 20821 10625 20855 10659
rect 22017 10625 22051 10659
rect 25237 10625 25271 10659
rect 28733 10625 28767 10659
rect 29377 10625 29411 10659
rect 29837 10625 29871 10659
rect 33977 10625 34011 10659
rect 1961 10557 1995 10591
rect 5365 10557 5399 10591
rect 7021 10557 7055 10591
rect 16865 10557 16899 10591
rect 17141 10557 17175 10591
rect 21005 10557 21039 10591
rect 23581 10557 23615 10591
rect 23857 10557 23891 10591
rect 30021 10557 30055 10591
rect 28549 10489 28583 10523
rect 14381 10421 14415 10455
rect 29193 10421 29227 10455
rect 30481 10421 30515 10455
rect 33793 10421 33827 10455
rect 22753 10217 22787 10251
rect 23489 10217 23523 10251
rect 29837 10217 29871 10251
rect 21465 10149 21499 10183
rect 4261 10081 4295 10115
rect 22109 10081 22143 10115
rect 24685 10081 24719 10115
rect 1777 10013 1811 10047
rect 3985 10013 4019 10047
rect 20453 10013 20487 10047
rect 21373 10013 21407 10047
rect 22017 10013 22051 10047
rect 22661 10013 22695 10047
rect 23673 10013 23707 10047
rect 30021 10013 30055 10047
rect 6009 9945 6043 9979
rect 6561 9945 6595 9979
rect 6653 9945 6687 9979
rect 7205 9945 7239 9979
rect 24777 9945 24811 9979
rect 25697 9945 25731 9979
rect 1593 9877 1627 9911
rect 20545 9877 20579 9911
rect 15761 9673 15795 9707
rect 23673 9673 23707 9707
rect 9413 9605 9447 9639
rect 20637 9605 20671 9639
rect 21281 9605 21315 9639
rect 20545 9537 20579 9571
rect 21189 9537 21223 9571
rect 22569 9537 22603 9571
rect 23581 9537 23615 9571
rect 29285 9537 29319 9571
rect 6745 9469 6779 9503
rect 8493 9469 8527 9503
rect 9137 9469 9171 9503
rect 11161 9469 11195 9503
rect 14013 9469 14047 9503
rect 14289 9469 14323 9503
rect 18245 9469 18279 9503
rect 18521 9469 18555 9503
rect 28641 9469 28675 9503
rect 28825 9469 28859 9503
rect 7008 9333 7042 9367
rect 19993 9333 20027 9367
rect 22661 9333 22695 9367
rect 28733 9129 28767 9163
rect 23581 9061 23615 9095
rect 25237 9061 25271 9095
rect 6653 8993 6687 9027
rect 11437 8993 11471 9027
rect 18613 8993 18647 9027
rect 1869 8925 1903 8959
rect 11345 8925 11379 8959
rect 11989 8925 12023 8959
rect 16589 8925 16623 8959
rect 20545 8925 20579 8959
rect 21649 8925 21683 8959
rect 22569 8925 22603 8959
rect 23489 8925 23523 8959
rect 25789 8925 25823 8959
rect 28181 8925 28215 8959
rect 28641 8925 28675 8959
rect 30573 8925 30607 8959
rect 38025 8925 38059 8959
rect 6009 8857 6043 8891
rect 6101 8857 6135 8891
rect 16865 8857 16899 8891
rect 22845 8857 22879 8891
rect 24685 8857 24719 8891
rect 24777 8857 24811 8891
rect 1961 8789 1995 8823
rect 12081 8789 12115 8823
rect 20637 8789 20671 8823
rect 21741 8789 21775 8823
rect 25881 8789 25915 8823
rect 26525 8789 26559 8823
rect 27997 8789 28031 8823
rect 30665 8789 30699 8823
rect 38209 8789 38243 8823
rect 2053 8585 2087 8619
rect 9965 8585 9999 8619
rect 15117 8585 15151 8619
rect 21097 8585 21131 8619
rect 8493 8517 8527 8551
rect 11989 8517 12023 8551
rect 12541 8517 12575 8551
rect 22201 8517 22235 8551
rect 23121 8517 23155 8551
rect 26065 8517 26099 8551
rect 30573 8517 30607 8551
rect 31125 8517 31159 8551
rect 1961 8449 1995 8483
rect 5733 8449 5767 8483
rect 8217 8449 8251 8483
rect 15025 8449 15059 8483
rect 21005 8449 21039 8483
rect 23581 8449 23615 8483
rect 27169 8449 27203 8483
rect 28457 8449 28491 8483
rect 29101 8449 29135 8483
rect 29745 8449 29779 8483
rect 32505 8449 32539 8483
rect 3709 8381 3743 8415
rect 3985 8381 4019 8415
rect 11897 8381 11931 8415
rect 18061 8381 18095 8415
rect 18337 8381 18371 8415
rect 22109 8381 22143 8415
rect 24685 8381 24719 8415
rect 24869 8381 24903 8415
rect 25973 8381 26007 8415
rect 27353 8381 27387 8415
rect 30481 8381 30515 8415
rect 25053 8313 25087 8347
rect 26525 8313 26559 8347
rect 27629 8313 27663 8347
rect 28917 8313 28951 8347
rect 29561 8313 29595 8347
rect 32321 8313 32355 8347
rect 19809 8245 19843 8279
rect 23673 8245 23707 8279
rect 28273 8245 28307 8279
rect 2605 8041 2639 8075
rect 5733 8041 5767 8075
rect 16037 8041 16071 8075
rect 21833 8041 21867 8075
rect 22477 8041 22511 8075
rect 23949 8041 23983 8075
rect 25973 8041 26007 8075
rect 29745 8041 29779 8075
rect 30389 8041 30423 8075
rect 31769 8041 31803 8075
rect 12909 7973 12943 8007
rect 21189 7973 21223 8007
rect 24593 7973 24627 8007
rect 2053 7905 2087 7939
rect 6837 7905 6871 7939
rect 8585 7905 8619 7939
rect 19441 7905 19475 7939
rect 28365 7905 28399 7939
rect 28641 7905 28675 7939
rect 1961 7837 1995 7871
rect 2789 7837 2823 7871
rect 3985 7837 4019 7871
rect 6561 7837 6595 7871
rect 11161 7837 11195 7871
rect 14289 7837 14323 7871
rect 18705 7837 18739 7871
rect 21741 7837 21775 7871
rect 22385 7837 22419 7871
rect 23857 7837 23891 7871
rect 24777 7837 24811 7871
rect 25421 7837 25455 7871
rect 25881 7837 25915 7871
rect 26893 7837 26927 7871
rect 29929 7837 29963 7871
rect 30573 7837 30607 7871
rect 31677 7837 31711 7871
rect 38301 7837 38335 7871
rect 4261 7769 4295 7803
rect 11437 7769 11471 7803
rect 14565 7769 14599 7803
rect 19717 7769 19751 7803
rect 28457 7769 28491 7803
rect 18797 7701 18831 7735
rect 25237 7701 25271 7735
rect 26709 7701 26743 7735
rect 38117 7701 38151 7735
rect 2053 7497 2087 7531
rect 22753 7497 22787 7531
rect 27169 7497 27203 7531
rect 14565 7429 14599 7463
rect 21373 7429 21407 7463
rect 24777 7429 24811 7463
rect 24869 7429 24903 7463
rect 29193 7429 29227 7463
rect 1961 7361 1995 7395
rect 7573 7361 7607 7395
rect 21281 7361 21315 7395
rect 22017 7361 22051 7395
rect 22661 7361 22695 7395
rect 23489 7361 23523 7395
rect 27353 7361 27387 7395
rect 30205 7361 30239 7395
rect 7849 7293 7883 7327
rect 14289 7293 14323 7327
rect 16313 7293 16347 7327
rect 17969 7293 18003 7327
rect 18245 7293 18279 7327
rect 19993 7293 20027 7327
rect 25421 7293 25455 7327
rect 29101 7293 29135 7327
rect 29377 7293 29411 7327
rect 22109 7225 22143 7259
rect 23581 7225 23615 7259
rect 9321 7157 9355 7191
rect 30297 7157 30331 7191
rect 6364 6953 6398 6987
rect 10136 6953 10170 6987
rect 21557 6885 21591 6919
rect 6101 6817 6135 6851
rect 11621 6817 11655 6851
rect 22570 6817 22604 6851
rect 28825 6817 28859 6851
rect 2237 6749 2271 6783
rect 2329 6749 2363 6783
rect 2973 6749 3007 6783
rect 9873 6749 9907 6783
rect 20821 6749 20855 6783
rect 21465 6749 21499 6783
rect 22385 6749 22419 6783
rect 23489 6749 23523 6783
rect 28733 6749 28767 6783
rect 23581 6681 23615 6715
rect 2789 6613 2823 6647
rect 7849 6613 7883 6647
rect 20913 6613 20947 6647
rect 23029 6613 23063 6647
rect 2053 6409 2087 6443
rect 10425 6409 10459 6443
rect 19993 6409 20027 6443
rect 24317 6409 24351 6443
rect 31309 6409 31343 6443
rect 23213 6341 23247 6375
rect 23765 6341 23799 6375
rect 25329 6341 25363 6375
rect 25881 6341 25915 6375
rect 27261 6341 27295 6375
rect 27353 6341 27387 6375
rect 28549 6341 28583 6375
rect 29101 6341 29135 6375
rect 1961 6273 1995 6307
rect 19073 6273 19107 6307
rect 19901 6273 19935 6307
rect 22017 6273 22051 6307
rect 24225 6273 24259 6307
rect 30205 6273 30239 6307
rect 38301 6273 38335 6307
rect 3985 6205 4019 6239
rect 4261 6205 4295 6239
rect 8677 6205 8711 6239
rect 8953 6205 8987 6239
rect 17969 6205 18003 6239
rect 18153 6205 18187 6239
rect 21005 6205 21039 6239
rect 23121 6205 23155 6239
rect 25237 6205 25271 6239
rect 28457 6205 28491 6239
rect 30665 6205 30699 6239
rect 30849 6205 30883 6239
rect 5733 6137 5767 6171
rect 22109 6137 22143 6171
rect 27813 6137 27847 6171
rect 30021 6137 30055 6171
rect 18613 6069 18647 6103
rect 19165 6069 19199 6103
rect 38117 6069 38151 6103
rect 1593 5865 1627 5899
rect 5733 5865 5767 5899
rect 13185 5865 13219 5899
rect 16392 5865 16426 5899
rect 22109 5865 22143 5899
rect 25237 5865 25271 5899
rect 26065 5865 26099 5899
rect 27629 5865 27663 5899
rect 28825 5865 28859 5899
rect 30021 5865 30055 5899
rect 30941 5865 30975 5899
rect 24685 5797 24719 5831
rect 22753 5729 22787 5763
rect 28181 5729 28215 5763
rect 1777 5661 1811 5695
rect 3985 5661 4019 5695
rect 11437 5661 11471 5695
rect 16129 5661 16163 5695
rect 22017 5661 22051 5695
rect 22661 5661 22695 5695
rect 23305 5661 23339 5695
rect 24593 5661 24627 5695
rect 25421 5661 25455 5695
rect 25973 5661 26007 5695
rect 27537 5661 27571 5695
rect 29009 5661 29043 5695
rect 30205 5661 30239 5695
rect 30849 5661 30883 5695
rect 4261 5593 4295 5627
rect 11713 5593 11747 5627
rect 18153 5593 18187 5627
rect 20913 5593 20947 5627
rect 21005 5593 21039 5627
rect 21557 5593 21591 5627
rect 23397 5593 23431 5627
rect 21373 5321 21407 5355
rect 23397 5321 23431 5355
rect 25881 5321 25915 5355
rect 27169 5321 27203 5355
rect 29837 5321 29871 5355
rect 14289 5253 14323 5287
rect 1593 5185 1627 5219
rect 2329 5185 2363 5219
rect 3709 5185 3743 5219
rect 9229 5185 9263 5219
rect 14002 5185 14036 5219
rect 17141 5185 17175 5219
rect 21281 5185 21315 5219
rect 22109 5185 22143 5219
rect 23305 5185 23339 5219
rect 23949 5185 23983 5219
rect 24593 5185 24627 5219
rect 26065 5185 26099 5219
rect 27353 5185 27387 5219
rect 27997 5185 28031 5219
rect 28457 5185 28491 5219
rect 29745 5185 29779 5219
rect 30573 5185 30607 5219
rect 31217 5185 31251 5219
rect 3985 5117 4019 5151
rect 9505 5117 9539 5151
rect 10977 5117 11011 5151
rect 17969 5117 18003 5151
rect 18245 5117 18279 5151
rect 25237 5117 25271 5151
rect 28549 5117 28583 5151
rect 5457 5049 5491 5083
rect 22201 5049 22235 5083
rect 30389 5049 30423 5083
rect 1777 4981 1811 5015
rect 2421 4981 2455 5015
rect 15761 4981 15795 5015
rect 16957 4981 16991 5015
rect 19717 4981 19751 5015
rect 24041 4981 24075 5015
rect 24685 4981 24719 5015
rect 27813 4981 27847 5015
rect 31033 4981 31067 5015
rect 12265 4777 12299 4811
rect 16957 4777 16991 4811
rect 26341 4777 26375 4811
rect 16037 4709 16071 4743
rect 18245 4709 18279 4743
rect 21465 4709 21499 4743
rect 24041 4709 24075 4743
rect 25605 4709 25639 4743
rect 27353 4709 27387 4743
rect 28273 4709 28307 4743
rect 4261 4641 4295 4675
rect 6009 4641 6043 4675
rect 23397 4641 23431 4675
rect 25421 4641 25455 4675
rect 28089 4641 28123 4675
rect 3985 4573 4019 4607
rect 10517 4573 10551 4607
rect 14289 4573 14323 4607
rect 16865 4573 16899 4607
rect 17509 4573 17543 4607
rect 18153 4573 18187 4607
rect 20453 4573 20487 4607
rect 21373 4573 21407 4607
rect 22017 4573 22051 4607
rect 23581 4573 23615 4607
rect 24593 4573 24627 4607
rect 25237 4573 25271 4607
rect 26525 4573 26559 4607
rect 27261 4573 27295 4607
rect 27905 4573 27939 4607
rect 29009 4573 29043 4607
rect 38025 4573 38059 4607
rect 10793 4505 10827 4539
rect 14565 4505 14599 4539
rect 20545 4505 20579 4539
rect 24685 4505 24719 4539
rect 17601 4437 17635 4471
rect 22109 4437 22143 4471
rect 29101 4437 29135 4471
rect 38209 4437 38243 4471
rect 16957 4233 16991 4267
rect 25789 4233 25823 4267
rect 28181 4233 28215 4267
rect 1777 4097 1811 4131
rect 8309 4097 8343 4131
rect 8401 4097 8435 4131
rect 16865 4097 16899 4131
rect 17785 4097 17819 4131
rect 20085 4097 20119 4131
rect 20177 4097 20211 4131
rect 21281 4097 21315 4131
rect 22017 4097 22051 4131
rect 22661 4097 22695 4131
rect 23305 4097 23339 4131
rect 24501 4097 24535 4131
rect 24593 4097 24627 4131
rect 25329 4097 25363 4131
rect 25973 4097 26007 4131
rect 26617 4097 26651 4131
rect 27353 4097 27387 4131
rect 28181 4097 28215 4131
rect 28733 4097 28767 4131
rect 28825 4097 28859 4131
rect 29561 4097 29595 4131
rect 30113 4097 30147 4131
rect 12725 4029 12759 4063
rect 13001 4029 13035 4063
rect 18061 4029 18095 4063
rect 19533 4029 19567 4063
rect 30757 4029 30791 4063
rect 1593 3961 1627 3995
rect 21373 3961 21407 3995
rect 25145 3961 25179 3995
rect 26433 3961 26467 3995
rect 27169 3961 27203 3995
rect 14473 3893 14507 3927
rect 22109 3893 22143 3927
rect 22753 3893 22787 3927
rect 23397 3893 23431 3927
rect 29377 3893 29411 3927
rect 30205 3893 30239 3927
rect 1593 3689 1627 3723
rect 17877 3689 17911 3723
rect 25881 3689 25915 3723
rect 26709 3689 26743 3723
rect 30849 3689 30883 3723
rect 38117 3689 38151 3723
rect 6745 3621 6779 3655
rect 4997 3553 5031 3587
rect 15117 3553 15151 3587
rect 25697 3553 25731 3587
rect 30665 3553 30699 3587
rect 1777 3485 1811 3519
rect 15025 3485 15059 3519
rect 17141 3485 17175 3519
rect 17785 3485 17819 3519
rect 18705 3481 18739 3515
rect 19901 3485 19935 3519
rect 20545 3485 20579 3519
rect 21189 3485 21223 3519
rect 22385 3485 22419 3519
rect 22661 3485 22695 3519
rect 24593 3485 24627 3519
rect 25521 3485 25555 3519
rect 26617 3485 26651 3519
rect 27261 3485 27295 3519
rect 28089 3485 28123 3519
rect 29745 3485 29779 3519
rect 30481 3485 30515 3519
rect 31769 3485 31803 3519
rect 32229 3485 32263 3519
rect 38301 3485 38335 3519
rect 5273 3417 5307 3451
rect 20637 3417 20671 3451
rect 23397 3417 23431 3451
rect 23489 3417 23523 3451
rect 24041 3417 24075 3451
rect 32321 3417 32355 3451
rect 17233 3349 17267 3383
rect 18521 3349 18555 3383
rect 19993 3349 20027 3383
rect 21281 3349 21315 3383
rect 24685 3349 24719 3383
rect 27353 3349 27387 3383
rect 27905 3349 27939 3383
rect 28549 3349 28583 3383
rect 29837 3349 29871 3383
rect 31585 3349 31619 3383
rect 2329 3145 2363 3179
rect 5917 3145 5951 3179
rect 13461 3145 13495 3179
rect 20637 3145 20671 3179
rect 23305 3145 23339 3179
rect 27813 3145 27847 3179
rect 31033 3145 31067 3179
rect 36737 3145 36771 3179
rect 7205 3077 7239 3111
rect 11161 3077 11195 3111
rect 11989 3077 12023 3111
rect 14381 3077 14415 3111
rect 18245 3077 18279 3111
rect 21373 3077 21407 3111
rect 22201 3077 22235 3111
rect 22753 3077 22787 3111
rect 25145 3077 25179 3111
rect 28825 3077 28859 3111
rect 30021 3077 30055 3111
rect 1593 3009 1627 3043
rect 2513 3009 2547 3043
rect 3341 3009 3375 3043
rect 4169 3009 4203 3043
rect 6929 3009 6963 3043
rect 9137 3009 9171 3043
rect 14105 3009 14139 3043
rect 18153 3009 18187 3043
rect 18889 3009 18923 3043
rect 21281 3009 21315 3043
rect 23213 3009 23247 3043
rect 24133 3009 24167 3043
rect 24593 3009 24627 3043
rect 25053 3009 25087 3043
rect 26065 3009 26099 3043
rect 27169 3009 27203 3043
rect 27353 3009 27387 3043
rect 31217 3009 31251 3043
rect 32505 3009 32539 3043
rect 36921 3009 36955 3043
rect 38025 3009 38059 3043
rect 4445 2941 4479 2975
rect 9413 2941 9447 2975
rect 11713 2941 11747 2975
rect 16129 2941 16163 2975
rect 19165 2941 19199 2975
rect 22109 2941 22143 2975
rect 23949 2941 23983 2975
rect 28733 2941 28767 2975
rect 29009 2941 29043 2975
rect 29929 2941 29963 2975
rect 30481 2873 30515 2907
rect 1777 2805 1811 2839
rect 3157 2805 3191 2839
rect 8677 2805 8711 2839
rect 26065 2805 26099 2839
rect 32321 2805 32355 2839
rect 38209 2805 38243 2839
rect 2605 2601 2639 2635
rect 3249 2601 3283 2635
rect 14289 2601 14323 2635
rect 20269 2601 20303 2635
rect 22201 2601 22235 2635
rect 23029 2601 23063 2635
rect 25881 2601 25915 2635
rect 28549 2601 28583 2635
rect 29745 2601 29779 2635
rect 30481 2601 30515 2635
rect 33701 2601 33735 2635
rect 5733 2533 5767 2567
rect 23581 2533 23615 2567
rect 27905 2533 27939 2567
rect 33057 2533 33091 2567
rect 34897 2533 34931 2567
rect 3985 2465 4019 2499
rect 4261 2465 4295 2499
rect 1593 2397 1627 2431
rect 2789 2397 2823 2431
rect 3433 2397 3467 2431
rect 6561 2397 6595 2431
rect 7757 2397 7791 2431
rect 9137 2397 9171 2431
rect 10425 2397 10459 2431
rect 11897 2397 11931 2431
rect 14473 2397 14507 2431
rect 15117 2397 15151 2431
rect 17049 2397 17083 2431
rect 18153 2397 18187 2431
rect 19441 2397 19475 2431
rect 20177 2397 20211 2431
rect 21465 2397 21499 2431
rect 22385 2397 22419 2431
rect 22937 2397 22971 2431
rect 23765 2397 23799 2431
rect 24593 2397 24627 2431
rect 26065 2397 26099 2431
rect 27169 2397 27203 2431
rect 28089 2397 28123 2431
rect 28733 2397 28767 2431
rect 29929 2397 29963 2431
rect 30389 2397 30423 2431
rect 31217 2397 31251 2431
rect 32321 2397 32355 2431
rect 33241 2397 33275 2431
rect 33885 2397 33919 2431
rect 35081 2397 35115 2431
rect 36369 2397 36403 2431
rect 38025 2397 38059 2431
rect 1777 2261 1811 2295
rect 6745 2261 6779 2295
rect 7573 2261 7607 2295
rect 9321 2261 9355 2295
rect 10609 2261 10643 2295
rect 11713 2261 11747 2295
rect 14933 2261 14967 2295
rect 16865 2261 16899 2295
rect 18337 2261 18371 2295
rect 19625 2261 19659 2295
rect 21281 2261 21315 2295
rect 24777 2261 24811 2295
rect 27353 2261 27387 2295
rect 31033 2261 31067 2295
rect 32505 2261 32539 2295
rect 36185 2261 36219 2295
rect 38209 2261 38243 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 37458 37312 37464 37324
rect 10336 37284 10548 37312
rect 37419 37284 37464 37312
rect 1581 37247 1639 37253
rect 1581 37213 1593 37247
rect 1627 37213 1639 37247
rect 1581 37207 1639 37213
rect 2501 37247 2559 37253
rect 2501 37213 2513 37247
rect 2547 37244 2559 37247
rect 2774 37244 2780 37256
rect 2547 37216 2780 37244
rect 2547 37213 2559 37216
rect 2501 37207 2559 37213
rect 1596 37176 1624 37207
rect 2774 37204 2780 37216
rect 2832 37204 2838 37256
rect 3142 37244 3148 37256
rect 3103 37216 3148 37244
rect 3142 37204 3148 37216
rect 3200 37204 3206 37256
rect 3234 37204 3240 37256
rect 3292 37244 3298 37256
rect 4157 37247 4215 37253
rect 4157 37244 4169 37247
rect 3292 37216 4169 37244
rect 3292 37204 3298 37216
rect 4157 37213 4169 37216
rect 4203 37213 4215 37247
rect 4157 37207 4215 37213
rect 4614 37204 4620 37256
rect 4672 37244 4678 37256
rect 4801 37247 4859 37253
rect 4801 37244 4813 37247
rect 4672 37216 4813 37244
rect 4672 37204 4678 37216
rect 4801 37213 4813 37216
rect 4847 37213 4859 37247
rect 4801 37207 4859 37213
rect 6549 37247 6607 37253
rect 6549 37213 6561 37247
rect 6595 37244 6607 37247
rect 7834 37244 7840 37256
rect 6595 37216 6914 37244
rect 7795 37216 7840 37244
rect 6595 37213 6607 37216
rect 6549 37207 6607 37213
rect 4062 37176 4068 37188
rect 1596 37148 4068 37176
rect 4062 37136 4068 37148
rect 4120 37136 4126 37188
rect 6886 37176 6914 37216
rect 7834 37204 7840 37216
rect 7892 37204 7898 37256
rect 9030 37204 9036 37256
rect 9088 37244 9094 37256
rect 9309 37247 9367 37253
rect 9309 37244 9321 37247
rect 9088 37216 9321 37244
rect 9088 37204 9094 37216
rect 9309 37213 9321 37216
rect 9355 37213 9367 37247
rect 9309 37207 9367 37213
rect 10336 37176 10364 37284
rect 10413 37247 10471 37253
rect 10413 37213 10425 37247
rect 10459 37213 10471 37247
rect 10520 37244 10548 37284
rect 37458 37272 37464 37284
rect 37516 37272 37522 37324
rect 11238 37244 11244 37256
rect 10520 37216 11244 37244
rect 10413 37207 10471 37213
rect 6886 37148 10364 37176
rect 10428 37176 10456 37207
rect 11238 37204 11244 37216
rect 11296 37204 11302 37256
rect 11698 37204 11704 37256
rect 11756 37244 11762 37256
rect 12345 37247 12403 37253
rect 12345 37244 12357 37247
rect 11756 37216 12357 37244
rect 11756 37204 11762 37216
rect 12345 37213 12357 37216
rect 12391 37213 12403 37247
rect 12345 37207 12403 37213
rect 13538 37204 13544 37256
rect 13596 37244 13602 37256
rect 14461 37247 14519 37253
rect 14461 37244 14473 37247
rect 13596 37216 14473 37244
rect 13596 37204 13602 37216
rect 14461 37213 14473 37216
rect 14507 37213 14519 37247
rect 15562 37244 15568 37256
rect 15523 37216 15568 37244
rect 14461 37207 14519 37213
rect 15562 37204 15568 37216
rect 15620 37204 15626 37256
rect 16850 37244 16856 37256
rect 16811 37216 16856 37244
rect 16850 37204 16856 37216
rect 16908 37204 16914 37256
rect 18046 37204 18052 37256
rect 18104 37244 18110 37256
rect 18325 37247 18383 37253
rect 18325 37244 18337 37247
rect 18104 37216 18337 37244
rect 18104 37204 18110 37216
rect 18325 37213 18337 37216
rect 18371 37213 18383 37247
rect 18325 37207 18383 37213
rect 20073 37247 20131 37253
rect 20073 37213 20085 37247
rect 20119 37213 20131 37247
rect 22002 37244 22008 37256
rect 21963 37216 22008 37244
rect 20073 37207 20131 37213
rect 13722 37176 13728 37188
rect 10428 37148 13728 37176
rect 13722 37136 13728 37148
rect 13780 37136 13786 37188
rect 17494 37136 17500 37188
rect 17552 37176 17558 37188
rect 20088 37176 20116 37207
rect 22002 37204 22008 37216
rect 22060 37204 22066 37256
rect 22554 37204 22560 37256
rect 22612 37244 22618 37256
rect 22925 37247 22983 37253
rect 22925 37244 22937 37247
rect 22612 37216 22937 37244
rect 22612 37204 22618 37216
rect 22925 37213 22937 37216
rect 22971 37213 22983 37247
rect 22925 37207 22983 37213
rect 24486 37204 24492 37256
rect 24544 37244 24550 37256
rect 24765 37247 24823 37253
rect 24765 37244 24777 37247
rect 24544 37216 24777 37244
rect 24544 37204 24550 37216
rect 24765 37213 24777 37216
rect 24811 37213 24823 37247
rect 24765 37207 24823 37213
rect 25774 37204 25780 37256
rect 25832 37244 25838 37256
rect 26053 37247 26111 37253
rect 26053 37244 26065 37247
rect 25832 37216 26065 37244
rect 25832 37204 25838 37216
rect 26053 37213 26065 37216
rect 26099 37213 26111 37247
rect 27798 37244 27804 37256
rect 27759 37216 27804 37244
rect 26053 37207 26111 37213
rect 27798 37204 27804 37216
rect 27856 37204 27862 37256
rect 28626 37204 28632 37256
rect 28684 37244 28690 37256
rect 29733 37247 29791 37253
rect 29733 37244 29745 37247
rect 28684 37216 29745 37244
rect 28684 37204 28690 37216
rect 29733 37213 29745 37216
rect 29779 37213 29791 37247
rect 29733 37207 29791 37213
rect 30374 37204 30380 37256
rect 30432 37244 30438 37256
rect 30653 37247 30711 37253
rect 30653 37244 30665 37247
rect 30432 37216 30665 37244
rect 30432 37204 30438 37216
rect 30653 37213 30665 37216
rect 30699 37213 30711 37247
rect 30653 37207 30711 37213
rect 32214 37204 32220 37256
rect 32272 37244 32278 37256
rect 32493 37247 32551 37253
rect 32493 37244 32505 37247
rect 32272 37216 32505 37244
rect 32272 37204 32278 37216
rect 32493 37213 32505 37216
rect 32539 37213 32551 37247
rect 32493 37207 32551 37213
rect 33502 37204 33508 37256
rect 33560 37244 33566 37256
rect 33781 37247 33839 37253
rect 33781 37244 33793 37247
rect 33560 37216 33793 37244
rect 33560 37204 33566 37216
rect 33781 37213 33793 37216
rect 33827 37213 33839 37247
rect 33781 37207 33839 37213
rect 33870 37204 33876 37256
rect 33928 37244 33934 37256
rect 34885 37247 34943 37253
rect 34885 37244 34897 37247
rect 33928 37216 34897 37244
rect 33928 37204 33934 37216
rect 34885 37213 34897 37216
rect 34931 37213 34943 37247
rect 36633 37247 36691 37253
rect 36633 37244 36645 37247
rect 34885 37207 34943 37213
rect 35866 37216 36645 37244
rect 17552 37148 20116 37176
rect 17552 37136 17558 37148
rect 28902 37136 28908 37188
rect 28960 37176 28966 37188
rect 28960 37148 30512 37176
rect 28960 37136 28966 37148
rect 1302 37068 1308 37120
rect 1360 37108 1366 37120
rect 1765 37111 1823 37117
rect 1765 37108 1777 37111
rect 1360 37080 1777 37108
rect 1360 37068 1366 37080
rect 1765 37077 1777 37080
rect 1811 37077 1823 37111
rect 2314 37108 2320 37120
rect 2275 37080 2320 37108
rect 1765 37071 1823 37077
rect 2314 37068 2320 37080
rect 2372 37068 2378 37120
rect 2958 37108 2964 37120
rect 2919 37080 2964 37108
rect 2958 37068 2964 37080
rect 3016 37068 3022 37120
rect 3970 37108 3976 37120
rect 3931 37080 3976 37108
rect 3970 37068 3976 37080
rect 4028 37068 4034 37120
rect 4614 37108 4620 37120
rect 4575 37080 4620 37108
rect 4614 37068 4620 37080
rect 4672 37068 4678 37120
rect 5810 37068 5816 37120
rect 5868 37108 5874 37120
rect 6733 37111 6791 37117
rect 6733 37108 6745 37111
rect 5868 37080 6745 37108
rect 5868 37068 5874 37080
rect 6733 37077 6745 37080
rect 6779 37077 6791 37111
rect 6733 37071 6791 37077
rect 7742 37068 7748 37120
rect 7800 37108 7806 37120
rect 8021 37111 8079 37117
rect 8021 37108 8033 37111
rect 7800 37080 8033 37108
rect 7800 37068 7806 37080
rect 8021 37077 8033 37080
rect 8067 37077 8079 37111
rect 8021 37071 8079 37077
rect 8938 37068 8944 37120
rect 8996 37108 9002 37120
rect 9125 37111 9183 37117
rect 9125 37108 9137 37111
rect 8996 37080 9137 37108
rect 8996 37068 9002 37080
rect 9125 37077 9137 37080
rect 9171 37077 9183 37111
rect 9125 37071 9183 37077
rect 10318 37068 10324 37120
rect 10376 37108 10382 37120
rect 10597 37111 10655 37117
rect 10597 37108 10609 37111
rect 10376 37080 10609 37108
rect 10376 37068 10382 37080
rect 10597 37077 10609 37080
rect 10643 37077 10655 37111
rect 10597 37071 10655 37077
rect 12434 37068 12440 37120
rect 12492 37108 12498 37120
rect 12529 37111 12587 37117
rect 12529 37108 12541 37111
rect 12492 37080 12541 37108
rect 12492 37068 12498 37080
rect 12529 37077 12541 37080
rect 12575 37077 12587 37111
rect 14274 37108 14280 37120
rect 14235 37080 14280 37108
rect 12529 37071 12587 37077
rect 14274 37068 14280 37080
rect 14332 37068 14338 37120
rect 15470 37068 15476 37120
rect 15528 37108 15534 37120
rect 15749 37111 15807 37117
rect 15749 37108 15761 37111
rect 15528 37080 15761 37108
rect 15528 37068 15534 37080
rect 15749 37077 15761 37080
rect 15795 37077 15807 37111
rect 15749 37071 15807 37077
rect 16758 37068 16764 37120
rect 16816 37108 16822 37120
rect 17037 37111 17095 37117
rect 17037 37108 17049 37111
rect 16816 37080 17049 37108
rect 16816 37068 16822 37080
rect 17037 37077 17049 37080
rect 17083 37077 17095 37111
rect 17037 37071 17095 37077
rect 17954 37068 17960 37120
rect 18012 37108 18018 37120
rect 18141 37111 18199 37117
rect 18141 37108 18153 37111
rect 18012 37080 18153 37108
rect 18012 37068 18018 37080
rect 18141 37077 18153 37080
rect 18187 37077 18199 37111
rect 18141 37071 18199 37077
rect 19978 37068 19984 37120
rect 20036 37108 20042 37120
rect 20257 37111 20315 37117
rect 20257 37108 20269 37111
rect 20036 37080 20269 37108
rect 20036 37068 20042 37080
rect 20257 37077 20269 37080
rect 20303 37077 20315 37111
rect 20257 37071 20315 37077
rect 21266 37068 21272 37120
rect 21324 37108 21330 37120
rect 22189 37111 22247 37117
rect 22189 37108 22201 37111
rect 21324 37080 22201 37108
rect 21324 37068 21330 37080
rect 22189 37077 22201 37080
rect 22235 37077 22247 37111
rect 22738 37108 22744 37120
rect 22699 37080 22744 37108
rect 22189 37071 22247 37077
rect 22738 37068 22744 37080
rect 22796 37068 22802 37120
rect 23106 37068 23112 37120
rect 23164 37108 23170 37120
rect 24581 37111 24639 37117
rect 24581 37108 24593 37111
rect 23164 37080 24593 37108
rect 23164 37068 23170 37080
rect 24581 37077 24593 37080
rect 24627 37077 24639 37111
rect 24581 37071 24639 37077
rect 25130 37068 25136 37120
rect 25188 37108 25194 37120
rect 25869 37111 25927 37117
rect 25869 37108 25881 37111
rect 25188 37080 25881 37108
rect 25188 37068 25194 37080
rect 25869 37077 25881 37080
rect 25915 37077 25927 37111
rect 25869 37071 25927 37077
rect 27706 37068 27712 37120
rect 27764 37108 27770 37120
rect 27985 37111 28043 37117
rect 27985 37108 27997 37111
rect 27764 37080 27997 37108
rect 27764 37068 27770 37080
rect 27985 37077 27997 37080
rect 28031 37077 28043 37111
rect 27985 37071 28043 37077
rect 28994 37068 29000 37120
rect 29052 37108 29058 37120
rect 30484 37117 30512 37148
rect 32122 37136 32128 37188
rect 32180 37176 32186 37188
rect 35866 37176 35894 37216
rect 36633 37213 36645 37216
rect 36679 37213 36691 37247
rect 37734 37244 37740 37256
rect 37695 37216 37740 37244
rect 36633 37207 36691 37213
rect 37734 37204 37740 37216
rect 37792 37204 37798 37256
rect 32180 37148 35894 37176
rect 32180 37136 32186 37148
rect 29917 37111 29975 37117
rect 29917 37108 29929 37111
rect 29052 37080 29929 37108
rect 29052 37068 29058 37080
rect 29917 37077 29929 37080
rect 29963 37077 29975 37111
rect 29917 37071 29975 37077
rect 30469 37111 30527 37117
rect 30469 37077 30481 37111
rect 30515 37077 30527 37111
rect 30469 37071 30527 37077
rect 32309 37111 32367 37117
rect 32309 37077 32321 37111
rect 32355 37108 32367 37111
rect 32398 37108 32404 37120
rect 32355 37080 32404 37108
rect 32355 37077 32367 37080
rect 32309 37071 32367 37077
rect 32398 37068 32404 37080
rect 32456 37068 32462 37120
rect 33318 37068 33324 37120
rect 33376 37108 33382 37120
rect 33597 37111 33655 37117
rect 33597 37108 33609 37111
rect 33376 37080 33609 37108
rect 33376 37068 33382 37080
rect 33597 37077 33609 37080
rect 33643 37077 33655 37111
rect 33597 37071 33655 37077
rect 34790 37068 34796 37120
rect 34848 37108 34854 37120
rect 35069 37111 35127 37117
rect 35069 37108 35081 37111
rect 34848 37080 35081 37108
rect 34848 37068 34854 37080
rect 35069 37077 35081 37080
rect 35115 37077 35127 37111
rect 35069 37071 35127 37077
rect 36722 37068 36728 37120
rect 36780 37108 36786 37120
rect 36817 37111 36875 37117
rect 36817 37108 36829 37111
rect 36780 37080 36829 37108
rect 36780 37068 36786 37080
rect 36817 37077 36829 37080
rect 36863 37077 36875 37111
rect 36817 37071 36875 37077
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 14 36864 20 36916
rect 72 36904 78 36916
rect 1765 36907 1823 36913
rect 1765 36904 1777 36907
rect 72 36876 1777 36904
rect 72 36864 78 36876
rect 1765 36873 1777 36876
rect 1811 36873 1823 36907
rect 1765 36867 1823 36873
rect 4614 36864 4620 36916
rect 4672 36904 4678 36916
rect 10686 36904 10692 36916
rect 4672 36876 10692 36904
rect 4672 36864 4678 36876
rect 10686 36864 10692 36876
rect 10744 36864 10750 36916
rect 15562 36864 15568 36916
rect 15620 36904 15626 36916
rect 18046 36904 18052 36916
rect 15620 36876 18052 36904
rect 15620 36864 15626 36876
rect 18046 36864 18052 36876
rect 18104 36864 18110 36916
rect 38197 36907 38255 36913
rect 38197 36873 38209 36907
rect 38243 36904 38255 36907
rect 39298 36904 39304 36916
rect 38243 36876 39304 36904
rect 38243 36873 38255 36876
rect 38197 36867 38255 36873
rect 39298 36864 39304 36876
rect 39356 36864 39362 36916
rect 2314 36796 2320 36848
rect 2372 36836 2378 36848
rect 7650 36836 7656 36848
rect 2372 36808 7656 36836
rect 2372 36796 2378 36808
rect 7650 36796 7656 36808
rect 7708 36796 7714 36848
rect 1581 36771 1639 36777
rect 1581 36737 1593 36771
rect 1627 36768 1639 36771
rect 4614 36768 4620 36780
rect 1627 36740 4620 36768
rect 1627 36737 1639 36740
rect 1581 36731 1639 36737
rect 4614 36728 4620 36740
rect 4672 36728 4678 36780
rect 36906 36768 36912 36780
rect 36867 36740 36912 36768
rect 36906 36728 36912 36740
rect 36964 36728 36970 36780
rect 36998 36728 37004 36780
rect 37056 36768 37062 36780
rect 38013 36771 38071 36777
rect 38013 36768 38025 36771
rect 37056 36740 38025 36768
rect 37056 36728 37062 36740
rect 38013 36737 38025 36740
rect 38059 36737 38071 36771
rect 38013 36731 38071 36737
rect 36722 36564 36728 36576
rect 36683 36536 36728 36564
rect 36722 36524 36728 36536
rect 36780 36524 36786 36576
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 38010 36116 38016 36168
rect 38068 36156 38074 36168
rect 38289 36159 38347 36165
rect 38289 36156 38301 36159
rect 38068 36128 38301 36156
rect 38068 36116 38074 36128
rect 38289 36125 38301 36128
rect 38335 36125 38347 36159
rect 38289 36119 38347 36125
rect 37274 35980 37280 36032
rect 37332 36020 37338 36032
rect 38105 36023 38163 36029
rect 38105 36020 38117 36023
rect 37332 35992 38117 36020
rect 37332 35980 37338 35992
rect 38105 35989 38117 35992
rect 38151 35989 38163 36023
rect 38105 35983 38163 35989
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 4062 35232 4068 35284
rect 4120 35272 4126 35284
rect 7009 35275 7067 35281
rect 7009 35272 7021 35275
rect 4120 35244 7021 35272
rect 4120 35232 4126 35244
rect 7009 35241 7021 35244
rect 7055 35241 7067 35275
rect 7009 35235 7067 35241
rect 7193 35071 7251 35077
rect 7193 35037 7205 35071
rect 7239 35068 7251 35071
rect 14090 35068 14096 35080
rect 7239 35040 14096 35068
rect 7239 35037 7251 35040
rect 7193 35031 7251 35037
rect 14090 35028 14096 35040
rect 14148 35028 14154 35080
rect 33410 35028 33416 35080
rect 33468 35068 33474 35080
rect 38013 35071 38071 35077
rect 38013 35068 38025 35071
rect 33468 35040 38025 35068
rect 33468 35028 33474 35040
rect 38013 35037 38025 35040
rect 38059 35037 38071 35071
rect 38013 35031 38071 35037
rect 38194 34932 38200 34944
rect 38155 34904 38200 34932
rect 38194 34892 38200 34904
rect 38252 34892 38258 34944
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 31481 34731 31539 34737
rect 31481 34697 31493 34731
rect 31527 34728 31539 34731
rect 32122 34728 32128 34740
rect 31527 34700 32128 34728
rect 31527 34697 31539 34700
rect 31481 34691 31539 34697
rect 32122 34688 32128 34700
rect 32180 34688 32186 34740
rect 32401 34731 32459 34737
rect 32401 34697 32413 34731
rect 32447 34728 32459 34731
rect 33870 34728 33876 34740
rect 32447 34700 33876 34728
rect 32447 34697 32459 34700
rect 32401 34691 32459 34697
rect 33870 34688 33876 34700
rect 33928 34688 33934 34740
rect 31662 34592 31668 34604
rect 31623 34564 31668 34592
rect 31662 34552 31668 34564
rect 31720 34552 31726 34604
rect 32585 34595 32643 34601
rect 32585 34561 32597 34595
rect 32631 34561 32643 34595
rect 32585 34555 32643 34561
rect 28534 34484 28540 34536
rect 28592 34524 28598 34536
rect 32600 34524 32628 34555
rect 28592 34496 32628 34524
rect 28592 34484 28598 34496
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 1762 33504 1768 33516
rect 1723 33476 1768 33504
rect 1762 33464 1768 33476
rect 1820 33464 1826 33516
rect 38286 33504 38292 33516
rect 38247 33476 38292 33504
rect 38286 33464 38292 33476
rect 38344 33464 38350 33516
rect 1581 33303 1639 33309
rect 1581 33269 1593 33303
rect 1627 33300 1639 33303
rect 7190 33300 7196 33312
rect 1627 33272 7196 33300
rect 1627 33269 1639 33272
rect 1581 33263 1639 33269
rect 7190 33260 7196 33272
rect 7248 33260 7254 33312
rect 38102 33300 38108 33312
rect 38063 33272 38108 33300
rect 38102 33260 38108 33272
rect 38160 33260 38166 33312
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 11238 33056 11244 33108
rect 11296 33096 11302 33108
rect 11885 33099 11943 33105
rect 11885 33096 11897 33099
rect 11296 33068 11897 33096
rect 11296 33056 11302 33068
rect 11885 33065 11897 33068
rect 11931 33065 11943 33099
rect 11885 33059 11943 33065
rect 31205 33099 31263 33105
rect 31205 33065 31217 33099
rect 31251 33096 31263 33099
rect 31662 33096 31668 33108
rect 31251 33068 31668 33096
rect 31251 33065 31263 33068
rect 31205 33059 31263 33065
rect 31662 33056 31668 33068
rect 31720 33056 31726 33108
rect 32769 33099 32827 33105
rect 32769 33065 32781 33099
rect 32815 33096 32827 33099
rect 36998 33096 37004 33108
rect 32815 33068 37004 33096
rect 32815 33065 32827 33068
rect 32769 33059 32827 33065
rect 36998 33056 37004 33068
rect 37056 33056 37062 33108
rect 12069 32895 12127 32901
rect 12069 32861 12081 32895
rect 12115 32892 12127 32895
rect 12526 32892 12532 32904
rect 12115 32864 12532 32892
rect 12115 32861 12127 32864
rect 12069 32855 12127 32861
rect 12526 32852 12532 32864
rect 12584 32852 12590 32904
rect 31110 32892 31116 32904
rect 31071 32864 31116 32892
rect 31110 32852 31116 32864
rect 31168 32852 31174 32904
rect 32950 32892 32956 32904
rect 32911 32864 32956 32892
rect 32950 32852 32956 32864
rect 33008 32852 33014 32904
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 4157 32555 4215 32561
rect 4157 32521 4169 32555
rect 4203 32552 4215 32555
rect 4614 32552 4620 32564
rect 4203 32524 4620 32552
rect 4203 32521 4215 32524
rect 4157 32515 4215 32521
rect 4614 32512 4620 32524
rect 4672 32512 4678 32564
rect 11698 32552 11704 32564
rect 11659 32524 11704 32552
rect 11698 32512 11704 32524
rect 11756 32512 11762 32564
rect 17494 32552 17500 32564
rect 17455 32524 17500 32552
rect 17494 32512 17500 32524
rect 17552 32512 17558 32564
rect 28626 32552 28632 32564
rect 28587 32524 28632 32552
rect 28626 32512 28632 32524
rect 28684 32512 28690 32564
rect 1762 32416 1768 32428
rect 1723 32388 1768 32416
rect 1762 32376 1768 32388
rect 1820 32376 1826 32428
rect 4341 32419 4399 32425
rect 4341 32385 4353 32419
rect 4387 32416 4399 32419
rect 4614 32416 4620 32428
rect 4387 32388 4620 32416
rect 4387 32385 4399 32388
rect 4341 32379 4399 32385
rect 4614 32376 4620 32388
rect 4672 32376 4678 32428
rect 11882 32416 11888 32428
rect 11843 32388 11888 32416
rect 11882 32376 11888 32388
rect 11940 32376 11946 32428
rect 16942 32376 16948 32428
rect 17000 32416 17006 32428
rect 17681 32419 17739 32425
rect 17681 32416 17693 32419
rect 17000 32388 17693 32416
rect 17000 32376 17006 32388
rect 17681 32385 17693 32388
rect 17727 32385 17739 32419
rect 28810 32416 28816 32428
rect 28771 32388 28816 32416
rect 17681 32379 17739 32385
rect 28810 32376 28816 32388
rect 28868 32376 28874 32428
rect 35434 32376 35440 32428
rect 35492 32416 35498 32428
rect 38013 32419 38071 32425
rect 38013 32416 38025 32419
rect 35492 32388 38025 32416
rect 35492 32376 35498 32388
rect 38013 32385 38025 32388
rect 38059 32385 38071 32419
rect 38013 32379 38071 32385
rect 1581 32215 1639 32221
rect 1581 32181 1593 32215
rect 1627 32212 1639 32215
rect 6270 32212 6276 32224
rect 1627 32184 6276 32212
rect 1627 32181 1639 32184
rect 1581 32175 1639 32181
rect 6270 32172 6276 32184
rect 6328 32172 6334 32224
rect 38194 32212 38200 32224
rect 38155 32184 38200 32212
rect 38194 32172 38200 32184
rect 38252 32172 38258 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 7834 31968 7840 32020
rect 7892 32008 7898 32020
rect 9953 32011 10011 32017
rect 9953 32008 9965 32011
rect 7892 31980 9965 32008
rect 7892 31968 7898 31980
rect 9953 31977 9965 31980
rect 9999 31977 10011 32011
rect 16850 32008 16856 32020
rect 16811 31980 16856 32008
rect 9953 31971 10011 31977
rect 16850 31968 16856 31980
rect 16908 31968 16914 32020
rect 14274 31900 14280 31952
rect 14332 31940 14338 31952
rect 14332 31912 21404 31940
rect 14332 31900 14338 31912
rect 10137 31807 10195 31813
rect 10137 31773 10149 31807
rect 10183 31804 10195 31807
rect 10594 31804 10600 31816
rect 10183 31776 10600 31804
rect 10183 31773 10195 31776
rect 10137 31767 10195 31773
rect 10594 31764 10600 31776
rect 10652 31764 10658 31816
rect 17034 31804 17040 31816
rect 16995 31776 17040 31804
rect 17034 31764 17040 31776
rect 17092 31764 17098 31816
rect 21376 31804 21404 31912
rect 27522 31832 27528 31884
rect 27580 31872 27586 31884
rect 30009 31875 30067 31881
rect 30009 31872 30021 31875
rect 27580 31844 30021 31872
rect 27580 31832 27586 31844
rect 30009 31841 30021 31844
rect 30055 31841 30067 31875
rect 30009 31835 30067 31841
rect 26973 31807 27031 31813
rect 26973 31804 26985 31807
rect 21376 31776 26985 31804
rect 26973 31773 26985 31776
rect 27019 31773 27031 31807
rect 26973 31767 27031 31773
rect 29917 31807 29975 31813
rect 29917 31773 29929 31807
rect 29963 31804 29975 31807
rect 36722 31804 36728 31816
rect 29963 31776 36728 31804
rect 29963 31773 29975 31776
rect 29917 31767 29975 31773
rect 36722 31764 36728 31776
rect 36780 31764 36786 31816
rect 26786 31668 26792 31680
rect 26747 31640 26792 31668
rect 26786 31628 26792 31640
rect 26844 31628 26850 31680
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 25961 31467 26019 31473
rect 25961 31433 25973 31467
rect 26007 31464 26019 31467
rect 27798 31464 27804 31476
rect 26007 31436 27804 31464
rect 26007 31433 26019 31436
rect 25961 31427 26019 31433
rect 27798 31424 27804 31436
rect 27856 31424 27862 31476
rect 15289 31331 15347 31337
rect 15289 31297 15301 31331
rect 15335 31328 15347 31331
rect 15562 31328 15568 31340
rect 15335 31300 15568 31328
rect 15335 31297 15347 31300
rect 15289 31291 15347 31297
rect 15562 31288 15568 31300
rect 15620 31288 15626 31340
rect 15933 31331 15991 31337
rect 15933 31297 15945 31331
rect 15979 31297 15991 31331
rect 15933 31291 15991 31297
rect 15948 31260 15976 31291
rect 19426 31288 19432 31340
rect 19484 31328 19490 31340
rect 19705 31331 19763 31337
rect 19705 31328 19717 31331
rect 19484 31300 19717 31328
rect 19484 31288 19490 31300
rect 19705 31297 19717 31300
rect 19751 31297 19763 31331
rect 26142 31328 26148 31340
rect 26103 31300 26148 31328
rect 19705 31291 19763 31297
rect 26142 31288 26148 31300
rect 26200 31288 26206 31340
rect 30653 31331 30711 31337
rect 30653 31297 30665 31331
rect 30699 31328 30711 31331
rect 37274 31328 37280 31340
rect 30699 31300 37280 31328
rect 30699 31297 30711 31300
rect 30653 31291 30711 31297
rect 37274 31288 37280 31300
rect 37332 31288 37338 31340
rect 15120 31232 15976 31260
rect 15120 31201 15148 31232
rect 19518 31220 19524 31272
rect 19576 31260 19582 31272
rect 20165 31263 20223 31269
rect 20165 31260 20177 31263
rect 19576 31232 20177 31260
rect 19576 31220 19582 31232
rect 20165 31229 20177 31232
rect 20211 31229 20223 31263
rect 20165 31223 20223 31229
rect 15105 31195 15163 31201
rect 15105 31161 15117 31195
rect 15151 31161 15163 31195
rect 15105 31155 15163 31161
rect 15286 31084 15292 31136
rect 15344 31124 15350 31136
rect 15749 31127 15807 31133
rect 15749 31124 15761 31127
rect 15344 31096 15761 31124
rect 15344 31084 15350 31096
rect 15749 31093 15761 31096
rect 15795 31093 15807 31127
rect 15749 31087 15807 31093
rect 19521 31127 19579 31133
rect 19521 31093 19533 31127
rect 19567 31124 19579 31127
rect 19702 31124 19708 31136
rect 19567 31096 19708 31124
rect 19567 31093 19579 31096
rect 19521 31087 19579 31093
rect 19702 31084 19708 31096
rect 19760 31084 19766 31136
rect 30466 31124 30472 31136
rect 30427 31096 30472 31124
rect 30466 31084 30472 31096
rect 30524 31084 30530 31136
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 13722 30880 13728 30932
rect 13780 30920 13786 30932
rect 14277 30923 14335 30929
rect 14277 30920 14289 30923
rect 13780 30892 14289 30920
rect 13780 30880 13786 30892
rect 14277 30889 14289 30892
rect 14323 30889 14335 30923
rect 14277 30883 14335 30889
rect 17034 30880 17040 30932
rect 17092 30920 17098 30932
rect 17405 30923 17463 30929
rect 17405 30920 17417 30923
rect 17092 30892 17417 30920
rect 17092 30880 17098 30892
rect 17405 30889 17417 30892
rect 17451 30889 17463 30923
rect 18046 30920 18052 30932
rect 18007 30892 18052 30920
rect 17405 30883 17463 30889
rect 18046 30880 18052 30892
rect 18104 30880 18110 30932
rect 19518 30784 19524 30796
rect 19479 30756 19524 30784
rect 19518 30744 19524 30756
rect 19576 30744 19582 30796
rect 19702 30784 19708 30796
rect 19663 30756 19708 30784
rect 19702 30744 19708 30756
rect 19760 30744 19766 30796
rect 23293 30787 23351 30793
rect 23293 30753 23305 30787
rect 23339 30784 23351 30787
rect 27522 30784 27528 30796
rect 23339 30756 27528 30784
rect 23339 30753 23351 30756
rect 23293 30747 23351 30753
rect 27522 30744 27528 30756
rect 27580 30744 27586 30796
rect 1578 30716 1584 30728
rect 1539 30688 1584 30716
rect 1578 30676 1584 30688
rect 1636 30676 1642 30728
rect 1854 30716 1860 30728
rect 1815 30688 1860 30716
rect 1854 30676 1860 30688
rect 1912 30676 1918 30728
rect 11238 30716 11244 30728
rect 11199 30688 11244 30716
rect 11238 30676 11244 30688
rect 11296 30676 11302 30728
rect 11885 30719 11943 30725
rect 11885 30685 11897 30719
rect 11931 30685 11943 30719
rect 14458 30716 14464 30728
rect 14419 30688 14464 30716
rect 11885 30679 11943 30685
rect 11900 30648 11928 30679
rect 14458 30676 14464 30688
rect 14516 30676 14522 30728
rect 17313 30719 17371 30725
rect 17313 30685 17325 30719
rect 17359 30685 17371 30719
rect 17313 30679 17371 30685
rect 18233 30719 18291 30725
rect 18233 30685 18245 30719
rect 18279 30716 18291 30719
rect 19978 30716 19984 30728
rect 18279 30688 19984 30716
rect 18279 30685 18291 30688
rect 18233 30679 18291 30685
rect 11072 30620 11928 30648
rect 17328 30648 17356 30679
rect 19978 30676 19984 30688
rect 20036 30676 20042 30728
rect 22554 30716 22560 30728
rect 22515 30688 22560 30716
rect 22554 30676 22560 30688
rect 22612 30676 22618 30728
rect 33318 30716 33324 30728
rect 33279 30688 33324 30716
rect 33318 30676 33324 30688
rect 33376 30676 33382 30728
rect 18874 30648 18880 30660
rect 17328 30620 18880 30648
rect 11072 30589 11100 30620
rect 18874 30608 18880 30620
rect 18932 30608 18938 30660
rect 23385 30651 23443 30657
rect 23385 30617 23397 30651
rect 23431 30617 23443 30651
rect 23385 30611 23443 30617
rect 23937 30651 23995 30657
rect 23937 30617 23949 30651
rect 23983 30648 23995 30651
rect 24026 30648 24032 30660
rect 23983 30620 24032 30648
rect 23983 30617 23995 30620
rect 23937 30611 23995 30617
rect 11057 30583 11115 30589
rect 11057 30549 11069 30583
rect 11103 30549 11115 30583
rect 11057 30543 11115 30549
rect 11701 30583 11759 30589
rect 11701 30549 11713 30583
rect 11747 30580 11759 30583
rect 11974 30580 11980 30592
rect 11747 30552 11980 30580
rect 11747 30549 11759 30552
rect 11701 30543 11759 30549
rect 11974 30540 11980 30552
rect 12032 30540 12038 30592
rect 20162 30580 20168 30592
rect 20123 30552 20168 30580
rect 20162 30540 20168 30552
rect 20220 30540 20226 30592
rect 22649 30583 22707 30589
rect 22649 30549 22661 30583
rect 22695 30580 22707 30583
rect 23400 30580 23428 30611
rect 24026 30608 24032 30620
rect 24084 30608 24090 30660
rect 22695 30552 23428 30580
rect 22695 30549 22707 30552
rect 22649 30543 22707 30549
rect 31754 30540 31760 30592
rect 31812 30580 31818 30592
rect 33413 30583 33471 30589
rect 33413 30580 33425 30583
rect 31812 30552 33425 30580
rect 31812 30540 31818 30552
rect 33413 30549 33425 30552
rect 33459 30549 33471 30583
rect 33413 30543 33471 30549
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 14458 30336 14464 30388
rect 14516 30376 14522 30388
rect 14921 30379 14979 30385
rect 14921 30376 14933 30379
rect 14516 30348 14933 30376
rect 14516 30336 14522 30348
rect 14921 30345 14933 30348
rect 14967 30345 14979 30379
rect 14921 30339 14979 30345
rect 19426 30336 19432 30388
rect 19484 30376 19490 30388
rect 19521 30379 19579 30385
rect 19521 30376 19533 30379
rect 19484 30348 19533 30376
rect 19484 30336 19490 30348
rect 19521 30345 19533 30348
rect 19567 30345 19579 30379
rect 22554 30376 22560 30388
rect 19521 30339 19579 30345
rect 22066 30348 22560 30376
rect 10594 30308 10600 30320
rect 10555 30280 10600 30308
rect 10594 30268 10600 30280
rect 10652 30268 10658 30320
rect 12526 30308 12532 30320
rect 12487 30280 12532 30308
rect 12526 30268 12532 30280
rect 12584 30268 12590 30320
rect 14090 30268 14096 30320
rect 14148 30308 14154 30320
rect 14277 30311 14335 30317
rect 14277 30308 14289 30311
rect 14148 30280 14289 30308
rect 14148 30268 14154 30280
rect 14277 30277 14289 30280
rect 14323 30277 14335 30311
rect 16942 30308 16948 30320
rect 16903 30280 16948 30308
rect 14277 30271 14335 30277
rect 16942 30268 16948 30280
rect 17000 30268 17006 30320
rect 10505 30243 10563 30249
rect 10505 30209 10517 30243
rect 10551 30240 10563 30243
rect 12250 30240 12256 30252
rect 10551 30212 12256 30240
rect 10551 30209 10563 30212
rect 10505 30203 10563 30209
rect 12250 30200 12256 30212
rect 12308 30200 12314 30252
rect 12434 30200 12440 30252
rect 12492 30240 12498 30252
rect 14182 30240 14188 30252
rect 12492 30212 12537 30240
rect 14143 30212 14188 30240
rect 12492 30200 12498 30212
rect 14182 30200 14188 30212
rect 14240 30200 14246 30252
rect 14829 30243 14887 30249
rect 14829 30209 14841 30243
rect 14875 30240 14887 30243
rect 15010 30240 15016 30252
rect 14875 30212 15016 30240
rect 14875 30209 14887 30212
rect 14829 30203 14887 30209
rect 15010 30200 15016 30212
rect 15068 30200 15074 30252
rect 16850 30240 16856 30252
rect 16811 30212 16856 30240
rect 16850 30200 16856 30212
rect 16908 30200 16914 30252
rect 19242 30200 19248 30252
rect 19300 30240 19306 30252
rect 19705 30243 19763 30249
rect 19705 30240 19717 30243
rect 19300 30212 19717 30240
rect 19300 30200 19306 30212
rect 19705 30209 19717 30212
rect 19751 30240 19763 30243
rect 22066 30240 22094 30348
rect 22554 30336 22560 30348
rect 22612 30376 22618 30388
rect 24946 30376 24952 30388
rect 22612 30348 24952 30376
rect 22612 30336 22618 30348
rect 24946 30336 24952 30348
rect 25004 30336 25010 30388
rect 28905 30311 28963 30317
rect 28905 30277 28917 30311
rect 28951 30308 28963 30311
rect 32950 30308 32956 30320
rect 28951 30280 32956 30308
rect 28951 30277 28963 30280
rect 28905 30271 28963 30277
rect 32950 30268 32956 30280
rect 33008 30268 33014 30320
rect 23106 30240 23112 30252
rect 19751 30212 22094 30240
rect 23067 30212 23112 30240
rect 19751 30209 19763 30212
rect 19705 30203 19763 30209
rect 23106 30200 23112 30212
rect 23164 30200 23170 30252
rect 24762 30200 24768 30252
rect 24820 30240 24826 30252
rect 28813 30243 28871 30249
rect 28813 30240 28825 30243
rect 24820 30212 28825 30240
rect 24820 30200 24826 30212
rect 28813 30209 28825 30212
rect 28859 30209 28871 30243
rect 33594 30240 33600 30252
rect 33555 30212 33600 30240
rect 28813 30203 28871 30209
rect 33594 30200 33600 30212
rect 33652 30200 33658 30252
rect 38013 30243 38071 30249
rect 38013 30240 38025 30243
rect 35866 30212 38025 30240
rect 5166 30132 5172 30184
rect 5224 30172 5230 30184
rect 7101 30175 7159 30181
rect 7101 30172 7113 30175
rect 5224 30144 7113 30172
rect 5224 30132 5230 30144
rect 7101 30141 7113 30144
rect 7147 30141 7159 30175
rect 7282 30172 7288 30184
rect 7243 30144 7288 30172
rect 7101 30135 7159 30141
rect 7282 30132 7288 30144
rect 7340 30132 7346 30184
rect 33318 30132 33324 30184
rect 33376 30172 33382 30184
rect 35866 30172 35894 30212
rect 38013 30209 38025 30212
rect 38059 30209 38071 30243
rect 38013 30203 38071 30209
rect 33376 30144 35894 30172
rect 33376 30132 33382 30144
rect 33410 30104 33416 30116
rect 33371 30076 33416 30104
rect 33410 30064 33416 30076
rect 33468 30064 33474 30116
rect 7745 30039 7803 30045
rect 7745 30005 7757 30039
rect 7791 30036 7803 30039
rect 8662 30036 8668 30048
rect 7791 30008 8668 30036
rect 7791 30005 7803 30008
rect 7745 29999 7803 30005
rect 8662 29996 8668 30008
rect 8720 29996 8726 30048
rect 23198 30036 23204 30048
rect 23159 30008 23204 30036
rect 23198 29996 23204 30008
rect 23256 29996 23262 30048
rect 38194 30036 38200 30048
rect 38155 30008 38200 30036
rect 38194 29996 38200 30008
rect 38252 29996 38258 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 5166 29832 5172 29844
rect 5127 29804 5172 29832
rect 5166 29792 5172 29804
rect 5224 29792 5230 29844
rect 7282 29832 7288 29844
rect 7243 29804 7288 29832
rect 7282 29792 7288 29804
rect 7340 29792 7346 29844
rect 11241 29835 11299 29841
rect 11241 29801 11253 29835
rect 11287 29832 11299 29835
rect 11882 29832 11888 29844
rect 11287 29804 11888 29832
rect 11287 29801 11299 29804
rect 11241 29795 11299 29801
rect 11882 29792 11888 29804
rect 11940 29792 11946 29844
rect 14182 29792 14188 29844
rect 14240 29832 14246 29844
rect 15013 29835 15071 29841
rect 15013 29832 15025 29835
rect 14240 29804 15025 29832
rect 14240 29792 14246 29804
rect 15013 29801 15025 29804
rect 15059 29832 15071 29835
rect 15102 29832 15108 29844
rect 15059 29804 15108 29832
rect 15059 29801 15071 29804
rect 15013 29795 15071 29801
rect 15102 29792 15108 29804
rect 15160 29792 15166 29844
rect 24857 29835 24915 29841
rect 24857 29801 24869 29835
rect 24903 29832 24915 29835
rect 26142 29832 26148 29844
rect 24903 29804 26148 29832
rect 24903 29801 24915 29804
rect 24857 29795 24915 29801
rect 26142 29792 26148 29804
rect 26200 29792 26206 29844
rect 28169 29835 28227 29841
rect 28169 29801 28181 29835
rect 28215 29832 28227 29835
rect 28810 29832 28816 29844
rect 28215 29804 28816 29832
rect 28215 29801 28227 29804
rect 28169 29795 28227 29801
rect 28810 29792 28816 29804
rect 28868 29792 28874 29844
rect 10597 29767 10655 29773
rect 10597 29733 10609 29767
rect 10643 29764 10655 29767
rect 12437 29767 12495 29773
rect 12437 29764 12449 29767
rect 10643 29736 12449 29764
rect 10643 29733 10655 29736
rect 10597 29727 10655 29733
rect 12437 29733 12449 29736
rect 12483 29764 12495 29767
rect 16850 29764 16856 29776
rect 12483 29736 16856 29764
rect 12483 29733 12495 29736
rect 12437 29727 12495 29733
rect 16850 29724 16856 29736
rect 16908 29724 16914 29776
rect 20073 29767 20131 29773
rect 20073 29764 20085 29767
rect 18432 29736 20085 29764
rect 14829 29699 14887 29705
rect 14829 29665 14841 29699
rect 14875 29696 14887 29699
rect 15286 29696 15292 29708
rect 14875 29668 15292 29696
rect 14875 29665 14887 29668
rect 14829 29659 14887 29665
rect 15286 29656 15292 29668
rect 15344 29656 15350 29708
rect 18432 29696 18460 29736
rect 20073 29733 20085 29736
rect 20119 29764 20131 29767
rect 20162 29764 20168 29776
rect 20119 29736 20168 29764
rect 20119 29733 20131 29736
rect 20073 29727 20131 29733
rect 20162 29724 20168 29736
rect 20220 29724 20226 29776
rect 15488 29668 18460 29696
rect 19705 29699 19763 29705
rect 2958 29588 2964 29640
rect 3016 29628 3022 29640
rect 5077 29631 5135 29637
rect 5077 29628 5089 29631
rect 3016 29600 5089 29628
rect 3016 29588 3022 29600
rect 5077 29597 5089 29600
rect 5123 29597 5135 29631
rect 5077 29591 5135 29597
rect 7193 29631 7251 29637
rect 7193 29597 7205 29631
rect 7239 29628 7251 29631
rect 8478 29628 8484 29640
rect 7239 29600 8484 29628
rect 7239 29597 7251 29600
rect 7193 29591 7251 29597
rect 8478 29588 8484 29600
rect 8536 29588 8542 29640
rect 10778 29588 10784 29640
rect 10836 29628 10842 29640
rect 11149 29631 11207 29637
rect 11149 29628 11161 29631
rect 10836 29600 11161 29628
rect 10836 29588 10842 29600
rect 11149 29597 11161 29600
rect 11195 29597 11207 29631
rect 11149 29591 11207 29597
rect 14645 29631 14703 29637
rect 14645 29597 14657 29631
rect 14691 29628 14703 29631
rect 15488 29628 15516 29668
rect 19705 29665 19717 29699
rect 19751 29696 19763 29699
rect 30466 29696 30472 29708
rect 19751 29668 30472 29696
rect 19751 29665 19763 29668
rect 19705 29659 19763 29665
rect 30466 29656 30472 29668
rect 30524 29656 30530 29708
rect 14691 29600 15516 29628
rect 14691 29597 14703 29600
rect 14645 29591 14703 29597
rect 15562 29588 15568 29640
rect 15620 29628 15626 29640
rect 15749 29631 15807 29637
rect 15749 29628 15761 29631
rect 15620 29600 15761 29628
rect 15620 29588 15626 29600
rect 15749 29597 15761 29600
rect 15795 29597 15807 29631
rect 15749 29591 15807 29597
rect 19334 29588 19340 29640
rect 19392 29628 19398 29640
rect 19889 29631 19947 29637
rect 19889 29628 19901 29631
rect 19392 29600 19901 29628
rect 19392 29588 19398 29600
rect 19889 29597 19901 29600
rect 19935 29597 19947 29631
rect 21082 29628 21088 29640
rect 21043 29600 21088 29628
rect 19889 29591 19947 29597
rect 21082 29588 21088 29600
rect 21140 29588 21146 29640
rect 24765 29631 24823 29637
rect 24765 29628 24777 29631
rect 22066 29600 24777 29628
rect 8662 29520 8668 29572
rect 8720 29560 8726 29572
rect 10045 29563 10103 29569
rect 10045 29560 10057 29563
rect 8720 29532 10057 29560
rect 8720 29520 8726 29532
rect 10045 29529 10057 29532
rect 10091 29529 10103 29563
rect 10045 29523 10103 29529
rect 10134 29520 10140 29572
rect 10192 29560 10198 29572
rect 11882 29560 11888 29572
rect 10192 29532 10237 29560
rect 11843 29532 11888 29560
rect 10192 29520 10198 29532
rect 11882 29520 11888 29532
rect 11940 29520 11946 29572
rect 11974 29520 11980 29572
rect 12032 29560 12038 29572
rect 18138 29560 18144 29572
rect 12032 29532 12077 29560
rect 18099 29532 18144 29560
rect 12032 29520 12038 29532
rect 18138 29520 18144 29532
rect 18196 29520 18202 29572
rect 18230 29520 18236 29572
rect 18288 29560 18294 29572
rect 18785 29563 18843 29569
rect 18288 29532 18333 29560
rect 18288 29520 18294 29532
rect 18785 29529 18797 29563
rect 18831 29560 18843 29563
rect 18874 29560 18880 29572
rect 18831 29532 18880 29560
rect 18831 29529 18843 29532
rect 18785 29523 18843 29529
rect 18874 29520 18880 29532
rect 18932 29520 18938 29572
rect 22066 29560 22094 29600
rect 24765 29597 24777 29600
rect 24811 29597 24823 29631
rect 24765 29591 24823 29597
rect 26234 29588 26240 29640
rect 26292 29628 26298 29640
rect 28077 29631 28135 29637
rect 28077 29628 28089 29631
rect 26292 29600 28089 29628
rect 26292 29588 26298 29600
rect 28077 29597 28089 29600
rect 28123 29597 28135 29631
rect 28077 29591 28135 29597
rect 18984 29532 22094 29560
rect 15838 29492 15844 29504
rect 15799 29464 15844 29492
rect 15838 29452 15844 29464
rect 15896 29452 15902 29504
rect 16574 29452 16580 29504
rect 16632 29492 16638 29504
rect 18984 29492 19012 29532
rect 16632 29464 19012 29492
rect 16632 29452 16638 29464
rect 20990 29452 20996 29504
rect 21048 29492 21054 29504
rect 21269 29495 21327 29501
rect 21269 29492 21281 29495
rect 21048 29464 21281 29492
rect 21048 29452 21054 29464
rect 21269 29461 21281 29464
rect 21315 29461 21327 29495
rect 21269 29455 21327 29461
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 8662 29288 8668 29300
rect 8623 29260 8668 29288
rect 8662 29248 8668 29260
rect 8720 29248 8726 29300
rect 10045 29291 10103 29297
rect 10045 29257 10057 29291
rect 10091 29288 10103 29291
rect 10134 29288 10140 29300
rect 10091 29260 10140 29288
rect 10091 29257 10103 29260
rect 10045 29251 10103 29257
rect 10134 29248 10140 29260
rect 10192 29248 10198 29300
rect 11882 29288 11888 29300
rect 11843 29260 11888 29288
rect 11882 29248 11888 29260
rect 11940 29248 11946 29300
rect 15102 29288 15108 29300
rect 15063 29260 15108 29288
rect 15102 29248 15108 29260
rect 15160 29248 15166 29300
rect 18138 29288 18144 29300
rect 18099 29260 18144 29288
rect 18138 29248 18144 29260
rect 18196 29248 18202 29300
rect 19334 29288 19340 29300
rect 19295 29260 19340 29288
rect 19334 29248 19340 29260
rect 19392 29248 19398 29300
rect 19978 29288 19984 29300
rect 19939 29260 19984 29288
rect 19978 29248 19984 29260
rect 20036 29248 20042 29300
rect 20809 29291 20867 29297
rect 20809 29257 20821 29291
rect 20855 29288 20867 29291
rect 22002 29288 22008 29300
rect 20855 29260 22008 29288
rect 20855 29257 20867 29260
rect 20809 29251 20867 29257
rect 22002 29248 22008 29260
rect 22060 29248 22066 29300
rect 24026 29220 24032 29232
rect 14476 29192 24032 29220
rect 1762 29152 1768 29164
rect 1723 29124 1768 29152
rect 1762 29112 1768 29124
rect 1820 29112 1826 29164
rect 9953 29155 10011 29161
rect 9953 29121 9965 29155
rect 9999 29152 10011 29155
rect 11238 29152 11244 29164
rect 9999 29124 11244 29152
rect 9999 29121 10011 29124
rect 9953 29115 10011 29121
rect 11238 29112 11244 29124
rect 11296 29112 11302 29164
rect 14476 29161 14504 29192
rect 24026 29180 24032 29192
rect 24084 29180 24090 29232
rect 14461 29155 14519 29161
rect 14461 29121 14473 29155
rect 14507 29121 14519 29155
rect 14461 29115 14519 29121
rect 14645 29155 14703 29161
rect 14645 29121 14657 29155
rect 14691 29152 14703 29155
rect 15838 29152 15844 29164
rect 14691 29124 15844 29152
rect 14691 29121 14703 29124
rect 14645 29115 14703 29121
rect 15838 29112 15844 29124
rect 15896 29112 15902 29164
rect 19242 29152 19248 29164
rect 19203 29124 19248 29152
rect 19242 29112 19248 29124
rect 19300 29112 19306 29164
rect 19889 29155 19947 29161
rect 19889 29121 19901 29155
rect 19935 29152 19947 29155
rect 20162 29152 20168 29164
rect 19935 29124 20168 29152
rect 19935 29121 19947 29124
rect 19889 29115 19947 29121
rect 20162 29112 20168 29124
rect 20220 29112 20226 29164
rect 20990 29152 20996 29164
rect 20951 29124 20996 29152
rect 20990 29112 20996 29124
rect 21048 29112 21054 29164
rect 38286 29152 38292 29164
rect 38247 29124 38292 29152
rect 38286 29112 38292 29124
rect 38344 29112 38350 29164
rect 8018 29084 8024 29096
rect 7979 29056 8024 29084
rect 8018 29044 8024 29056
rect 8076 29044 8082 29096
rect 8202 29084 8208 29096
rect 8163 29056 8208 29084
rect 8202 29044 8208 29056
rect 8260 29044 8266 29096
rect 1581 29019 1639 29025
rect 1581 28985 1593 29019
rect 1627 29016 1639 29019
rect 5718 29016 5724 29028
rect 1627 28988 5724 29016
rect 1627 28985 1639 28988
rect 1581 28979 1639 28985
rect 5718 28976 5724 28988
rect 5776 28976 5782 29028
rect 34514 28976 34520 29028
rect 34572 29016 34578 29028
rect 38105 29019 38163 29025
rect 38105 29016 38117 29019
rect 34572 28988 38117 29016
rect 34572 28976 34578 28988
rect 38105 28985 38117 28988
rect 38151 28985 38163 29019
rect 38105 28979 38163 28985
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 12434 28704 12440 28756
rect 12492 28744 12498 28756
rect 13081 28747 13139 28753
rect 13081 28744 13093 28747
rect 12492 28716 13093 28744
rect 12492 28704 12498 28716
rect 13081 28713 13093 28716
rect 13127 28744 13139 28747
rect 13262 28744 13268 28756
rect 13127 28716 13268 28744
rect 13127 28713 13139 28716
rect 13081 28707 13139 28713
rect 13262 28704 13268 28716
rect 13320 28704 13326 28756
rect 13446 28704 13452 28756
rect 13504 28744 13510 28756
rect 22094 28744 22100 28756
rect 13504 28716 22100 28744
rect 13504 28704 13510 28716
rect 22094 28704 22100 28716
rect 22152 28704 22158 28756
rect 28997 28747 29055 28753
rect 28997 28713 29009 28747
rect 29043 28744 29055 28747
rect 33594 28744 33600 28756
rect 29043 28716 33600 28744
rect 29043 28713 29055 28716
rect 28997 28707 29055 28713
rect 33594 28704 33600 28716
rect 33652 28704 33658 28756
rect 7745 28679 7803 28685
rect 7745 28645 7757 28679
rect 7791 28676 7803 28679
rect 8018 28676 8024 28688
rect 7791 28648 8024 28676
rect 7791 28645 7803 28648
rect 7745 28639 7803 28645
rect 8018 28636 8024 28648
rect 8076 28676 8082 28688
rect 14734 28676 14740 28688
rect 8076 28648 14740 28676
rect 8076 28636 8082 28648
rect 14734 28636 14740 28648
rect 14792 28636 14798 28688
rect 13998 28568 14004 28620
rect 14056 28608 14062 28620
rect 14056 28580 16068 28608
rect 14056 28568 14062 28580
rect 7650 28540 7656 28552
rect 7611 28512 7656 28540
rect 7650 28500 7656 28512
rect 7708 28500 7714 28552
rect 8478 28540 8484 28552
rect 8439 28512 8484 28540
rect 8478 28500 8484 28512
rect 8536 28500 8542 28552
rect 10226 28540 10232 28552
rect 10187 28512 10232 28540
rect 10226 28500 10232 28512
rect 10284 28500 10290 28552
rect 10686 28540 10692 28552
rect 10647 28512 10692 28540
rect 10686 28500 10692 28512
rect 10744 28500 10750 28552
rect 12713 28543 12771 28549
rect 12713 28509 12725 28543
rect 12759 28509 12771 28543
rect 12894 28540 12900 28552
rect 12855 28512 12900 28540
rect 12713 28503 12771 28509
rect 12728 28472 12756 28503
rect 12894 28500 12900 28512
rect 12952 28500 12958 28552
rect 16040 28549 16068 28580
rect 15381 28543 15439 28549
rect 15381 28509 15393 28543
rect 15427 28540 15439 28543
rect 16025 28543 16083 28549
rect 15427 28512 15884 28540
rect 15427 28509 15439 28512
rect 15381 28503 15439 28509
rect 15286 28472 15292 28484
rect 12728 28444 15292 28472
rect 15286 28432 15292 28444
rect 15344 28432 15350 28484
rect 8297 28407 8355 28413
rect 8297 28373 8309 28407
rect 8343 28404 8355 28407
rect 8386 28404 8392 28416
rect 8343 28376 8392 28404
rect 8343 28373 8355 28376
rect 8297 28367 8355 28373
rect 8386 28364 8392 28376
rect 8444 28364 8450 28416
rect 10042 28404 10048 28416
rect 10003 28376 10048 28404
rect 10042 28364 10048 28376
rect 10100 28364 10106 28416
rect 10781 28407 10839 28413
rect 10781 28373 10793 28407
rect 10827 28404 10839 28407
rect 11698 28404 11704 28416
rect 10827 28376 11704 28404
rect 10827 28373 10839 28376
rect 10781 28367 10839 28373
rect 11698 28364 11704 28376
rect 11756 28364 11762 28416
rect 14458 28364 14464 28416
rect 14516 28404 14522 28416
rect 14553 28407 14611 28413
rect 14553 28404 14565 28407
rect 14516 28376 14565 28404
rect 14516 28364 14522 28376
rect 14553 28373 14565 28376
rect 14599 28373 14611 28407
rect 15194 28404 15200 28416
rect 15155 28376 15200 28404
rect 14553 28367 14611 28373
rect 15194 28364 15200 28376
rect 15252 28364 15258 28416
rect 15856 28413 15884 28512
rect 16025 28509 16037 28543
rect 16071 28509 16083 28543
rect 16025 28503 16083 28509
rect 26418 28500 26424 28552
rect 26476 28540 26482 28552
rect 28905 28543 28963 28549
rect 28905 28540 28917 28543
rect 26476 28512 28917 28540
rect 26476 28500 26482 28512
rect 28905 28509 28917 28512
rect 28951 28509 28963 28543
rect 28905 28503 28963 28509
rect 31021 28543 31079 28549
rect 31021 28509 31033 28543
rect 31067 28540 31079 28543
rect 34514 28540 34520 28552
rect 31067 28512 34520 28540
rect 31067 28509 31079 28512
rect 31021 28503 31079 28509
rect 34514 28500 34520 28512
rect 34572 28500 34578 28552
rect 15841 28407 15899 28413
rect 15841 28373 15853 28407
rect 15887 28373 15899 28407
rect 15841 28367 15899 28373
rect 19889 28407 19947 28413
rect 19889 28373 19901 28407
rect 19935 28404 19947 28407
rect 19978 28404 19984 28416
rect 19935 28376 19984 28404
rect 19935 28373 19947 28376
rect 19889 28367 19947 28373
rect 19978 28364 19984 28376
rect 20036 28364 20042 28416
rect 29454 28364 29460 28416
rect 29512 28404 29518 28416
rect 31113 28407 31171 28413
rect 31113 28404 31125 28407
rect 29512 28376 31125 28404
rect 29512 28364 29518 28376
rect 31113 28373 31125 28376
rect 31159 28373 31171 28407
rect 31113 28367 31171 28373
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 8202 28200 8208 28212
rect 8163 28172 8208 28200
rect 8202 28160 8208 28172
rect 8260 28160 8266 28212
rect 12069 28203 12127 28209
rect 12069 28169 12081 28203
rect 12115 28200 12127 28203
rect 12894 28200 12900 28212
rect 12115 28172 12900 28200
rect 12115 28169 12127 28172
rect 12069 28163 12127 28169
rect 12894 28160 12900 28172
rect 12952 28160 12958 28212
rect 13262 28200 13268 28212
rect 13223 28172 13268 28200
rect 13262 28160 13268 28172
rect 13320 28160 13326 28212
rect 19978 28200 19984 28212
rect 19628 28172 19984 28200
rect 14458 28132 14464 28144
rect 14419 28104 14464 28132
rect 14458 28092 14464 28104
rect 14516 28092 14522 28144
rect 14553 28135 14611 28141
rect 14553 28101 14565 28135
rect 14599 28132 14611 28135
rect 16114 28132 16120 28144
rect 14599 28104 16120 28132
rect 14599 28101 14611 28104
rect 14553 28095 14611 28101
rect 16114 28092 16120 28104
rect 16172 28092 16178 28144
rect 19628 28141 19656 28172
rect 19978 28160 19984 28172
rect 20036 28160 20042 28212
rect 23477 28203 23535 28209
rect 23477 28169 23489 28203
rect 23523 28169 23535 28203
rect 28534 28200 28540 28212
rect 28495 28172 28540 28200
rect 23477 28163 23535 28169
rect 19613 28135 19671 28141
rect 19613 28101 19625 28135
rect 19659 28101 19671 28135
rect 19613 28095 19671 28101
rect 19705 28135 19763 28141
rect 19705 28101 19717 28135
rect 19751 28132 19763 28135
rect 20070 28132 20076 28144
rect 19751 28104 20076 28132
rect 19751 28101 19763 28104
rect 19705 28095 19763 28101
rect 20070 28092 20076 28104
rect 20128 28092 20134 28144
rect 20898 28132 20904 28144
rect 20859 28104 20904 28132
rect 20898 28092 20904 28104
rect 20956 28092 20962 28144
rect 21910 28092 21916 28144
rect 21968 28132 21974 28144
rect 23492 28132 23520 28163
rect 28534 28160 28540 28172
rect 28592 28160 28598 28212
rect 35434 28200 35440 28212
rect 35395 28172 35440 28200
rect 35434 28160 35440 28172
rect 35492 28160 35498 28212
rect 21968 28104 23428 28132
rect 23492 28104 24348 28132
rect 21968 28092 21974 28104
rect 3970 28024 3976 28076
rect 4028 28064 4034 28076
rect 6917 28067 6975 28073
rect 6917 28064 6929 28067
rect 4028 28036 6929 28064
rect 4028 28024 4034 28036
rect 6917 28033 6929 28036
rect 6963 28033 6975 28067
rect 8386 28064 8392 28076
rect 8347 28036 8392 28064
rect 6917 28027 6975 28033
rect 8386 28024 8392 28036
rect 8444 28024 8450 28076
rect 8938 28064 8944 28076
rect 8899 28036 8944 28064
rect 8938 28024 8944 28036
rect 8996 28024 9002 28076
rect 10042 28064 10048 28076
rect 10003 28036 10048 28064
rect 10042 28024 10048 28036
rect 10100 28024 10106 28076
rect 11977 28067 12035 28073
rect 11977 28033 11989 28067
rect 12023 28064 12035 28067
rect 13998 28064 14004 28076
rect 12023 28036 14004 28064
rect 12023 28033 12035 28036
rect 11977 28027 12035 28033
rect 13998 28024 14004 28036
rect 14056 28024 14062 28076
rect 22005 28067 22063 28073
rect 22005 28033 22017 28067
rect 22051 28064 22063 28067
rect 22738 28064 22744 28076
rect 22051 28036 22744 28064
rect 22051 28033 22063 28036
rect 22005 28027 22063 28033
rect 22738 28024 22744 28036
rect 22796 28024 22802 28076
rect 23400 28064 23428 28104
rect 24320 28073 24348 28104
rect 27798 28092 27804 28144
rect 27856 28132 27862 28144
rect 27856 28104 28488 28132
rect 27856 28092 27862 28104
rect 23661 28067 23719 28073
rect 23661 28064 23673 28067
rect 23400 28036 23673 28064
rect 23661 28033 23673 28036
rect 23707 28033 23719 28067
rect 23661 28027 23719 28033
rect 24305 28067 24363 28073
rect 24305 28033 24317 28067
rect 24351 28033 24363 28067
rect 24305 28027 24363 28033
rect 27341 28067 27399 28073
rect 27341 28033 27353 28067
rect 27387 28033 27399 28067
rect 27982 28064 27988 28076
rect 27943 28036 27988 28064
rect 27341 28027 27399 28033
rect 9033 27999 9091 28005
rect 9033 27965 9045 27999
rect 9079 27996 9091 27999
rect 9858 27996 9864 28008
rect 9079 27968 9864 27996
rect 9079 27965 9091 27968
rect 9033 27959 9091 27965
rect 9858 27956 9864 27968
rect 9916 27956 9922 28008
rect 12618 27996 12624 28008
rect 12579 27968 12624 27996
rect 12618 27956 12624 27968
rect 12676 27956 12682 28008
rect 12805 27999 12863 28005
rect 12805 27965 12817 27999
rect 12851 27996 12863 27999
rect 15194 27996 15200 28008
rect 12851 27968 15200 27996
rect 12851 27965 12863 27968
rect 12805 27959 12863 27965
rect 15194 27956 15200 27968
rect 15252 27956 15258 28008
rect 15286 27956 15292 28008
rect 15344 27996 15350 28008
rect 20809 27999 20867 28005
rect 15344 27968 20300 27996
rect 15344 27956 15350 27968
rect 15013 27931 15071 27937
rect 15013 27897 15025 27931
rect 15059 27928 15071 27931
rect 15102 27928 15108 27940
rect 15059 27900 15108 27928
rect 15059 27897 15071 27900
rect 15013 27891 15071 27897
rect 15102 27888 15108 27900
rect 15160 27888 15166 27940
rect 20162 27928 20168 27940
rect 20123 27900 20168 27928
rect 20162 27888 20168 27900
rect 20220 27888 20226 27940
rect 20272 27928 20300 27968
rect 20809 27965 20821 27999
rect 20855 27996 20867 27999
rect 23198 27996 23204 28008
rect 20855 27968 23204 27996
rect 20855 27965 20867 27968
rect 20809 27959 20867 27965
rect 23198 27956 23204 27968
rect 23256 27956 23262 28008
rect 24857 27999 24915 28005
rect 24857 27996 24869 27999
rect 23308 27968 24869 27996
rect 20622 27928 20628 27940
rect 20272 27900 20628 27928
rect 20622 27888 20628 27900
rect 20680 27928 20686 27940
rect 21361 27931 21419 27937
rect 21361 27928 21373 27931
rect 20680 27900 21373 27928
rect 20680 27888 20686 27900
rect 21361 27897 21373 27900
rect 21407 27897 21419 27931
rect 21361 27891 21419 27897
rect 22094 27888 22100 27940
rect 22152 27928 22158 27940
rect 23308 27928 23336 27968
rect 24857 27965 24869 27968
rect 24903 27965 24915 27999
rect 24857 27959 24915 27965
rect 25041 27999 25099 28005
rect 25041 27965 25053 27999
rect 25087 27965 25099 27999
rect 25041 27959 25099 27965
rect 22152 27900 23336 27928
rect 24121 27931 24179 27937
rect 22152 27888 22158 27900
rect 24121 27897 24133 27931
rect 24167 27928 24179 27931
rect 25056 27928 25084 27959
rect 24167 27900 25084 27928
rect 25501 27931 25559 27937
rect 24167 27897 24179 27900
rect 24121 27891 24179 27897
rect 25501 27897 25513 27931
rect 25547 27928 25559 27931
rect 27356 27928 27384 28027
rect 27982 28024 27988 28036
rect 28040 28024 28046 28076
rect 28460 28073 28488 28104
rect 28445 28067 28503 28073
rect 28445 28033 28457 28067
rect 28491 28033 28503 28067
rect 29454 28064 29460 28076
rect 29415 28036 29460 28064
rect 28445 28027 28503 28033
rect 29454 28024 29460 28036
rect 29512 28024 29518 28076
rect 33134 28024 33140 28076
rect 33192 28064 33198 28076
rect 35621 28067 35679 28073
rect 35621 28064 35633 28067
rect 33192 28036 35633 28064
rect 33192 28024 33198 28036
rect 35621 28033 35633 28036
rect 35667 28033 35679 28067
rect 35621 28027 35679 28033
rect 29638 27996 29644 28008
rect 29599 27968 29644 27996
rect 29638 27956 29644 27968
rect 29696 27956 29702 28008
rect 27801 27931 27859 27937
rect 27801 27928 27813 27931
rect 25547 27900 27292 27928
rect 27356 27900 27813 27928
rect 25547 27897 25559 27900
rect 25501 27891 25559 27897
rect 27264 27872 27292 27900
rect 27801 27897 27813 27900
rect 27847 27897 27859 27931
rect 27801 27891 27859 27897
rect 6822 27820 6828 27872
rect 6880 27860 6886 27872
rect 7009 27863 7067 27869
rect 7009 27860 7021 27863
rect 6880 27832 7021 27860
rect 6880 27820 6886 27832
rect 7009 27829 7021 27832
rect 7055 27829 7067 27863
rect 10502 27860 10508 27872
rect 10463 27832 10508 27860
rect 7009 27823 7067 27829
rect 10502 27820 10508 27832
rect 10560 27820 10566 27872
rect 27154 27860 27160 27872
rect 27115 27832 27160 27860
rect 27154 27820 27160 27832
rect 27212 27820 27218 27872
rect 27246 27820 27252 27872
rect 27304 27860 27310 27872
rect 29825 27863 29883 27869
rect 29825 27860 29837 27863
rect 27304 27832 29837 27860
rect 27304 27820 27310 27832
rect 29825 27829 29837 27832
rect 29871 27829 29883 27863
rect 29825 27823 29883 27829
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 5902 27616 5908 27668
rect 5960 27656 5966 27668
rect 6822 27656 6828 27668
rect 5960 27628 6828 27656
rect 5960 27616 5966 27628
rect 6822 27616 6828 27628
rect 6880 27656 6886 27668
rect 6880 27616 6914 27656
rect 9858 27616 9864 27668
rect 9916 27656 9922 27668
rect 19426 27656 19432 27668
rect 9916 27628 19432 27656
rect 9916 27616 9922 27628
rect 19426 27616 19432 27628
rect 19484 27616 19490 27668
rect 29638 27616 29644 27668
rect 29696 27656 29702 27668
rect 29825 27659 29883 27665
rect 29825 27656 29837 27659
rect 29696 27628 29837 27656
rect 29696 27616 29702 27628
rect 29825 27625 29837 27628
rect 29871 27625 29883 27659
rect 29825 27619 29883 27625
rect 6549 27591 6607 27597
rect 6549 27557 6561 27591
rect 6595 27557 6607 27591
rect 6886 27588 6914 27616
rect 10502 27588 10508 27600
rect 6886 27560 9260 27588
rect 6549 27551 6607 27557
rect 6564 27520 6592 27551
rect 6564 27492 8064 27520
rect 1762 27452 1768 27464
rect 1723 27424 1768 27452
rect 1762 27412 1768 27424
rect 1820 27412 1826 27464
rect 5718 27452 5724 27464
rect 5679 27424 5724 27452
rect 5718 27412 5724 27424
rect 5776 27412 5782 27464
rect 6730 27452 6736 27464
rect 6691 27424 6736 27452
rect 6730 27412 6736 27424
rect 6788 27412 6794 27464
rect 7190 27452 7196 27464
rect 7151 27424 7196 27452
rect 7190 27412 7196 27424
rect 7248 27412 7254 27464
rect 8036 27461 8064 27492
rect 8021 27455 8079 27461
rect 8021 27421 8033 27455
rect 8067 27421 8079 27455
rect 8021 27415 8079 27421
rect 7285 27387 7343 27393
rect 7285 27353 7297 27387
rect 7331 27384 7343 27387
rect 8938 27384 8944 27396
rect 7331 27356 8944 27384
rect 7331 27353 7343 27356
rect 7285 27347 7343 27353
rect 8938 27344 8944 27356
rect 8996 27344 9002 27396
rect 1581 27319 1639 27325
rect 1581 27285 1593 27319
rect 1627 27316 1639 27319
rect 5350 27316 5356 27328
rect 1627 27288 5356 27316
rect 1627 27285 1639 27288
rect 1581 27279 1639 27285
rect 5350 27276 5356 27288
rect 5408 27276 5414 27328
rect 5810 27316 5816 27328
rect 5771 27288 5816 27316
rect 5810 27276 5816 27288
rect 5868 27276 5874 27328
rect 7834 27316 7840 27328
rect 7795 27288 7840 27316
rect 7834 27276 7840 27288
rect 7892 27276 7898 27328
rect 9122 27316 9128 27328
rect 9083 27288 9128 27316
rect 9122 27276 9128 27288
rect 9180 27276 9186 27328
rect 9232 27316 9260 27560
rect 10152 27560 10508 27588
rect 10152 27529 10180 27560
rect 10502 27548 10508 27560
rect 10560 27588 10566 27600
rect 11609 27591 11667 27597
rect 11609 27588 11621 27591
rect 10560 27560 11621 27588
rect 10560 27548 10566 27560
rect 11609 27557 11621 27560
rect 11655 27557 11667 27591
rect 11609 27551 11667 27557
rect 26786 27548 26792 27600
rect 26844 27588 26850 27600
rect 32953 27591 33011 27597
rect 26844 27560 32904 27588
rect 26844 27548 26850 27560
rect 10137 27523 10195 27529
rect 10137 27489 10149 27523
rect 10183 27489 10195 27523
rect 11514 27520 11520 27532
rect 10137 27483 10195 27489
rect 10244 27492 11520 27520
rect 9309 27455 9367 27461
rect 9309 27421 9321 27455
rect 9355 27452 9367 27455
rect 10244 27452 10272 27492
rect 11514 27480 11520 27492
rect 11572 27480 11578 27532
rect 12618 27480 12624 27532
rect 12676 27520 12682 27532
rect 12713 27523 12771 27529
rect 12713 27520 12725 27523
rect 12676 27492 12725 27520
rect 12676 27480 12682 27492
rect 12713 27489 12725 27492
rect 12759 27489 12771 27523
rect 12713 27483 12771 27489
rect 26421 27523 26479 27529
rect 26421 27489 26433 27523
rect 26467 27520 26479 27523
rect 27246 27520 27252 27532
rect 26467 27492 27252 27520
rect 26467 27489 26479 27492
rect 26421 27483 26479 27489
rect 27246 27480 27252 27492
rect 27304 27480 27310 27532
rect 27982 27480 27988 27532
rect 28040 27520 28046 27532
rect 32876 27520 32904 27560
rect 32953 27557 32965 27591
rect 32999 27588 33011 27591
rect 33134 27588 33140 27600
rect 32999 27560 33140 27588
rect 32999 27557 33011 27560
rect 32953 27551 33011 27557
rect 33134 27548 33140 27560
rect 33192 27548 33198 27600
rect 28040 27492 29776 27520
rect 32876 27492 35894 27520
rect 28040 27480 28046 27492
rect 9355 27424 10272 27452
rect 9355 27421 9367 27424
rect 9309 27415 9367 27421
rect 10318 27412 10324 27464
rect 10376 27452 10382 27464
rect 10778 27452 10784 27464
rect 10376 27424 10421 27452
rect 10739 27424 10784 27452
rect 10376 27412 10382 27424
rect 10778 27412 10784 27424
rect 10836 27412 10842 27464
rect 11241 27455 11299 27461
rect 11241 27421 11253 27455
rect 11287 27421 11299 27455
rect 11422 27452 11428 27464
rect 11383 27424 11428 27452
rect 11241 27415 11299 27421
rect 11256 27316 11284 27415
rect 11422 27412 11428 27424
rect 11480 27412 11486 27464
rect 16758 27452 16764 27464
rect 16719 27424 16764 27452
rect 16758 27412 16764 27424
rect 16816 27412 16822 27464
rect 26602 27452 26608 27464
rect 26563 27424 26608 27452
rect 26602 27412 26608 27424
rect 26660 27412 26666 27464
rect 28813 27455 28871 27461
rect 28813 27421 28825 27455
rect 28859 27452 28871 27455
rect 28902 27452 28908 27464
rect 28859 27424 28908 27452
rect 28859 27421 28871 27424
rect 28813 27415 28871 27421
rect 28902 27412 28908 27424
rect 28960 27412 28966 27464
rect 29748 27461 29776 27492
rect 29733 27455 29791 27461
rect 29733 27421 29745 27455
rect 29779 27421 29791 27455
rect 29733 27415 29791 27421
rect 32861 27455 32919 27461
rect 32861 27421 32873 27455
rect 32907 27421 32919 27455
rect 35866 27452 35894 27492
rect 38013 27455 38071 27461
rect 38013 27452 38025 27455
rect 35866 27424 38025 27452
rect 32861 27415 32919 27421
rect 38013 27421 38025 27424
rect 38059 27421 38071 27455
rect 38013 27415 38071 27421
rect 17494 27384 17500 27396
rect 17455 27356 17500 27384
rect 17494 27344 17500 27356
rect 17552 27344 17558 27396
rect 17589 27387 17647 27393
rect 17589 27353 17601 27387
rect 17635 27353 17647 27387
rect 18138 27384 18144 27396
rect 18099 27356 18144 27384
rect 17589 27347 17647 27353
rect 13262 27316 13268 27328
rect 9232 27288 13268 27316
rect 13262 27276 13268 27288
rect 13320 27276 13326 27328
rect 16853 27319 16911 27325
rect 16853 27285 16865 27319
rect 16899 27316 16911 27319
rect 17604 27316 17632 27347
rect 18138 27344 18144 27356
rect 18196 27344 18202 27396
rect 23842 27344 23848 27396
rect 23900 27384 23906 27396
rect 32876 27384 32904 27415
rect 23900 27356 32904 27384
rect 23900 27344 23906 27356
rect 16899 27288 17632 27316
rect 27065 27319 27123 27325
rect 16899 27285 16911 27288
rect 16853 27279 16911 27285
rect 27065 27285 27077 27319
rect 27111 27316 27123 27319
rect 27798 27316 27804 27328
rect 27111 27288 27804 27316
rect 27111 27285 27123 27288
rect 27065 27279 27123 27285
rect 27798 27276 27804 27288
rect 27856 27276 27862 27328
rect 28258 27276 28264 27328
rect 28316 27316 28322 27328
rect 28905 27319 28963 27325
rect 28905 27316 28917 27319
rect 28316 27288 28917 27316
rect 28316 27276 28322 27288
rect 28905 27285 28917 27288
rect 28951 27285 28963 27319
rect 38194 27316 38200 27328
rect 38155 27288 38200 27316
rect 28905 27279 28963 27285
rect 38194 27276 38200 27288
rect 38252 27276 38258 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 10229 27115 10287 27121
rect 10229 27081 10241 27115
rect 10275 27112 10287 27115
rect 11422 27112 11428 27124
rect 10275 27084 11428 27112
rect 10275 27081 10287 27084
rect 10229 27075 10287 27081
rect 11422 27072 11428 27084
rect 11480 27072 11486 27124
rect 11793 27115 11851 27121
rect 11793 27081 11805 27115
rect 11839 27081 11851 27115
rect 11793 27075 11851 27081
rect 6730 27004 6736 27056
rect 6788 27044 6794 27056
rect 6788 27016 10180 27044
rect 6788 27004 6794 27016
rect 5810 26936 5816 26988
rect 5868 26976 5874 26988
rect 7101 26979 7159 26985
rect 7101 26976 7113 26979
rect 5868 26948 7113 26976
rect 5868 26936 5874 26948
rect 7101 26945 7113 26948
rect 7147 26945 7159 26979
rect 9122 26976 9128 26988
rect 9083 26948 9128 26976
rect 7101 26939 7159 26945
rect 9122 26936 9128 26948
rect 9180 26936 9186 26988
rect 10152 26985 10180 27016
rect 10318 27004 10324 27056
rect 10376 27044 10382 27056
rect 11808 27044 11836 27075
rect 17494 27072 17500 27124
rect 17552 27112 17558 27124
rect 18141 27115 18199 27121
rect 18141 27112 18153 27115
rect 17552 27084 18153 27112
rect 17552 27072 17558 27084
rect 18141 27081 18153 27084
rect 18187 27081 18199 27115
rect 18141 27075 18199 27081
rect 18230 27072 18236 27124
rect 18288 27112 18294 27124
rect 19153 27115 19211 27121
rect 19153 27112 19165 27115
rect 18288 27084 19165 27112
rect 18288 27072 18294 27084
rect 19153 27081 19165 27084
rect 19199 27081 19211 27115
rect 19153 27075 19211 27081
rect 22005 27115 22063 27121
rect 22005 27081 22017 27115
rect 22051 27081 22063 27115
rect 22005 27075 22063 27081
rect 23293 27115 23351 27121
rect 23293 27081 23305 27115
rect 23339 27081 23351 27115
rect 23293 27075 23351 27081
rect 25869 27115 25927 27121
rect 25869 27081 25881 27115
rect 25915 27112 25927 27115
rect 26602 27112 26608 27124
rect 25915 27084 26608 27112
rect 25915 27081 25927 27084
rect 25869 27075 25927 27081
rect 13262 27044 13268 27056
rect 10376 27016 11836 27044
rect 13223 27016 13268 27044
rect 10376 27004 10382 27016
rect 13262 27004 13268 27016
rect 13320 27004 13326 27056
rect 13357 27047 13415 27053
rect 13357 27013 13369 27047
rect 13403 27044 13415 27047
rect 13538 27044 13544 27056
rect 13403 27016 13544 27044
rect 13403 27013 13415 27016
rect 13357 27007 13415 27013
rect 13538 27004 13544 27016
rect 13596 27004 13602 27056
rect 16758 27004 16764 27056
rect 16816 27044 16822 27056
rect 22020 27044 22048 27075
rect 23308 27044 23336 27075
rect 26602 27072 26608 27084
rect 26660 27072 26666 27124
rect 16816 27016 21312 27044
rect 22020 27016 22876 27044
rect 23308 27016 24164 27044
rect 16816 27004 16822 27016
rect 10137 26979 10195 26985
rect 10137 26945 10149 26979
rect 10183 26976 10195 26979
rect 10965 26979 11023 26985
rect 10965 26976 10977 26979
rect 10183 26948 10977 26976
rect 10183 26945 10195 26948
rect 10137 26939 10195 26945
rect 10965 26945 10977 26948
rect 11011 26945 11023 26979
rect 10965 26939 11023 26945
rect 11514 26936 11520 26988
rect 11572 26976 11578 26988
rect 11701 26979 11759 26985
rect 11701 26976 11713 26979
rect 11572 26948 11713 26976
rect 11572 26936 11578 26948
rect 11701 26945 11713 26948
rect 11747 26945 11759 26979
rect 14734 26976 14740 26988
rect 14695 26948 14740 26976
rect 11701 26939 11759 26945
rect 14734 26936 14740 26948
rect 14792 26936 14798 26988
rect 17405 26979 17463 26985
rect 17405 26945 17417 26979
rect 17451 26976 17463 26979
rect 17586 26976 17592 26988
rect 17451 26948 17592 26976
rect 17451 26945 17463 26948
rect 17405 26939 17463 26945
rect 17586 26936 17592 26948
rect 17644 26936 17650 26988
rect 17954 26976 17960 26988
rect 17915 26948 17960 26976
rect 17954 26936 17960 26948
rect 18012 26936 18018 26988
rect 19334 26976 19340 26988
rect 19295 26948 19340 26976
rect 19334 26936 19340 26948
rect 19392 26936 19398 26988
rect 21174 26976 21180 26988
rect 21135 26948 21180 26976
rect 21174 26936 21180 26948
rect 21232 26936 21238 26988
rect 21284 26976 21312 27016
rect 22848 26985 22876 27016
rect 24136 26985 24164 27016
rect 22189 26979 22247 26985
rect 22189 26976 22201 26979
rect 21284 26948 22201 26976
rect 22189 26945 22201 26948
rect 22235 26945 22247 26979
rect 22189 26939 22247 26945
rect 22833 26979 22891 26985
rect 22833 26945 22845 26979
rect 22879 26945 22891 26979
rect 22833 26939 22891 26945
rect 23477 26979 23535 26985
rect 23477 26945 23489 26979
rect 23523 26945 23535 26979
rect 23477 26939 23535 26945
rect 24121 26979 24179 26985
rect 24121 26945 24133 26979
rect 24167 26945 24179 26979
rect 25130 26976 25136 26988
rect 25091 26948 25136 26976
rect 24121 26939 24179 26945
rect 7285 26911 7343 26917
rect 7285 26877 7297 26911
rect 7331 26908 7343 26911
rect 8294 26908 8300 26920
rect 7331 26880 8300 26908
rect 7331 26877 7343 26880
rect 7285 26871 7343 26877
rect 8294 26868 8300 26880
rect 8352 26868 8358 26920
rect 14918 26908 14924 26920
rect 14879 26880 14924 26908
rect 14918 26868 14924 26880
rect 14976 26868 14982 26920
rect 16117 26911 16175 26917
rect 16117 26877 16129 26911
rect 16163 26908 16175 26911
rect 16482 26908 16488 26920
rect 16163 26880 16488 26908
rect 16163 26877 16175 26880
rect 16117 26871 16175 26877
rect 16482 26868 16488 26880
rect 16540 26868 16546 26920
rect 18690 26868 18696 26920
rect 18748 26908 18754 26920
rect 23492 26908 23520 26939
rect 25130 26936 25136 26948
rect 25188 26936 25194 26988
rect 25314 26936 25320 26988
rect 25372 26976 25378 26988
rect 25777 26979 25835 26985
rect 25777 26976 25789 26979
rect 25372 26948 25789 26976
rect 25372 26936 25378 26948
rect 25777 26945 25789 26948
rect 25823 26945 25835 26979
rect 32398 26976 32404 26988
rect 32359 26948 32404 26976
rect 25777 26939 25835 26945
rect 32398 26936 32404 26948
rect 32456 26936 32462 26988
rect 18748 26880 23520 26908
rect 18748 26868 18754 26880
rect 25958 26868 25964 26920
rect 26016 26908 26022 26920
rect 26421 26911 26479 26917
rect 26421 26908 26433 26911
rect 26016 26880 26433 26908
rect 26016 26868 26022 26880
rect 26421 26877 26433 26880
rect 26467 26877 26479 26911
rect 26421 26871 26479 26877
rect 10226 26800 10232 26852
rect 10284 26840 10290 26852
rect 10781 26843 10839 26849
rect 10781 26840 10793 26843
rect 10284 26812 10793 26840
rect 10284 26800 10290 26812
rect 10781 26809 10793 26812
rect 10827 26809 10839 26843
rect 10781 26803 10839 26809
rect 13817 26843 13875 26849
rect 13817 26809 13829 26843
rect 13863 26840 13875 26843
rect 20806 26840 20812 26852
rect 13863 26812 20812 26840
rect 13863 26809 13875 26812
rect 13817 26803 13875 26809
rect 20806 26800 20812 26812
rect 20864 26800 20870 26852
rect 22649 26843 22707 26849
rect 22649 26809 22661 26843
rect 22695 26840 22707 26843
rect 24302 26840 24308 26852
rect 22695 26812 24308 26840
rect 22695 26809 22707 26812
rect 22649 26803 22707 26809
rect 24302 26800 24308 26812
rect 24360 26800 24366 26852
rect 7742 26772 7748 26784
rect 7703 26744 7748 26772
rect 7742 26732 7748 26744
rect 7800 26732 7806 26784
rect 8941 26775 8999 26781
rect 8941 26741 8953 26775
rect 8987 26772 8999 26775
rect 9306 26772 9312 26784
rect 8987 26744 9312 26772
rect 8987 26741 8999 26744
rect 8941 26735 8999 26741
rect 9306 26732 9312 26744
rect 9364 26732 9370 26784
rect 15378 26772 15384 26784
rect 15339 26744 15384 26772
rect 15378 26732 15384 26744
rect 15436 26732 15442 26784
rect 16666 26732 16672 26784
rect 16724 26772 16730 26784
rect 17221 26775 17279 26781
rect 17221 26772 17233 26775
rect 16724 26744 17233 26772
rect 16724 26732 16730 26744
rect 17221 26741 17233 26744
rect 17267 26741 17279 26775
rect 20990 26772 20996 26784
rect 20951 26744 20996 26772
rect 17221 26735 17279 26741
rect 20990 26732 20996 26744
rect 21048 26732 21054 26784
rect 23934 26772 23940 26784
rect 23895 26744 23940 26772
rect 23934 26732 23940 26744
rect 23992 26732 23998 26784
rect 25038 26732 25044 26784
rect 25096 26772 25102 26784
rect 25225 26775 25283 26781
rect 25225 26772 25237 26775
rect 25096 26744 25237 26772
rect 25096 26732 25102 26744
rect 25225 26741 25237 26744
rect 25271 26741 25283 26775
rect 25225 26735 25283 26741
rect 31846 26732 31852 26784
rect 31904 26772 31910 26784
rect 32493 26775 32551 26781
rect 32493 26772 32505 26775
rect 31904 26744 32505 26772
rect 31904 26732 31910 26744
rect 32493 26741 32505 26744
rect 32539 26741 32551 26775
rect 32493 26735 32551 26741
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 9769 26571 9827 26577
rect 9769 26537 9781 26571
rect 9815 26568 9827 26571
rect 10778 26568 10784 26580
rect 9815 26540 10784 26568
rect 9815 26537 9827 26540
rect 9769 26531 9827 26537
rect 10778 26528 10784 26540
rect 10836 26528 10842 26580
rect 12069 26571 12127 26577
rect 12069 26537 12081 26571
rect 12115 26568 12127 26571
rect 12894 26568 12900 26580
rect 12115 26540 12900 26568
rect 12115 26537 12127 26540
rect 12069 26531 12127 26537
rect 12894 26528 12900 26540
rect 12952 26528 12958 26580
rect 13538 26568 13544 26580
rect 13499 26540 13544 26568
rect 13538 26528 13544 26540
rect 13596 26528 13602 26580
rect 14553 26571 14611 26577
rect 14553 26537 14565 26571
rect 14599 26568 14611 26571
rect 14918 26568 14924 26580
rect 14599 26540 14924 26568
rect 14599 26537 14611 26540
rect 14553 26531 14611 26537
rect 14918 26528 14924 26540
rect 14976 26528 14982 26580
rect 17586 26568 17592 26580
rect 17547 26540 17592 26568
rect 17586 26528 17592 26540
rect 17644 26528 17650 26580
rect 20070 26528 20076 26580
rect 20128 26568 20134 26580
rect 20165 26571 20223 26577
rect 20165 26568 20177 26571
rect 20128 26540 20177 26568
rect 20128 26528 20134 26540
rect 20165 26537 20177 26540
rect 20211 26537 20223 26571
rect 27798 26568 27804 26580
rect 27759 26540 27804 26568
rect 20165 26531 20223 26537
rect 27798 26528 27804 26540
rect 27856 26528 27862 26580
rect 12713 26503 12771 26509
rect 12713 26500 12725 26503
rect 12406 26472 12725 26500
rect 7742 26392 7748 26444
rect 7800 26432 7806 26444
rect 9125 26435 9183 26441
rect 9125 26432 9137 26435
rect 7800 26404 9137 26432
rect 7800 26392 7806 26404
rect 9125 26401 9137 26404
rect 9171 26401 9183 26435
rect 9306 26432 9312 26444
rect 9267 26404 9312 26432
rect 9125 26395 9183 26401
rect 9306 26392 9312 26404
rect 9364 26392 9370 26444
rect 12253 26367 12311 26373
rect 12253 26333 12265 26367
rect 12299 26364 12311 26367
rect 12406 26364 12434 26472
rect 12713 26469 12725 26472
rect 12759 26469 12771 26503
rect 12713 26463 12771 26469
rect 15378 26460 15384 26512
rect 15436 26500 15442 26512
rect 15436 26472 17172 26500
rect 15436 26460 15442 26472
rect 16482 26432 16488 26444
rect 16443 26404 16488 26432
rect 16482 26392 16488 26404
rect 16540 26392 16546 26444
rect 16666 26432 16672 26444
rect 16627 26404 16672 26432
rect 16666 26392 16672 26404
rect 16724 26392 16730 26444
rect 17144 26441 17172 26472
rect 18138 26460 18144 26512
rect 18196 26500 18202 26512
rect 24486 26500 24492 26512
rect 18196 26472 24492 26500
rect 18196 26460 18202 26472
rect 24486 26460 24492 26472
rect 24544 26460 24550 26512
rect 24949 26503 25007 26509
rect 24949 26469 24961 26503
rect 24995 26500 25007 26503
rect 26326 26500 26332 26512
rect 24995 26472 26332 26500
rect 24995 26469 25007 26472
rect 24949 26463 25007 26469
rect 26326 26460 26332 26472
rect 26384 26460 26390 26512
rect 17129 26435 17187 26441
rect 17129 26401 17141 26435
rect 17175 26432 17187 26435
rect 20901 26435 20959 26441
rect 20901 26432 20913 26435
rect 17175 26404 20913 26432
rect 17175 26401 17187 26404
rect 17129 26395 17187 26401
rect 20901 26401 20913 26404
rect 20947 26401 20959 26435
rect 20901 26395 20959 26401
rect 21545 26435 21603 26441
rect 21545 26401 21557 26435
rect 21591 26432 21603 26435
rect 24210 26432 24216 26444
rect 21591 26404 24216 26432
rect 21591 26401 21603 26404
rect 21545 26395 21603 26401
rect 24210 26392 24216 26404
rect 24268 26432 24274 26444
rect 24762 26432 24768 26444
rect 24268 26404 24768 26432
rect 24268 26392 24274 26404
rect 24762 26392 24768 26404
rect 24820 26392 24826 26444
rect 25958 26432 25964 26444
rect 25919 26404 25964 26432
rect 25958 26392 25964 26404
rect 26016 26392 26022 26444
rect 26145 26435 26203 26441
rect 26145 26401 26157 26435
rect 26191 26432 26203 26435
rect 27154 26432 27160 26444
rect 26191 26404 27160 26432
rect 26191 26401 26203 26404
rect 26145 26395 26203 26401
rect 27154 26392 27160 26404
rect 27212 26392 27218 26444
rect 12299 26336 12434 26364
rect 12897 26367 12955 26373
rect 12299 26333 12311 26336
rect 12253 26327 12311 26333
rect 12897 26333 12909 26367
rect 12943 26364 12955 26367
rect 13078 26364 13084 26376
rect 12943 26336 13084 26364
rect 12943 26333 12955 26336
rect 12897 26327 12955 26333
rect 13078 26324 13084 26336
rect 13136 26324 13142 26376
rect 13725 26367 13783 26373
rect 13725 26333 13737 26367
rect 13771 26364 13783 26367
rect 14366 26364 14372 26376
rect 13771 26336 14372 26364
rect 13771 26333 13783 26336
rect 13725 26327 13783 26333
rect 14366 26324 14372 26336
rect 14424 26324 14430 26376
rect 14461 26367 14519 26373
rect 14461 26333 14473 26367
rect 14507 26364 14519 26367
rect 14642 26364 14648 26376
rect 14507 26336 14648 26364
rect 14507 26333 14519 26336
rect 14461 26327 14519 26333
rect 14642 26324 14648 26336
rect 14700 26364 14706 26376
rect 17773 26367 17831 26373
rect 17773 26364 17785 26367
rect 14700 26336 17785 26364
rect 14700 26324 14706 26336
rect 17773 26333 17785 26336
rect 17819 26333 17831 26367
rect 20346 26364 20352 26376
rect 20307 26336 20352 26364
rect 17773 26327 17831 26333
rect 20346 26324 20352 26336
rect 20404 26324 20410 26376
rect 25133 26367 25191 26373
rect 25133 26333 25145 26367
rect 25179 26364 25191 26367
rect 25314 26364 25320 26376
rect 25179 26336 25320 26364
rect 25179 26333 25191 26336
rect 25133 26327 25191 26333
rect 25314 26324 25320 26336
rect 25372 26324 25378 26376
rect 26605 26367 26663 26373
rect 26605 26333 26617 26367
rect 26651 26364 26663 26367
rect 27433 26367 27491 26373
rect 27433 26364 27445 26367
rect 26651 26336 27445 26364
rect 26651 26333 26663 26336
rect 26605 26327 26663 26333
rect 27433 26333 27445 26336
rect 27479 26333 27491 26367
rect 27433 26327 27491 26333
rect 20990 26256 20996 26308
rect 21048 26296 21054 26308
rect 27448 26296 27476 26327
rect 27522 26324 27528 26376
rect 27580 26364 27586 26376
rect 27617 26367 27675 26373
rect 27617 26364 27629 26367
rect 27580 26336 27629 26364
rect 27580 26324 27586 26336
rect 27617 26333 27629 26336
rect 27663 26333 27675 26367
rect 27617 26327 27675 26333
rect 28813 26367 28871 26373
rect 28813 26333 28825 26367
rect 28859 26364 28871 26367
rect 37734 26364 37740 26376
rect 28859 26336 37740 26364
rect 28859 26333 28871 26336
rect 28813 26327 28871 26333
rect 37734 26324 37740 26336
rect 37792 26324 37798 26376
rect 27798 26296 27804 26308
rect 21048 26268 21093 26296
rect 27448 26268 27804 26296
rect 21048 26256 21054 26268
rect 27798 26256 27804 26268
rect 27856 26256 27862 26308
rect 27890 26256 27896 26308
rect 27948 26296 27954 26308
rect 28905 26299 28963 26305
rect 28905 26296 28917 26299
rect 27948 26268 28917 26296
rect 27948 26256 27954 26268
rect 28905 26265 28917 26268
rect 28951 26265 28963 26299
rect 28905 26259 28963 26265
rect 7282 26228 7288 26240
rect 7243 26200 7288 26228
rect 7282 26188 7288 26200
rect 7340 26188 7346 26240
rect 23014 26188 23020 26240
rect 23072 26228 23078 26240
rect 23109 26231 23167 26237
rect 23109 26228 23121 26231
rect 23072 26200 23121 26228
rect 23072 26188 23078 26200
rect 23109 26197 23121 26200
rect 23155 26197 23167 26231
rect 23109 26191 23167 26197
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 7742 25984 7748 26036
rect 7800 26024 7806 26036
rect 7929 26027 7987 26033
rect 7929 26024 7941 26027
rect 7800 25996 7941 26024
rect 7800 25984 7806 25996
rect 7929 25993 7941 25996
rect 7975 25993 7987 26027
rect 14366 26024 14372 26036
rect 14327 25996 14372 26024
rect 7929 25987 7987 25993
rect 14366 25984 14372 25996
rect 14424 25984 14430 26036
rect 18877 26027 18935 26033
rect 15304 25996 15700 26024
rect 8938 25956 8944 25968
rect 8899 25928 8944 25956
rect 8938 25916 8944 25928
rect 8996 25916 9002 25968
rect 9033 25959 9091 25965
rect 9033 25925 9045 25959
rect 9079 25956 9091 25959
rect 9766 25956 9772 25968
rect 9079 25928 9772 25956
rect 9079 25925 9091 25928
rect 9033 25919 9091 25925
rect 9766 25916 9772 25928
rect 9824 25916 9830 25968
rect 7282 25888 7288 25900
rect 7243 25860 7288 25888
rect 7282 25848 7288 25860
rect 7340 25848 7346 25900
rect 7469 25891 7527 25897
rect 7469 25857 7481 25891
rect 7515 25888 7527 25891
rect 7834 25888 7840 25900
rect 7515 25860 7840 25888
rect 7515 25857 7527 25860
rect 7469 25851 7527 25857
rect 7834 25848 7840 25860
rect 7892 25848 7898 25900
rect 11149 25891 11207 25897
rect 11149 25857 11161 25891
rect 11195 25888 11207 25891
rect 11514 25888 11520 25900
rect 11195 25860 11520 25888
rect 11195 25857 11207 25860
rect 11149 25851 11207 25857
rect 11514 25848 11520 25860
rect 11572 25848 11578 25900
rect 11698 25888 11704 25900
rect 11659 25860 11704 25888
rect 11698 25848 11704 25860
rect 11756 25848 11762 25900
rect 13630 25888 13636 25900
rect 11808 25860 13492 25888
rect 13591 25860 13636 25888
rect 9585 25823 9643 25829
rect 9585 25789 9597 25823
rect 9631 25820 9643 25823
rect 11808 25820 11836 25860
rect 9631 25792 11836 25820
rect 11885 25823 11943 25829
rect 9631 25789 9643 25792
rect 9585 25783 9643 25789
rect 11885 25789 11897 25823
rect 11931 25789 11943 25823
rect 11885 25783 11943 25789
rect 10962 25684 10968 25696
rect 10923 25656 10968 25684
rect 10962 25644 10968 25656
rect 11020 25644 11026 25696
rect 11900 25684 11928 25783
rect 12710 25780 12716 25832
rect 12768 25820 12774 25832
rect 12805 25823 12863 25829
rect 12805 25820 12817 25823
rect 12768 25792 12817 25820
rect 12768 25780 12774 25792
rect 12805 25789 12817 25792
rect 12851 25789 12863 25823
rect 12805 25783 12863 25789
rect 12345 25755 12403 25761
rect 12345 25721 12357 25755
rect 12391 25752 12403 25755
rect 13354 25752 13360 25764
rect 12391 25724 13360 25752
rect 12391 25721 12403 25724
rect 12345 25715 12403 25721
rect 13354 25712 13360 25724
rect 13412 25712 13418 25764
rect 13464 25752 13492 25860
rect 13630 25848 13636 25860
rect 13688 25848 13694 25900
rect 14274 25848 14280 25900
rect 14332 25888 14338 25900
rect 14553 25891 14611 25897
rect 14553 25888 14565 25891
rect 14332 25860 14565 25888
rect 14332 25848 14338 25860
rect 14553 25857 14565 25860
rect 14599 25888 14611 25891
rect 15304 25888 15332 25996
rect 15470 25916 15476 25968
rect 15528 25956 15534 25968
rect 15565 25959 15623 25965
rect 15565 25956 15577 25959
rect 15528 25928 15577 25956
rect 15528 25916 15534 25928
rect 15565 25925 15577 25928
rect 15611 25925 15623 25959
rect 15672 25956 15700 25996
rect 18877 25993 18889 26027
rect 18923 26024 18935 26027
rect 19334 26024 19340 26036
rect 18923 25996 19340 26024
rect 18923 25993 18935 25996
rect 18877 25987 18935 25993
rect 19334 25984 19340 25996
rect 19392 25984 19398 26036
rect 20165 26027 20223 26033
rect 20165 25993 20177 26027
rect 20211 26024 20223 26027
rect 20346 26024 20352 26036
rect 20211 25996 20352 26024
rect 20211 25993 20223 25996
rect 20165 25987 20223 25993
rect 20346 25984 20352 25996
rect 20404 25984 20410 26036
rect 20809 26027 20867 26033
rect 20809 25993 20821 26027
rect 20855 26024 20867 26027
rect 21174 26024 21180 26036
rect 20855 25996 21180 26024
rect 20855 25993 20867 25996
rect 20809 25987 20867 25993
rect 21174 25984 21180 25996
rect 21232 25984 21238 26036
rect 26145 26027 26203 26033
rect 24044 25996 24440 26024
rect 21266 25956 21272 25968
rect 15672 25928 21272 25956
rect 15565 25919 15623 25925
rect 21266 25916 21272 25928
rect 21324 25916 21330 25968
rect 23014 25956 23020 25968
rect 22975 25928 23020 25956
rect 23014 25916 23020 25928
rect 23072 25916 23078 25968
rect 23109 25959 23167 25965
rect 23109 25925 23121 25959
rect 23155 25956 23167 25959
rect 23934 25956 23940 25968
rect 23155 25928 23940 25956
rect 23155 25925 23167 25928
rect 23109 25919 23167 25925
rect 23934 25916 23940 25928
rect 23992 25916 23998 25968
rect 14599 25860 15332 25888
rect 16117 25891 16175 25897
rect 14599 25857 14611 25860
rect 14553 25851 14611 25857
rect 16117 25857 16129 25891
rect 16163 25888 16175 25891
rect 16574 25888 16580 25900
rect 16163 25860 16580 25888
rect 16163 25857 16175 25860
rect 16117 25851 16175 25857
rect 16574 25848 16580 25860
rect 16632 25848 16638 25900
rect 19061 25891 19119 25897
rect 19061 25857 19073 25891
rect 19107 25888 19119 25891
rect 19334 25888 19340 25900
rect 19107 25860 19340 25888
rect 19107 25857 19119 25860
rect 19061 25851 19119 25857
rect 19334 25848 19340 25860
rect 19392 25848 19398 25900
rect 20346 25888 20352 25900
rect 20307 25860 20352 25888
rect 20346 25848 20352 25860
rect 20404 25848 20410 25900
rect 20993 25891 21051 25897
rect 20993 25857 21005 25891
rect 21039 25888 21051 25891
rect 22830 25888 22836 25900
rect 21039 25860 22836 25888
rect 21039 25857 21051 25860
rect 20993 25851 21051 25857
rect 22830 25848 22836 25860
rect 22888 25848 22894 25900
rect 23661 25891 23719 25897
rect 23661 25857 23673 25891
rect 23707 25888 23719 25891
rect 24044 25888 24072 25996
rect 24302 25956 24308 25968
rect 24263 25928 24308 25956
rect 24302 25916 24308 25928
rect 24360 25916 24366 25968
rect 24412 25956 24440 25996
rect 26145 25993 26157 26027
rect 26191 26024 26203 26027
rect 27522 26024 27528 26036
rect 26191 25996 27528 26024
rect 26191 25993 26203 25996
rect 26145 25987 26203 25993
rect 27522 25984 27528 25996
rect 27580 25984 27586 26036
rect 27798 26024 27804 26036
rect 27759 25996 27804 26024
rect 27798 25984 27804 25996
rect 27856 25984 27862 26036
rect 26418 25956 26424 25968
rect 24412 25928 26424 25956
rect 26418 25916 26424 25928
rect 26476 25916 26482 25968
rect 26326 25888 26332 25900
rect 23707 25860 24072 25888
rect 26287 25860 26332 25888
rect 23707 25857 23719 25860
rect 23661 25851 23719 25857
rect 15194 25780 15200 25832
rect 15252 25820 15258 25832
rect 15473 25823 15531 25829
rect 15473 25820 15485 25823
rect 15252 25792 15485 25820
rect 15252 25780 15258 25792
rect 15473 25789 15485 25792
rect 15519 25820 15531 25823
rect 16206 25820 16212 25832
rect 15519 25792 16212 25820
rect 15519 25789 15531 25792
rect 15473 25783 15531 25789
rect 16206 25780 16212 25792
rect 16264 25780 16270 25832
rect 23474 25780 23480 25832
rect 23532 25820 23538 25832
rect 23676 25820 23704 25851
rect 26326 25848 26332 25860
rect 26384 25848 26390 25900
rect 27157 25891 27215 25897
rect 27157 25857 27169 25891
rect 27203 25888 27215 25891
rect 27798 25888 27804 25900
rect 27203 25860 27804 25888
rect 27203 25857 27215 25860
rect 27157 25851 27215 25857
rect 27798 25848 27804 25860
rect 27856 25848 27862 25900
rect 23532 25792 23704 25820
rect 24213 25823 24271 25829
rect 23532 25780 23538 25792
rect 24213 25789 24225 25823
rect 24259 25789 24271 25823
rect 24486 25820 24492 25832
rect 24447 25792 24492 25820
rect 24213 25783 24271 25789
rect 24228 25752 24256 25783
rect 24486 25780 24492 25792
rect 24544 25780 24550 25832
rect 27338 25820 27344 25832
rect 27299 25792 27344 25820
rect 27338 25780 27344 25792
rect 27396 25780 27402 25832
rect 27706 25752 27712 25764
rect 13464 25724 15976 25752
rect 24228 25724 27712 25752
rect 13449 25687 13507 25693
rect 13449 25684 13461 25687
rect 11900 25656 13461 25684
rect 13449 25653 13461 25656
rect 13495 25653 13507 25687
rect 15948 25684 15976 25724
rect 27706 25712 27712 25724
rect 27764 25752 27770 25764
rect 28442 25752 28448 25764
rect 27764 25724 28448 25752
rect 27764 25712 27770 25724
rect 28442 25712 28448 25724
rect 28500 25712 28506 25764
rect 19978 25684 19984 25696
rect 15948 25656 19984 25684
rect 13449 25647 13507 25653
rect 19978 25644 19984 25656
rect 20036 25644 20042 25696
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 8294 25480 8300 25492
rect 8255 25452 8300 25480
rect 8294 25440 8300 25452
rect 8352 25440 8358 25492
rect 9766 25480 9772 25492
rect 9727 25452 9772 25480
rect 9766 25440 9772 25452
rect 9824 25440 9830 25492
rect 11514 25480 11520 25492
rect 11475 25452 11520 25480
rect 11514 25440 11520 25452
rect 11572 25440 11578 25492
rect 13357 25483 13415 25489
rect 13357 25449 13369 25483
rect 13403 25480 13415 25483
rect 15194 25480 15200 25492
rect 13403 25452 15200 25480
rect 13403 25449 13415 25452
rect 13357 25443 13415 25449
rect 15194 25440 15200 25452
rect 15252 25440 15258 25492
rect 15470 25480 15476 25492
rect 15431 25452 15476 25480
rect 15470 25440 15476 25452
rect 15528 25440 15534 25492
rect 16114 25480 16120 25492
rect 16075 25452 16120 25480
rect 16114 25440 16120 25452
rect 16172 25440 16178 25492
rect 38102 25480 38108 25492
rect 28368 25452 38108 25480
rect 16761 25415 16819 25421
rect 16761 25381 16773 25415
rect 16807 25381 16819 25415
rect 16761 25375 16819 25381
rect 20073 25415 20131 25421
rect 20073 25381 20085 25415
rect 20119 25412 20131 25415
rect 23474 25412 23480 25424
rect 20119 25384 23480 25412
rect 20119 25381 20131 25384
rect 20073 25375 20131 25381
rect 12710 25344 12716 25356
rect 12671 25316 12716 25344
rect 12710 25304 12716 25316
rect 12768 25304 12774 25356
rect 12894 25344 12900 25356
rect 12855 25316 12900 25344
rect 12894 25304 12900 25316
rect 12952 25304 12958 25356
rect 16776 25344 16804 25375
rect 23474 25372 23480 25384
rect 23532 25372 23538 25424
rect 25038 25344 25044 25356
rect 15672 25316 16804 25344
rect 24999 25316 25044 25344
rect 1762 25276 1768 25288
rect 1723 25248 1768 25276
rect 1762 25236 1768 25248
rect 1820 25236 1826 25288
rect 6178 25236 6184 25288
rect 6236 25276 6242 25288
rect 6730 25276 6736 25288
rect 6236 25248 6736 25276
rect 6236 25236 6242 25248
rect 6730 25236 6736 25248
rect 6788 25276 6794 25288
rect 8205 25279 8263 25285
rect 8205 25276 8217 25279
rect 6788 25248 8217 25276
rect 6788 25236 6794 25248
rect 8205 25245 8217 25248
rect 8251 25245 8263 25279
rect 9950 25276 9956 25288
rect 9911 25248 9956 25276
rect 8205 25239 8263 25245
rect 9950 25236 9956 25248
rect 10008 25236 10014 25288
rect 11698 25276 11704 25288
rect 11659 25248 11704 25276
rect 11698 25236 11704 25248
rect 11756 25236 11762 25288
rect 15672 25285 15700 25316
rect 25038 25304 25044 25316
rect 25096 25304 25102 25356
rect 15657 25279 15715 25285
rect 15657 25245 15669 25279
rect 15703 25245 15715 25279
rect 15657 25239 15715 25245
rect 16301 25279 16359 25285
rect 16301 25245 16313 25279
rect 16347 25276 16359 25279
rect 16758 25276 16764 25288
rect 16347 25248 16764 25276
rect 16347 25245 16359 25248
rect 16301 25239 16359 25245
rect 16758 25236 16764 25248
rect 16816 25236 16822 25288
rect 16850 25236 16856 25288
rect 16908 25276 16914 25288
rect 16945 25279 17003 25285
rect 16945 25276 16957 25279
rect 16908 25248 16957 25276
rect 16908 25236 16914 25248
rect 16945 25245 16957 25248
rect 16991 25245 17003 25279
rect 16945 25239 17003 25245
rect 18414 25236 18420 25288
rect 18472 25276 18478 25288
rect 18690 25276 18696 25288
rect 18472 25248 18696 25276
rect 18472 25236 18478 25248
rect 18690 25236 18696 25248
rect 18748 25236 18754 25288
rect 28368 25285 28396 25452
rect 38102 25440 38108 25452
rect 38160 25440 38166 25492
rect 28442 25372 28448 25424
rect 28500 25412 28506 25424
rect 32122 25412 32128 25424
rect 28500 25384 28545 25412
rect 32083 25384 32128 25412
rect 28500 25372 28506 25384
rect 32122 25372 32128 25384
rect 32180 25372 32186 25424
rect 31754 25344 31760 25356
rect 31715 25316 31760 25344
rect 31754 25304 31760 25316
rect 31812 25304 31818 25356
rect 28353 25279 28411 25285
rect 28353 25245 28365 25279
rect 28399 25245 28411 25279
rect 31938 25276 31944 25288
rect 31899 25248 31944 25276
rect 28353 25239 28411 25245
rect 31938 25236 31944 25248
rect 31996 25236 32002 25288
rect 38286 25276 38292 25288
rect 38247 25248 38292 25276
rect 38286 25236 38292 25248
rect 38344 25236 38350 25288
rect 13354 25168 13360 25220
rect 13412 25208 13418 25220
rect 17862 25208 17868 25220
rect 13412 25180 17868 25208
rect 13412 25168 13418 25180
rect 17862 25168 17868 25180
rect 17920 25208 17926 25220
rect 19521 25211 19579 25217
rect 19521 25208 19533 25211
rect 17920 25180 19533 25208
rect 17920 25168 17926 25180
rect 19521 25177 19533 25180
rect 19567 25177 19579 25211
rect 19521 25171 19579 25177
rect 19613 25211 19671 25217
rect 19613 25177 19625 25211
rect 19659 25177 19671 25211
rect 19613 25171 19671 25177
rect 1581 25143 1639 25149
rect 1581 25109 1593 25143
rect 1627 25140 1639 25143
rect 3142 25140 3148 25152
rect 1627 25112 3148 25140
rect 1627 25109 1639 25112
rect 1581 25103 1639 25109
rect 3142 25100 3148 25112
rect 3200 25100 3206 25152
rect 18785 25143 18843 25149
rect 18785 25109 18797 25143
rect 18831 25140 18843 25143
rect 19628 25140 19656 25171
rect 25130 25168 25136 25220
rect 25188 25208 25194 25220
rect 25685 25211 25743 25217
rect 25188 25180 25233 25208
rect 25188 25168 25194 25180
rect 25685 25177 25697 25211
rect 25731 25208 25743 25211
rect 27614 25208 27620 25220
rect 25731 25180 27620 25208
rect 25731 25177 25743 25180
rect 25685 25171 25743 25177
rect 27614 25168 27620 25180
rect 27672 25168 27678 25220
rect 38102 25140 38108 25152
rect 18831 25112 19656 25140
rect 38063 25112 38108 25140
rect 18831 25109 18843 25112
rect 18785 25103 18843 25109
rect 38102 25100 38108 25112
rect 38160 25100 38166 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 9950 24896 9956 24948
rect 10008 24936 10014 24948
rect 10873 24939 10931 24945
rect 10873 24936 10885 24939
rect 10008 24908 10885 24936
rect 10008 24896 10014 24908
rect 10873 24905 10885 24908
rect 10919 24905 10931 24939
rect 10873 24899 10931 24905
rect 12345 24939 12403 24945
rect 12345 24905 12357 24939
rect 12391 24936 12403 24939
rect 13630 24936 13636 24948
rect 12391 24908 13636 24936
rect 12391 24905 12403 24908
rect 12345 24899 12403 24905
rect 13630 24896 13636 24908
rect 13688 24896 13694 24948
rect 21910 24896 21916 24948
rect 21968 24936 21974 24948
rect 27249 24939 27307 24945
rect 21968 24908 27200 24936
rect 21968 24896 21974 24908
rect 14918 24868 14924 24880
rect 14879 24840 14924 24868
rect 14918 24828 14924 24840
rect 14976 24828 14982 24880
rect 22186 24868 22192 24880
rect 22147 24840 22192 24868
rect 22186 24828 22192 24840
rect 22244 24828 22250 24880
rect 27172 24868 27200 24908
rect 27249 24905 27261 24939
rect 27295 24936 27307 24939
rect 27338 24936 27344 24948
rect 27295 24908 27344 24936
rect 27295 24905 27307 24908
rect 27249 24899 27307 24905
rect 27338 24896 27344 24908
rect 27396 24896 27402 24948
rect 27982 24868 27988 24880
rect 27172 24840 27988 24868
rect 5350 24800 5356 24812
rect 5311 24772 5356 24800
rect 5350 24760 5356 24772
rect 5408 24760 5414 24812
rect 6270 24760 6276 24812
rect 6328 24800 6334 24812
rect 7561 24803 7619 24809
rect 7561 24800 7573 24803
rect 6328 24772 7573 24800
rect 6328 24760 6334 24772
rect 7561 24769 7573 24772
rect 7607 24769 7619 24803
rect 7561 24763 7619 24769
rect 10778 24760 10784 24812
rect 10836 24800 10842 24812
rect 11057 24803 11115 24809
rect 11057 24800 11069 24803
rect 10836 24772 11069 24800
rect 10836 24760 10842 24772
rect 11057 24769 11069 24772
rect 11103 24769 11115 24803
rect 11057 24763 11115 24769
rect 12529 24803 12587 24809
rect 12529 24769 12541 24803
rect 12575 24800 12587 24803
rect 12894 24800 12900 24812
rect 12575 24772 12900 24800
rect 12575 24769 12587 24772
rect 12529 24763 12587 24769
rect 12894 24760 12900 24772
rect 12952 24760 12958 24812
rect 12989 24803 13047 24809
rect 12989 24769 13001 24803
rect 13035 24800 13047 24803
rect 13446 24800 13452 24812
rect 13035 24772 13452 24800
rect 13035 24769 13047 24772
rect 12989 24763 13047 24769
rect 12618 24692 12624 24744
rect 12676 24732 12682 24744
rect 13004 24732 13032 24763
rect 13446 24760 13452 24772
rect 13504 24760 13510 24812
rect 27172 24809 27200 24840
rect 27982 24828 27988 24840
rect 28040 24828 28046 24880
rect 27157 24803 27215 24809
rect 27157 24769 27169 24803
rect 27203 24769 27215 24803
rect 27157 24763 27215 24769
rect 12676 24704 13032 24732
rect 13173 24735 13231 24741
rect 12676 24692 12682 24704
rect 13173 24701 13185 24735
rect 13219 24732 13231 24735
rect 13354 24732 13360 24744
rect 13219 24704 13360 24732
rect 13219 24701 13231 24704
rect 13173 24695 13231 24701
rect 13354 24692 13360 24704
rect 13412 24692 13418 24744
rect 14826 24732 14832 24744
rect 14787 24704 14832 24732
rect 14826 24692 14832 24704
rect 14884 24692 14890 24744
rect 15470 24732 15476 24744
rect 15431 24704 15476 24732
rect 15470 24692 15476 24704
rect 15528 24692 15534 24744
rect 19610 24692 19616 24744
rect 19668 24732 19674 24744
rect 22097 24735 22155 24741
rect 22097 24732 22109 24735
rect 19668 24704 22109 24732
rect 19668 24692 19674 24704
rect 22097 24701 22109 24704
rect 22143 24732 22155 24735
rect 28258 24732 28264 24744
rect 22143 24704 28264 24732
rect 22143 24701 22155 24704
rect 22097 24695 22155 24701
rect 28258 24692 28264 24704
rect 28316 24692 28322 24744
rect 14550 24624 14556 24676
rect 14608 24664 14614 24676
rect 21910 24664 21916 24676
rect 14608 24636 21916 24664
rect 14608 24624 14614 24636
rect 21910 24624 21916 24636
rect 21968 24624 21974 24676
rect 22646 24664 22652 24676
rect 22607 24636 22652 24664
rect 22646 24624 22652 24636
rect 22704 24624 22710 24676
rect 5350 24556 5356 24608
rect 5408 24596 5414 24608
rect 5445 24599 5503 24605
rect 5445 24596 5457 24599
rect 5408 24568 5457 24596
rect 5408 24556 5414 24568
rect 5445 24565 5457 24568
rect 5491 24565 5503 24599
rect 5445 24559 5503 24565
rect 7653 24599 7711 24605
rect 7653 24565 7665 24599
rect 7699 24596 7711 24599
rect 8386 24596 8392 24608
rect 7699 24568 8392 24596
rect 7699 24565 7711 24568
rect 7653 24559 7711 24565
rect 8386 24556 8392 24568
rect 8444 24556 8450 24608
rect 12802 24556 12808 24608
rect 12860 24596 12866 24608
rect 13357 24599 13415 24605
rect 13357 24596 13369 24599
rect 12860 24568 13369 24596
rect 12860 24556 12866 24568
rect 13357 24565 13369 24568
rect 13403 24565 13415 24599
rect 13357 24559 13415 24565
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 4249 24395 4307 24401
rect 4249 24361 4261 24395
rect 4295 24392 4307 24395
rect 4614 24392 4620 24404
rect 4295 24364 4620 24392
rect 4295 24361 4307 24364
rect 4249 24355 4307 24361
rect 4614 24352 4620 24364
rect 4672 24352 4678 24404
rect 14918 24352 14924 24404
rect 14976 24392 14982 24404
rect 15933 24395 15991 24401
rect 15933 24392 15945 24395
rect 14976 24364 15945 24392
rect 14976 24352 14982 24364
rect 15933 24361 15945 24364
rect 15979 24361 15991 24395
rect 15933 24355 15991 24361
rect 20809 24395 20867 24401
rect 20809 24361 20821 24395
rect 20855 24392 20867 24395
rect 20898 24392 20904 24404
rect 20855 24364 20904 24392
rect 20855 24361 20867 24364
rect 20809 24355 20867 24361
rect 20898 24352 20904 24364
rect 20956 24352 20962 24404
rect 24765 24395 24823 24401
rect 24765 24361 24777 24395
rect 24811 24392 24823 24395
rect 25130 24392 25136 24404
rect 24811 24364 25136 24392
rect 24811 24361 24823 24364
rect 24765 24355 24823 24361
rect 25130 24352 25136 24364
rect 25188 24352 25194 24404
rect 31938 24352 31944 24404
rect 31996 24392 32002 24404
rect 32033 24395 32091 24401
rect 32033 24392 32045 24395
rect 31996 24364 32045 24392
rect 31996 24352 32002 24364
rect 32033 24361 32045 24364
rect 32079 24361 32091 24395
rect 32033 24355 32091 24361
rect 13449 24327 13507 24333
rect 13449 24293 13461 24327
rect 13495 24293 13507 24327
rect 22554 24324 22560 24336
rect 13449 24287 13507 24293
rect 18248 24296 22560 24324
rect 1578 24188 1584 24200
rect 1539 24160 1584 24188
rect 1578 24148 1584 24160
rect 1636 24148 1642 24200
rect 4157 24191 4215 24197
rect 4157 24157 4169 24191
rect 4203 24157 4215 24191
rect 4157 24151 4215 24157
rect 4172 24120 4200 24151
rect 6362 24148 6368 24200
rect 6420 24188 6426 24200
rect 7561 24191 7619 24197
rect 7561 24188 7573 24191
rect 6420 24160 7573 24188
rect 6420 24148 6426 24160
rect 7561 24157 7573 24160
rect 7607 24157 7619 24191
rect 7742 24188 7748 24200
rect 7703 24160 7748 24188
rect 7561 24151 7619 24157
rect 7742 24148 7748 24160
rect 7800 24148 7806 24200
rect 10778 24148 10784 24200
rect 10836 24188 10842 24200
rect 11149 24191 11207 24197
rect 11149 24188 11161 24191
rect 10836 24160 11161 24188
rect 10836 24148 10842 24160
rect 11149 24157 11161 24160
rect 11195 24157 11207 24191
rect 11149 24151 11207 24157
rect 12989 24191 13047 24197
rect 12989 24157 13001 24191
rect 13035 24188 13047 24191
rect 13464 24188 13492 24287
rect 16666 24256 16672 24268
rect 13648 24228 16672 24256
rect 13648 24200 13676 24228
rect 16666 24216 16672 24228
rect 16724 24216 16730 24268
rect 18248 24265 18276 24296
rect 22554 24284 22560 24296
rect 22612 24284 22618 24336
rect 18233 24259 18291 24265
rect 18233 24225 18245 24259
rect 18279 24225 18291 24259
rect 18874 24256 18880 24268
rect 18835 24228 18880 24256
rect 18233 24219 18291 24225
rect 18874 24216 18880 24228
rect 18932 24216 18938 24268
rect 19610 24256 19616 24268
rect 19571 24228 19616 24256
rect 19610 24216 19616 24228
rect 19668 24216 19674 24268
rect 19978 24256 19984 24268
rect 19939 24228 19984 24256
rect 19978 24216 19984 24228
rect 20036 24216 20042 24268
rect 20806 24216 20812 24268
rect 20864 24256 20870 24268
rect 22646 24256 22652 24268
rect 20864 24228 22652 24256
rect 20864 24216 20870 24228
rect 22646 24216 22652 24228
rect 22704 24256 22710 24268
rect 25409 24259 25467 24265
rect 25409 24256 25421 24259
rect 22704 24228 25421 24256
rect 22704 24216 22710 24228
rect 25409 24225 25421 24228
rect 25455 24225 25467 24259
rect 25409 24219 25467 24225
rect 26053 24259 26111 24265
rect 26053 24225 26065 24259
rect 26099 24256 26111 24259
rect 26234 24256 26240 24268
rect 26099 24228 26240 24256
rect 26099 24225 26111 24228
rect 26053 24219 26111 24225
rect 26234 24216 26240 24228
rect 26292 24216 26298 24268
rect 38102 24256 38108 24268
rect 28460 24228 38108 24256
rect 13035 24160 13492 24188
rect 13035 24157 13047 24160
rect 12989 24151 13047 24157
rect 13630 24148 13636 24200
rect 13688 24188 13694 24200
rect 16117 24191 16175 24197
rect 13688 24160 13781 24188
rect 13688 24148 13694 24160
rect 16117 24157 16129 24191
rect 16163 24188 16175 24191
rect 16942 24188 16948 24200
rect 16163 24160 16948 24188
rect 16163 24157 16175 24160
rect 16117 24151 16175 24157
rect 16942 24148 16948 24160
rect 17000 24148 17006 24200
rect 20714 24188 20720 24200
rect 20675 24160 20720 24188
rect 20714 24148 20720 24160
rect 20772 24148 20778 24200
rect 21174 24148 21180 24200
rect 21232 24188 21238 24200
rect 22189 24191 22247 24197
rect 22189 24188 22201 24191
rect 21232 24160 22201 24188
rect 21232 24148 21238 24160
rect 22189 24157 22201 24160
rect 22235 24157 22247 24191
rect 22189 24151 22247 24157
rect 24673 24191 24731 24197
rect 24673 24157 24685 24191
rect 24719 24188 24731 24191
rect 24854 24188 24860 24200
rect 24719 24160 24860 24188
rect 24719 24157 24731 24160
rect 24673 24151 24731 24157
rect 24854 24148 24860 24160
rect 24912 24148 24918 24200
rect 28460 24197 28488 24228
rect 38102 24216 38108 24228
rect 38160 24216 38166 24268
rect 28445 24191 28503 24197
rect 28445 24157 28457 24191
rect 28491 24157 28503 24191
rect 28445 24151 28503 24157
rect 31297 24191 31355 24197
rect 31297 24157 31309 24191
rect 31343 24157 31355 24191
rect 31297 24151 31355 24157
rect 7282 24120 7288 24132
rect 4172 24092 7288 24120
rect 7282 24080 7288 24092
rect 7340 24080 7346 24132
rect 11241 24123 11299 24129
rect 11241 24089 11253 24123
rect 11287 24120 11299 24123
rect 11287 24092 16068 24120
rect 11287 24089 11299 24092
rect 11241 24083 11299 24089
rect 1762 24052 1768 24064
rect 1723 24024 1768 24052
rect 1762 24012 1768 24024
rect 1820 24012 1826 24064
rect 8202 24052 8208 24064
rect 8163 24024 8208 24052
rect 8202 24012 8208 24024
rect 8260 24012 8266 24064
rect 10502 24052 10508 24064
rect 10463 24024 10508 24052
rect 10502 24012 10508 24024
rect 10560 24012 10566 24064
rect 12342 24012 12348 24064
rect 12400 24052 12406 24064
rect 12805 24055 12863 24061
rect 12805 24052 12817 24055
rect 12400 24024 12817 24052
rect 12400 24012 12406 24024
rect 12805 24021 12817 24024
rect 12851 24021 12863 24055
rect 16040 24052 16068 24092
rect 18322 24080 18328 24132
rect 18380 24120 18386 24132
rect 19705 24123 19763 24129
rect 18380 24092 18425 24120
rect 18380 24080 18386 24092
rect 19705 24089 19717 24123
rect 19751 24089 19763 24123
rect 19705 24083 19763 24089
rect 25501 24123 25559 24129
rect 25501 24089 25513 24123
rect 25547 24089 25559 24123
rect 31312 24120 31340 24151
rect 31386 24148 31392 24200
rect 31444 24188 31450 24200
rect 31941 24191 31999 24197
rect 31941 24188 31953 24191
rect 31444 24160 31953 24188
rect 31444 24148 31450 24160
rect 31941 24157 31953 24160
rect 31987 24157 31999 24191
rect 38286 24188 38292 24200
rect 38247 24160 38292 24188
rect 31941 24151 31999 24157
rect 38286 24148 38292 24160
rect 38344 24148 38350 24200
rect 25501 24083 25559 24089
rect 25976 24092 31340 24120
rect 19720 24052 19748 24083
rect 16040 24024 19748 24052
rect 22005 24055 22063 24061
rect 12805 24015 12863 24021
rect 22005 24021 22017 24055
rect 22051 24052 22063 24055
rect 22646 24052 22652 24064
rect 22051 24024 22652 24052
rect 22051 24021 22063 24024
rect 22005 24015 22063 24021
rect 22646 24012 22652 24024
rect 22704 24012 22710 24064
rect 24670 24012 24676 24064
rect 24728 24052 24734 24064
rect 25516 24052 25544 24083
rect 25976 24064 26004 24092
rect 24728 24024 25544 24052
rect 24728 24012 24734 24024
rect 25958 24012 25964 24064
rect 26016 24012 26022 24064
rect 28442 24052 28448 24064
rect 28403 24024 28448 24052
rect 28442 24012 28448 24024
rect 28500 24012 28506 24064
rect 31389 24055 31447 24061
rect 31389 24021 31401 24055
rect 31435 24052 31447 24055
rect 33502 24052 33508 24064
rect 31435 24024 33508 24052
rect 31435 24021 31447 24024
rect 31389 24015 31447 24021
rect 33502 24012 33508 24024
rect 33560 24012 33566 24064
rect 36998 24012 37004 24064
rect 37056 24052 37062 24064
rect 38105 24055 38163 24061
rect 38105 24052 38117 24055
rect 37056 24024 38117 24052
rect 37056 24012 37062 24024
rect 38105 24021 38117 24024
rect 38151 24021 38163 24055
rect 38105 24015 38163 24021
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 1578 23808 1584 23860
rect 1636 23848 1642 23860
rect 7101 23851 7159 23857
rect 7101 23848 7113 23851
rect 1636 23820 7113 23848
rect 1636 23808 1642 23820
rect 7101 23817 7113 23820
rect 7147 23817 7159 23851
rect 7101 23811 7159 23817
rect 8202 23808 8208 23860
rect 8260 23848 8266 23860
rect 11149 23851 11207 23857
rect 11149 23848 11161 23851
rect 8260 23820 11161 23848
rect 8260 23808 8266 23820
rect 11149 23817 11161 23820
rect 11195 23817 11207 23851
rect 12802 23848 12808 23860
rect 12763 23820 12808 23848
rect 11149 23811 11207 23817
rect 11164 23780 11192 23811
rect 12802 23808 12808 23820
rect 12860 23808 12866 23860
rect 13354 23848 13360 23860
rect 13315 23820 13360 23848
rect 13354 23808 13360 23820
rect 13412 23808 13418 23860
rect 21361 23851 21419 23857
rect 21361 23817 21373 23851
rect 21407 23848 21419 23851
rect 22186 23848 22192 23860
rect 21407 23820 22192 23848
rect 21407 23817 21419 23820
rect 21361 23811 21419 23817
rect 22186 23808 22192 23820
rect 22244 23808 22250 23860
rect 27798 23848 27804 23860
rect 22388 23820 27804 23848
rect 14366 23780 14372 23792
rect 11164 23752 14372 23780
rect 14366 23740 14372 23752
rect 14424 23740 14430 23792
rect 17034 23780 17040 23792
rect 16995 23752 17040 23780
rect 17034 23740 17040 23752
rect 17092 23740 17098 23792
rect 7285 23715 7343 23721
rect 7285 23681 7297 23715
rect 7331 23712 7343 23715
rect 9214 23712 9220 23724
rect 7331 23684 9220 23712
rect 7331 23681 7343 23684
rect 7285 23675 7343 23681
rect 9214 23672 9220 23684
rect 9272 23672 9278 23724
rect 10502 23712 10508 23724
rect 10463 23684 10508 23712
rect 10502 23672 10508 23684
rect 10560 23672 10566 23724
rect 10689 23715 10747 23721
rect 10689 23681 10701 23715
rect 10735 23712 10747 23715
rect 10962 23712 10968 23724
rect 10735 23684 10968 23712
rect 10735 23681 10747 23684
rect 10689 23675 10747 23681
rect 10962 23672 10968 23684
rect 11020 23672 11026 23724
rect 12342 23712 12348 23724
rect 12303 23684 12348 23712
rect 12342 23672 12348 23684
rect 12400 23672 12406 23724
rect 13265 23715 13323 23721
rect 13265 23681 13277 23715
rect 13311 23712 13323 23715
rect 13630 23712 13636 23724
rect 13311 23684 13636 23712
rect 13311 23681 13323 23684
rect 13265 23675 13323 23681
rect 13630 23672 13636 23684
rect 13688 23672 13694 23724
rect 15010 23712 15016 23724
rect 14971 23684 15016 23712
rect 15010 23672 15016 23684
rect 15068 23672 15074 23724
rect 21266 23712 21272 23724
rect 21227 23684 21272 23712
rect 21266 23672 21272 23684
rect 21324 23672 21330 23724
rect 12158 23644 12164 23656
rect 12119 23616 12164 23644
rect 12158 23604 12164 23616
rect 12216 23604 12222 23656
rect 16666 23604 16672 23656
rect 16724 23644 16730 23656
rect 16945 23647 17003 23653
rect 16945 23644 16957 23647
rect 16724 23616 16957 23644
rect 16724 23604 16730 23616
rect 16945 23613 16957 23616
rect 16991 23644 17003 23647
rect 22388 23644 22416 23820
rect 27798 23808 27804 23820
rect 27856 23848 27862 23860
rect 28534 23848 28540 23860
rect 27856 23820 28540 23848
rect 27856 23808 27862 23820
rect 28534 23808 28540 23820
rect 28592 23808 28598 23860
rect 31757 23851 31815 23857
rect 31757 23817 31769 23851
rect 31803 23848 31815 23851
rect 32122 23848 32128 23860
rect 31803 23820 32128 23848
rect 31803 23817 31815 23820
rect 31757 23811 31815 23817
rect 32122 23808 32128 23820
rect 32180 23808 32186 23860
rect 33318 23848 33324 23860
rect 33279 23820 33324 23848
rect 33318 23808 33324 23820
rect 33376 23808 33382 23860
rect 22646 23780 22652 23792
rect 22607 23752 22652 23780
rect 22646 23740 22652 23752
rect 22704 23740 22710 23792
rect 29178 23712 29184 23724
rect 29139 23684 29184 23712
rect 29178 23672 29184 23684
rect 29236 23672 29242 23724
rect 32490 23712 32496 23724
rect 32451 23684 32496 23712
rect 32490 23672 32496 23684
rect 32548 23672 32554 23724
rect 33502 23712 33508 23724
rect 33463 23684 33508 23712
rect 33502 23672 33508 23684
rect 33560 23672 33566 23724
rect 22557 23647 22615 23653
rect 22557 23644 22569 23647
rect 16991 23616 22094 23644
rect 22388 23616 22569 23644
rect 16991 23613 17003 23616
rect 16945 23607 17003 23613
rect 16574 23536 16580 23588
rect 16632 23576 16638 23588
rect 17497 23579 17555 23585
rect 17497 23576 17509 23579
rect 16632 23548 17509 23576
rect 16632 23536 16638 23548
rect 17497 23545 17509 23548
rect 17543 23545 17555 23579
rect 22066 23576 22094 23616
rect 22557 23613 22569 23616
rect 22603 23613 22615 23647
rect 22557 23607 22615 23613
rect 22833 23647 22891 23653
rect 22833 23613 22845 23647
rect 22879 23613 22891 23647
rect 22833 23607 22891 23613
rect 30469 23647 30527 23653
rect 30469 23613 30481 23647
rect 30515 23644 30527 23647
rect 31113 23647 31171 23653
rect 31113 23644 31125 23647
rect 30515 23616 31125 23644
rect 30515 23613 30527 23616
rect 30469 23607 30527 23613
rect 31113 23613 31125 23616
rect 31159 23613 31171 23647
rect 31113 23607 31171 23613
rect 31297 23647 31355 23653
rect 31297 23613 31309 23647
rect 31343 23644 31355 23647
rect 31343 23616 32352 23644
rect 31343 23613 31355 23616
rect 31297 23607 31355 23613
rect 22848 23576 22876 23607
rect 32324 23585 32352 23616
rect 22066 23548 22876 23576
rect 32309 23579 32367 23585
rect 17497 23539 17555 23545
rect 32309 23545 32321 23579
rect 32355 23545 32367 23579
rect 32309 23539 32367 23545
rect 14458 23468 14464 23520
rect 14516 23508 14522 23520
rect 14829 23511 14887 23517
rect 14829 23508 14841 23511
rect 14516 23480 14841 23508
rect 14516 23468 14522 23480
rect 14829 23477 14841 23480
rect 14875 23477 14887 23511
rect 14829 23471 14887 23477
rect 19978 23468 19984 23520
rect 20036 23508 20042 23520
rect 27246 23508 27252 23520
rect 20036 23480 27252 23508
rect 20036 23468 20042 23480
rect 27246 23468 27252 23480
rect 27304 23468 27310 23520
rect 29270 23508 29276 23520
rect 29231 23480 29276 23508
rect 29270 23468 29276 23480
rect 29328 23468 29334 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 7742 23264 7748 23316
rect 7800 23304 7806 23316
rect 7929 23307 7987 23313
rect 7929 23304 7941 23307
rect 7800 23276 7941 23304
rect 7800 23264 7806 23276
rect 7929 23273 7941 23276
rect 7975 23273 7987 23307
rect 7929 23267 7987 23273
rect 11698 23264 11704 23316
rect 11756 23304 11762 23316
rect 14918 23304 14924 23316
rect 11756 23276 14924 23304
rect 11756 23264 11762 23276
rect 14918 23264 14924 23276
rect 14976 23264 14982 23316
rect 16206 23304 16212 23316
rect 16167 23276 16212 23304
rect 16206 23264 16212 23276
rect 16264 23264 16270 23316
rect 16758 23264 16764 23316
rect 16816 23304 16822 23316
rect 17129 23307 17187 23313
rect 17129 23304 17141 23307
rect 16816 23276 17141 23304
rect 16816 23264 16822 23276
rect 17129 23273 17141 23276
rect 17175 23273 17187 23307
rect 17129 23267 17187 23273
rect 18049 23307 18107 23313
rect 18049 23273 18061 23307
rect 18095 23304 18107 23307
rect 18322 23304 18328 23316
rect 18095 23276 18328 23304
rect 18095 23273 18107 23276
rect 18049 23267 18107 23273
rect 18322 23264 18328 23276
rect 18380 23264 18386 23316
rect 20349 23307 20407 23313
rect 20349 23273 20361 23307
rect 20395 23304 20407 23307
rect 21174 23304 21180 23316
rect 20395 23276 21180 23304
rect 20395 23273 20407 23276
rect 20349 23267 20407 23273
rect 21174 23264 21180 23276
rect 21232 23264 21238 23316
rect 22066 23276 27016 23304
rect 22066 23248 22094 23276
rect 9398 23196 9404 23248
rect 9456 23236 9462 23248
rect 16666 23236 16672 23248
rect 9456 23208 16672 23236
rect 9456 23196 9462 23208
rect 16666 23196 16672 23208
rect 16724 23196 16730 23248
rect 19426 23196 19432 23248
rect 19484 23236 19490 23248
rect 22002 23236 22008 23248
rect 19484 23208 22008 23236
rect 19484 23196 19490 23208
rect 22002 23196 22008 23208
rect 22060 23208 22094 23248
rect 25409 23239 25467 23245
rect 22060 23196 22066 23208
rect 25409 23205 25421 23239
rect 25455 23205 25467 23239
rect 25409 23199 25467 23205
rect 12158 23168 12164 23180
rect 12119 23140 12164 23168
rect 12158 23128 12164 23140
rect 12216 23128 12222 23180
rect 14366 23168 14372 23180
rect 14327 23140 14372 23168
rect 14366 23128 14372 23140
rect 14424 23128 14430 23180
rect 15381 23171 15439 23177
rect 15381 23137 15393 23171
rect 15427 23168 15439 23171
rect 19334 23168 19340 23180
rect 15427 23140 17908 23168
rect 15427 23137 15439 23140
rect 15381 23131 15439 23137
rect 6454 23060 6460 23112
rect 6512 23100 6518 23112
rect 7837 23103 7895 23109
rect 7837 23100 7849 23103
rect 6512 23072 7849 23100
rect 6512 23060 6518 23072
rect 7837 23069 7849 23072
rect 7883 23100 7895 23103
rect 11698 23100 11704 23112
rect 7883 23072 11704 23100
rect 7883 23069 7895 23072
rect 7837 23063 7895 23069
rect 11698 23060 11704 23072
rect 11756 23060 11762 23112
rect 15841 23103 15899 23109
rect 15841 23069 15853 23103
rect 15887 23069 15899 23103
rect 16022 23100 16028 23112
rect 15983 23072 16028 23100
rect 15841 23063 15899 23069
rect 14458 22992 14464 23044
rect 14516 23032 14522 23044
rect 14516 23004 14561 23032
rect 14516 22992 14522 23004
rect 11330 22924 11336 22976
rect 11388 22964 11394 22976
rect 15856 22964 15884 23063
rect 16022 23060 16028 23072
rect 16080 23060 16086 23112
rect 17313 23103 17371 23109
rect 17313 23069 17325 23103
rect 17359 23069 17371 23103
rect 17313 23063 17371 23069
rect 11388 22936 15884 22964
rect 17328 22964 17356 23063
rect 17880 23032 17908 23140
rect 17972 23140 19340 23168
rect 17972 23109 18000 23140
rect 19334 23128 19340 23140
rect 19392 23168 19398 23180
rect 20806 23168 20812 23180
rect 19392 23140 20812 23168
rect 19392 23128 19398 23140
rect 20806 23128 20812 23140
rect 20864 23128 20870 23180
rect 25424 23168 25452 23199
rect 26988 23177 27016 23276
rect 27430 23264 27436 23316
rect 27488 23304 27494 23316
rect 29178 23304 29184 23316
rect 27488 23276 29184 23304
rect 27488 23264 27494 23276
rect 29178 23264 29184 23276
rect 29236 23304 29242 23316
rect 31205 23307 31263 23313
rect 29236 23276 30236 23304
rect 29236 23264 29242 23276
rect 28905 23239 28963 23245
rect 28905 23205 28917 23239
rect 28951 23236 28963 23239
rect 29730 23236 29736 23248
rect 28951 23208 29736 23236
rect 28951 23205 28963 23208
rect 28905 23199 28963 23205
rect 29730 23196 29736 23208
rect 29788 23236 29794 23248
rect 30101 23239 30159 23245
rect 30101 23236 30113 23239
rect 29788 23208 30113 23236
rect 29788 23196 29794 23208
rect 30101 23205 30113 23208
rect 30147 23205 30159 23239
rect 30101 23199 30159 23205
rect 26973 23171 27031 23177
rect 25424 23140 26280 23168
rect 17957 23103 18015 23109
rect 17957 23069 17969 23103
rect 18003 23069 18015 23103
rect 17957 23063 18015 23069
rect 19889 23103 19947 23109
rect 19889 23069 19901 23103
rect 19935 23100 19947 23103
rect 19978 23100 19984 23112
rect 19935 23072 19984 23100
rect 19935 23069 19947 23072
rect 19889 23063 19947 23069
rect 19978 23060 19984 23072
rect 20036 23060 20042 23112
rect 20533 23103 20591 23109
rect 20533 23069 20545 23103
rect 20579 23069 20591 23103
rect 20533 23063 20591 23069
rect 18506 23032 18512 23044
rect 17880 23004 18512 23032
rect 18506 22992 18512 23004
rect 18564 22992 18570 23044
rect 19334 22992 19340 23044
rect 19392 23032 19398 23044
rect 20548 23032 20576 23063
rect 21266 23060 21272 23112
rect 21324 23100 21330 23112
rect 21821 23103 21879 23109
rect 21821 23100 21833 23103
rect 21324 23072 21833 23100
rect 21324 23060 21330 23072
rect 21821 23069 21833 23072
rect 21867 23069 21879 23103
rect 21821 23063 21879 23069
rect 24854 23060 24860 23112
rect 24912 23100 24918 23112
rect 26252 23109 26280 23140
rect 26973 23137 26985 23171
rect 27019 23137 27031 23171
rect 28258 23168 28264 23180
rect 28219 23140 28264 23168
rect 26973 23131 27031 23137
rect 28258 23128 28264 23140
rect 28316 23128 28322 23180
rect 29270 23128 29276 23180
rect 29328 23168 29334 23180
rect 29917 23171 29975 23177
rect 29917 23168 29929 23171
rect 29328 23140 29929 23168
rect 29328 23128 29334 23140
rect 29917 23137 29929 23140
rect 29963 23137 29975 23171
rect 29917 23131 29975 23137
rect 25593 23103 25651 23109
rect 25593 23100 25605 23103
rect 24912 23072 25605 23100
rect 24912 23060 24918 23072
rect 25593 23069 25605 23072
rect 25639 23069 25651 23103
rect 25593 23063 25651 23069
rect 26237 23103 26295 23109
rect 26237 23069 26249 23103
rect 26283 23069 26295 23103
rect 27154 23100 27160 23112
rect 27115 23072 27160 23100
rect 26237 23063 26295 23069
rect 19392 23004 20576 23032
rect 25608 23032 25636 23063
rect 27154 23060 27160 23072
rect 27212 23060 27218 23112
rect 28350 23060 28356 23112
rect 28408 23100 28414 23112
rect 28445 23103 28503 23109
rect 28445 23100 28457 23103
rect 28408 23072 28457 23100
rect 28408 23060 28414 23072
rect 28445 23069 28457 23072
rect 28491 23069 28503 23103
rect 28445 23063 28503 23069
rect 29733 23103 29791 23109
rect 29733 23069 29745 23103
rect 29779 23069 29791 23103
rect 30208 23100 30236 23276
rect 31205 23273 31217 23307
rect 31251 23304 31263 23307
rect 32490 23304 32496 23316
rect 31251 23276 32496 23304
rect 31251 23273 31263 23276
rect 31205 23267 31263 23273
rect 32490 23264 32496 23276
rect 32548 23264 32554 23316
rect 31386 23100 31392 23112
rect 30208 23072 31392 23100
rect 29733 23063 29791 23069
rect 26418 23032 26424 23044
rect 25608 23004 26424 23032
rect 19392 22992 19398 23004
rect 26418 22992 26424 23004
rect 26476 22992 26482 23044
rect 29748 23032 29776 23063
rect 31386 23060 31392 23072
rect 31444 23060 31450 23112
rect 34885 23103 34943 23109
rect 34885 23069 34897 23103
rect 34931 23100 34943 23103
rect 36998 23100 37004 23112
rect 34931 23072 37004 23100
rect 34931 23069 34943 23072
rect 34885 23063 34943 23069
rect 36998 23060 37004 23072
rect 37056 23060 37062 23112
rect 31846 23032 31852 23044
rect 29748 23004 31852 23032
rect 31846 22992 31852 23004
rect 31904 22992 31910 23044
rect 19426 22964 19432 22976
rect 17328 22936 19432 22964
rect 11388 22924 11394 22936
rect 19426 22924 19432 22936
rect 19484 22924 19490 22976
rect 19705 22967 19763 22973
rect 19705 22933 19717 22967
rect 19751 22964 19763 22967
rect 20070 22964 20076 22976
rect 19751 22936 20076 22964
rect 19751 22933 19763 22936
rect 19705 22927 19763 22933
rect 20070 22924 20076 22936
rect 20128 22924 20134 22976
rect 21637 22967 21695 22973
rect 21637 22933 21649 22967
rect 21683 22964 21695 22967
rect 22094 22964 22100 22976
rect 21683 22936 22100 22964
rect 21683 22933 21695 22936
rect 21637 22927 21695 22933
rect 22094 22924 22100 22936
rect 22152 22924 22158 22976
rect 25866 22924 25872 22976
rect 25924 22964 25930 22976
rect 26053 22967 26111 22973
rect 26053 22964 26065 22967
rect 25924 22936 26065 22964
rect 25924 22924 25930 22936
rect 26053 22933 26065 22936
rect 26099 22933 26111 22967
rect 26053 22927 26111 22933
rect 27617 22967 27675 22973
rect 27617 22933 27629 22967
rect 27663 22964 27675 22967
rect 28258 22964 28264 22976
rect 27663 22936 28264 22964
rect 27663 22933 27675 22936
rect 27617 22927 27675 22933
rect 28258 22924 28264 22936
rect 28316 22924 28322 22976
rect 30558 22924 30564 22976
rect 30616 22964 30622 22976
rect 34977 22967 35035 22973
rect 34977 22964 34989 22967
rect 30616 22936 34989 22964
rect 30616 22924 30622 22936
rect 34977 22933 34989 22936
rect 35023 22933 35035 22967
rect 34977 22927 35035 22933
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 15010 22720 15016 22772
rect 15068 22760 15074 22772
rect 15105 22763 15163 22769
rect 15105 22760 15117 22763
rect 15068 22732 15117 22760
rect 15068 22720 15074 22732
rect 15105 22729 15117 22732
rect 15151 22729 15163 22763
rect 15105 22723 15163 22729
rect 16209 22763 16267 22769
rect 16209 22729 16221 22763
rect 16255 22760 16267 22763
rect 17034 22760 17040 22772
rect 16255 22732 17040 22760
rect 16255 22729 16267 22732
rect 16209 22723 16267 22729
rect 17034 22720 17040 22732
rect 17092 22720 17098 22772
rect 18506 22720 18512 22772
rect 18564 22760 18570 22772
rect 19797 22763 19855 22769
rect 18564 22732 19748 22760
rect 18564 22720 18570 22732
rect 5350 22692 5356 22704
rect 5311 22664 5356 22692
rect 5350 22652 5356 22664
rect 5408 22652 5414 22704
rect 5445 22695 5503 22701
rect 5445 22661 5457 22695
rect 5491 22692 5503 22695
rect 5718 22692 5724 22704
rect 5491 22664 5724 22692
rect 5491 22661 5503 22664
rect 5445 22655 5503 22661
rect 5718 22652 5724 22664
rect 5776 22652 5782 22704
rect 8846 22692 8852 22704
rect 8807 22664 8852 22692
rect 8846 22652 8852 22664
rect 8904 22652 8910 22704
rect 9398 22692 9404 22704
rect 9359 22664 9404 22692
rect 9398 22652 9404 22664
rect 9456 22652 9462 22704
rect 11882 22692 11888 22704
rect 11843 22664 11888 22692
rect 11882 22652 11888 22664
rect 11940 22652 11946 22704
rect 14182 22692 14188 22704
rect 13464 22664 14188 22692
rect 1762 22624 1768 22636
rect 1723 22596 1768 22624
rect 1762 22584 1768 22596
rect 1820 22584 1826 22636
rect 3142 22624 3148 22636
rect 3103 22596 3148 22624
rect 3142 22584 3148 22596
rect 3200 22584 3206 22636
rect 13464 22633 13492 22664
rect 14182 22652 14188 22664
rect 14240 22692 14246 22704
rect 19720 22692 19748 22732
rect 19797 22729 19809 22763
rect 19843 22760 19855 22763
rect 19978 22760 19984 22772
rect 19843 22732 19984 22760
rect 19843 22729 19855 22732
rect 19797 22723 19855 22729
rect 19978 22720 19984 22732
rect 20036 22720 20042 22772
rect 21266 22760 21272 22772
rect 21227 22732 21272 22760
rect 21266 22720 21272 22732
rect 21324 22720 21330 22772
rect 27801 22763 27859 22769
rect 22066 22732 23428 22760
rect 22066 22692 22094 22732
rect 22370 22692 22376 22704
rect 14240 22664 18920 22692
rect 19720 22664 22094 22692
rect 22331 22664 22376 22692
rect 14240 22652 14246 22664
rect 13449 22627 13507 22633
rect 13449 22593 13461 22627
rect 13495 22593 13507 22627
rect 13449 22587 13507 22593
rect 15289 22627 15347 22633
rect 15289 22593 15301 22627
rect 15335 22624 15347 22627
rect 15654 22624 15660 22636
rect 15335 22596 15660 22624
rect 15335 22593 15347 22596
rect 15289 22587 15347 22593
rect 15654 22584 15660 22596
rect 15712 22584 15718 22636
rect 16114 22624 16120 22636
rect 16075 22596 16120 22624
rect 16114 22584 16120 22596
rect 16172 22624 16178 22636
rect 16850 22624 16856 22636
rect 16172 22596 16856 22624
rect 16172 22584 16178 22596
rect 16850 22584 16856 22596
rect 16908 22584 16914 22636
rect 17129 22627 17187 22633
rect 17129 22593 17141 22627
rect 17175 22624 17187 22627
rect 17770 22624 17776 22636
rect 17175 22596 17776 22624
rect 17175 22593 17187 22596
rect 17129 22587 17187 22593
rect 17770 22584 17776 22596
rect 17828 22584 17834 22636
rect 18892 22633 18920 22664
rect 22370 22652 22376 22664
rect 22428 22652 22434 22704
rect 18233 22627 18291 22633
rect 18233 22593 18245 22627
rect 18279 22624 18291 22627
rect 18877 22627 18935 22633
rect 18279 22596 18736 22624
rect 18279 22593 18291 22596
rect 18233 22587 18291 22593
rect 5994 22516 6000 22568
rect 6052 22556 6058 22568
rect 8757 22559 8815 22565
rect 8757 22556 8769 22559
rect 6052 22528 8769 22556
rect 6052 22516 6058 22528
rect 8757 22525 8769 22528
rect 8803 22525 8815 22559
rect 8757 22519 8815 22525
rect 10134 22516 10140 22568
rect 10192 22556 10198 22568
rect 10229 22559 10287 22565
rect 10229 22556 10241 22559
rect 10192 22528 10241 22556
rect 10192 22516 10198 22528
rect 10229 22525 10241 22528
rect 10275 22525 10287 22559
rect 11790 22556 11796 22568
rect 11751 22528 11796 22556
rect 10229 22519 10287 22525
rect 11790 22516 11796 22528
rect 11848 22516 11854 22568
rect 11974 22516 11980 22568
rect 12032 22556 12038 22568
rect 12069 22559 12127 22565
rect 12069 22556 12081 22559
rect 12032 22528 12081 22556
rect 12032 22516 12038 22528
rect 12069 22525 12081 22528
rect 12115 22556 12127 22559
rect 12250 22556 12256 22568
rect 12115 22528 12256 22556
rect 12115 22525 12127 22528
rect 12069 22519 12127 22525
rect 12250 22516 12256 22528
rect 12308 22516 12314 22568
rect 1581 22491 1639 22497
rect 1581 22457 1593 22491
rect 1627 22488 1639 22491
rect 5810 22488 5816 22500
rect 1627 22460 5816 22488
rect 1627 22457 1639 22460
rect 1581 22451 1639 22457
rect 5810 22448 5816 22460
rect 5868 22448 5874 22500
rect 5905 22491 5963 22497
rect 5905 22457 5917 22491
rect 5951 22488 5963 22491
rect 8110 22488 8116 22500
rect 5951 22460 8116 22488
rect 5951 22457 5963 22460
rect 5905 22451 5963 22457
rect 8110 22448 8116 22460
rect 8168 22448 8174 22500
rect 16942 22488 16948 22500
rect 16903 22460 16948 22488
rect 16942 22448 16948 22460
rect 17000 22448 17006 22500
rect 18708 22497 18736 22596
rect 18877 22593 18889 22627
rect 18923 22593 18935 22627
rect 18877 22587 18935 22593
rect 19150 22584 19156 22636
rect 19208 22624 19214 22636
rect 19981 22627 20039 22633
rect 19981 22624 19993 22627
rect 19208 22596 19993 22624
rect 19208 22584 19214 22596
rect 19981 22593 19993 22596
rect 20027 22624 20039 22627
rect 20714 22624 20720 22636
rect 20027 22596 20720 22624
rect 20027 22593 20039 22596
rect 19981 22587 20039 22593
rect 20714 22584 20720 22596
rect 20772 22584 20778 22636
rect 20990 22584 20996 22636
rect 21048 22624 21054 22636
rect 21453 22627 21511 22633
rect 21453 22624 21465 22627
rect 21048 22596 21465 22624
rect 21048 22584 21054 22596
rect 21453 22593 21465 22596
rect 21499 22593 21511 22627
rect 21453 22587 21511 22593
rect 22002 22516 22008 22568
rect 22060 22556 22066 22568
rect 22281 22559 22339 22565
rect 22281 22556 22293 22559
rect 22060 22528 22293 22556
rect 22060 22516 22066 22528
rect 22281 22525 22293 22528
rect 22327 22525 22339 22559
rect 22554 22556 22560 22568
rect 22515 22528 22560 22556
rect 22281 22519 22339 22525
rect 22554 22516 22560 22528
rect 22612 22516 22618 22568
rect 18693 22491 18751 22497
rect 18693 22457 18705 22491
rect 18739 22457 18751 22491
rect 18693 22451 18751 22457
rect 3234 22420 3240 22432
rect 3195 22392 3240 22420
rect 3234 22380 3240 22392
rect 3292 22380 3298 22432
rect 13262 22420 13268 22432
rect 13223 22392 13268 22420
rect 13262 22380 13268 22392
rect 13320 22380 13326 22432
rect 17954 22380 17960 22432
rect 18012 22420 18018 22432
rect 18049 22423 18107 22429
rect 18049 22420 18061 22423
rect 18012 22392 18061 22420
rect 18012 22380 18018 22392
rect 18049 22389 18061 22392
rect 18095 22389 18107 22423
rect 23400 22420 23428 22732
rect 27801 22729 27813 22763
rect 27847 22760 27859 22763
rect 28350 22760 28356 22772
rect 27847 22732 28356 22760
rect 27847 22729 27859 22732
rect 27801 22723 27859 22729
rect 28350 22720 28356 22732
rect 28408 22720 28414 22772
rect 23658 22692 23664 22704
rect 23619 22664 23664 22692
rect 23658 22652 23664 22664
rect 23716 22652 23722 22704
rect 24210 22692 24216 22704
rect 24171 22664 24216 22692
rect 24210 22652 24216 22664
rect 24268 22652 24274 22704
rect 25866 22692 25872 22704
rect 25827 22664 25872 22692
rect 25866 22652 25872 22664
rect 25924 22652 25930 22704
rect 26421 22695 26479 22701
rect 26421 22661 26433 22695
rect 26467 22692 26479 22695
rect 27614 22692 27620 22704
rect 26467 22664 27620 22692
rect 26467 22661 26479 22664
rect 26421 22655 26479 22661
rect 27614 22652 27620 22664
rect 27672 22692 27678 22704
rect 27890 22692 27896 22704
rect 27672 22664 27896 22692
rect 27672 22652 27678 22664
rect 27890 22652 27896 22664
rect 27948 22652 27954 22704
rect 27341 22627 27399 22633
rect 27341 22593 27353 22627
rect 27387 22624 27399 22627
rect 27430 22624 27436 22636
rect 27387 22596 27436 22624
rect 27387 22593 27399 22596
rect 27341 22587 27399 22593
rect 27430 22584 27436 22596
rect 27488 22584 27494 22636
rect 27985 22627 28043 22633
rect 27985 22593 27997 22627
rect 28031 22593 28043 22627
rect 28442 22624 28448 22636
rect 28403 22596 28448 22624
rect 27985 22587 28043 22593
rect 23569 22559 23627 22565
rect 23569 22525 23581 22559
rect 23615 22556 23627 22559
rect 25498 22556 25504 22568
rect 23615 22528 25504 22556
rect 23615 22525 23627 22528
rect 23569 22519 23627 22525
rect 25498 22516 25504 22528
rect 25556 22516 25562 22568
rect 25774 22556 25780 22568
rect 25735 22528 25780 22556
rect 25774 22516 25780 22528
rect 25832 22516 25838 22568
rect 28000 22556 28028 22587
rect 28442 22584 28448 22596
rect 28500 22584 28506 22636
rect 30469 22627 30527 22633
rect 30469 22593 30481 22627
rect 30515 22624 30527 22627
rect 32122 22624 32128 22636
rect 30515 22596 32128 22624
rect 30515 22593 30527 22596
rect 30469 22587 30527 22593
rect 32122 22584 32128 22596
rect 32180 22584 32186 22636
rect 28626 22556 28632 22568
rect 27172 22528 28028 22556
rect 28587 22528 28632 22556
rect 27172 22497 27200 22528
rect 28626 22516 28632 22528
rect 28684 22516 28690 22568
rect 30650 22556 30656 22568
rect 30611 22528 30656 22556
rect 30650 22516 30656 22528
rect 30708 22516 30714 22568
rect 27157 22491 27215 22497
rect 27157 22457 27169 22491
rect 27203 22457 27215 22491
rect 31110 22488 31116 22500
rect 27157 22451 27215 22457
rect 27264 22460 31116 22488
rect 27264 22420 27292 22460
rect 31110 22448 31116 22460
rect 31168 22448 31174 22500
rect 28994 22420 29000 22432
rect 23400 22392 27292 22420
rect 28955 22392 29000 22420
rect 18049 22383 18107 22389
rect 28994 22380 29000 22392
rect 29052 22380 29058 22432
rect 30374 22380 30380 22432
rect 30432 22420 30438 22432
rect 30837 22423 30895 22429
rect 30837 22420 30849 22423
rect 30432 22392 30849 22420
rect 30432 22380 30438 22392
rect 30837 22389 30849 22392
rect 30883 22389 30895 22423
rect 30837 22383 30895 22389
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 8846 22176 8852 22228
rect 8904 22216 8910 22228
rect 9217 22219 9275 22225
rect 9217 22216 9229 22219
rect 8904 22188 9229 22216
rect 8904 22176 8910 22188
rect 9217 22185 9229 22188
rect 9263 22185 9275 22219
rect 9217 22179 9275 22185
rect 16022 22176 16028 22228
rect 16080 22216 16086 22228
rect 16209 22219 16267 22225
rect 16209 22216 16221 22219
rect 16080 22188 16221 22216
rect 16080 22176 16086 22188
rect 16209 22185 16221 22188
rect 16255 22185 16267 22219
rect 16209 22179 16267 22185
rect 26605 22219 26663 22225
rect 26605 22185 26617 22219
rect 26651 22216 26663 22219
rect 27154 22216 27160 22228
rect 26651 22188 27160 22216
rect 26651 22185 26663 22188
rect 26605 22179 26663 22185
rect 27154 22176 27160 22188
rect 27212 22176 27218 22228
rect 28626 22176 28632 22228
rect 28684 22216 28690 22228
rect 28813 22219 28871 22225
rect 28813 22216 28825 22219
rect 28684 22188 28825 22216
rect 28684 22176 28690 22188
rect 28813 22185 28825 22188
rect 28859 22185 28871 22219
rect 30374 22216 30380 22228
rect 30335 22188 30380 22216
rect 28813 22179 28871 22185
rect 30374 22176 30380 22188
rect 30432 22176 30438 22228
rect 30650 22176 30656 22228
rect 30708 22216 30714 22228
rect 30837 22219 30895 22225
rect 30837 22216 30849 22219
rect 30708 22188 30849 22216
rect 30708 22176 30714 22188
rect 30837 22185 30849 22188
rect 30883 22185 30895 22219
rect 30837 22179 30895 22185
rect 5258 22108 5264 22160
rect 5316 22148 5322 22160
rect 16114 22148 16120 22160
rect 5316 22120 16120 22148
rect 5316 22108 5322 22120
rect 16114 22108 16120 22120
rect 16172 22108 16178 22160
rect 17770 22108 17776 22160
rect 17828 22148 17834 22160
rect 17828 22120 18000 22148
rect 17828 22108 17834 22120
rect 6362 22080 6368 22092
rect 6323 22052 6368 22080
rect 6362 22040 6368 22052
rect 6420 22040 6426 22092
rect 7009 22083 7067 22089
rect 7009 22049 7021 22083
rect 7055 22080 7067 22083
rect 9950 22080 9956 22092
rect 7055 22052 9956 22080
rect 7055 22049 7067 22052
rect 7009 22043 7067 22049
rect 9950 22040 9956 22052
rect 10008 22040 10014 22092
rect 10134 22080 10140 22092
rect 10095 22052 10140 22080
rect 10134 22040 10140 22052
rect 10192 22040 10198 22092
rect 11517 22083 11575 22089
rect 11517 22049 11529 22083
rect 11563 22080 11575 22083
rect 11790 22080 11796 22092
rect 11563 22052 11796 22080
rect 11563 22049 11575 22052
rect 11517 22043 11575 22049
rect 11790 22040 11796 22052
rect 11848 22040 11854 22092
rect 13078 22080 13084 22092
rect 12991 22052 13084 22080
rect 13078 22040 13084 22052
rect 13136 22080 13142 22092
rect 17405 22083 17463 22089
rect 13136 22052 16160 22080
rect 13136 22040 13142 22052
rect 5810 21972 5816 22024
rect 5868 22012 5874 22024
rect 6273 22015 6331 22021
rect 6273 22012 6285 22015
rect 5868 21984 6285 22012
rect 5868 21972 5874 21984
rect 6273 21981 6285 21984
rect 6319 21981 6331 22015
rect 6273 21975 6331 21981
rect 8481 22015 8539 22021
rect 8481 21981 8493 22015
rect 8527 22012 8539 22015
rect 8662 22012 8668 22024
rect 8527 21984 8668 22012
rect 8527 21981 8539 21984
rect 8481 21975 8539 21981
rect 8662 21972 8668 21984
rect 8720 21972 8726 22024
rect 9125 22015 9183 22021
rect 9125 21981 9137 22015
rect 9171 21981 9183 22015
rect 9125 21975 9183 21981
rect 10321 22015 10379 22021
rect 10321 21981 10333 22015
rect 10367 22012 10379 22015
rect 10870 22012 10876 22024
rect 10367 21984 10876 22012
rect 10367 21981 10379 21984
rect 10321 21975 10379 21981
rect 7098 21904 7104 21956
rect 7156 21944 7162 21956
rect 7156 21916 7201 21944
rect 7156 21904 7162 21916
rect 7282 21904 7288 21956
rect 7340 21944 7346 21956
rect 7653 21947 7711 21953
rect 7653 21944 7665 21947
rect 7340 21916 7665 21944
rect 7340 21904 7346 21916
rect 7653 21913 7665 21916
rect 7699 21913 7711 21947
rect 9140 21944 9168 21975
rect 10870 21972 10876 21984
rect 10928 21972 10934 22024
rect 13096 22012 13124 22040
rect 13262 22012 13268 22024
rect 11164 21984 13124 22012
rect 13223 21984 13268 22012
rect 11164 21944 11192 21984
rect 13262 21972 13268 21984
rect 13320 21972 13326 22024
rect 16132 22021 16160 22052
rect 17405 22049 17417 22083
rect 17451 22080 17463 22083
rect 17862 22080 17868 22092
rect 17451 22052 17868 22080
rect 17451 22049 17463 22052
rect 17405 22043 17463 22049
rect 17862 22040 17868 22052
rect 17920 22040 17926 22092
rect 17972 22080 18000 22120
rect 21008 22120 22416 22148
rect 21008 22080 21036 22120
rect 17972 22052 21036 22080
rect 21082 22040 21088 22092
rect 21140 22080 21146 22092
rect 21818 22080 21824 22092
rect 21140 22052 21824 22080
rect 21140 22040 21146 22052
rect 21818 22040 21824 22052
rect 21876 22080 21882 22092
rect 22281 22083 22339 22089
rect 22281 22080 22293 22083
rect 21876 22052 22293 22080
rect 21876 22040 21882 22052
rect 22281 22049 22293 22052
rect 22327 22049 22339 22083
rect 22388 22080 22416 22120
rect 23201 22083 23259 22089
rect 22388 22052 22876 22080
rect 22281 22043 22339 22049
rect 16117 22015 16175 22021
rect 16117 21981 16129 22015
rect 16163 21981 16175 22015
rect 16758 22012 16764 22024
rect 16719 21984 16764 22012
rect 16117 21975 16175 21981
rect 9140 21916 11192 21944
rect 16132 21944 16160 21975
rect 16758 21972 16764 21984
rect 16816 21972 16822 22024
rect 16942 22012 16948 22024
rect 16903 21984 16948 22012
rect 16942 21972 16948 21984
rect 17000 21972 17006 22024
rect 20441 22015 20499 22021
rect 20441 21981 20453 22015
rect 20487 22012 20499 22015
rect 20530 22012 20536 22024
rect 20487 21984 20536 22012
rect 20487 21981 20499 21984
rect 20441 21975 20499 21981
rect 20530 21972 20536 21984
rect 20588 21972 20594 22024
rect 20901 22015 20959 22021
rect 20901 21981 20913 22015
rect 20947 22012 20959 22015
rect 20990 22012 20996 22024
rect 20947 21984 20996 22012
rect 20947 21981 20959 21984
rect 20901 21975 20959 21981
rect 20990 21972 20996 21984
rect 21048 21972 21054 22024
rect 19334 21944 19340 21956
rect 16132 21916 19340 21944
rect 7653 21907 7711 21913
rect 19334 21904 19340 21916
rect 19392 21944 19398 21956
rect 19978 21944 19984 21956
rect 19392 21916 19984 21944
rect 19392 21904 19398 21916
rect 19978 21904 19984 21916
rect 20036 21904 20042 21956
rect 22002 21944 22008 21956
rect 21963 21916 22008 21944
rect 22002 21904 22008 21916
rect 22060 21904 22066 21956
rect 22094 21904 22100 21956
rect 22152 21944 22158 21956
rect 22848 21944 22876 22052
rect 23201 22049 23213 22083
rect 23247 22080 23259 22083
rect 23658 22080 23664 22092
rect 23247 22052 23664 22080
rect 23247 22049 23259 22052
rect 23201 22043 23259 22049
rect 23658 22040 23664 22052
rect 23716 22040 23722 22092
rect 24670 22080 24676 22092
rect 24631 22052 24676 22080
rect 24670 22040 24676 22052
rect 24728 22040 24734 22092
rect 25774 22040 25780 22092
rect 25832 22080 25838 22092
rect 25869 22083 25927 22089
rect 25869 22080 25881 22083
rect 25832 22052 25881 22080
rect 25832 22040 25838 22052
rect 25869 22049 25881 22052
rect 25915 22049 25927 22083
rect 29730 22080 29736 22092
rect 29691 22052 29736 22080
rect 25869 22043 25927 22049
rect 29730 22040 29736 22052
rect 29788 22040 29794 22092
rect 22922 21972 22928 22024
rect 22980 22012 22986 22024
rect 23109 22015 23167 22021
rect 23109 22012 23121 22015
rect 22980 21984 23121 22012
rect 22980 21972 22986 21984
rect 23109 21981 23121 21984
rect 23155 21981 23167 22015
rect 23109 21975 23167 21981
rect 24581 22015 24639 22021
rect 24581 21981 24593 22015
rect 24627 22012 24639 22015
rect 25682 22012 25688 22024
rect 24627 21984 25688 22012
rect 24627 21981 24639 21984
rect 24581 21975 24639 21981
rect 25682 21972 25688 21984
rect 25740 21972 25746 22024
rect 26418 21972 26424 22024
rect 26476 22012 26482 22024
rect 26513 22015 26571 22021
rect 26513 22012 26525 22015
rect 26476 21984 26525 22012
rect 26476 21972 26482 21984
rect 26513 21981 26525 21984
rect 26559 21981 26571 22015
rect 26513 21975 26571 21981
rect 27798 21972 27804 22024
rect 27856 22012 27862 22024
rect 28721 22015 28779 22021
rect 28721 22012 28733 22015
rect 27856 21984 28733 22012
rect 27856 21972 27862 21984
rect 28721 21981 28733 21984
rect 28767 21981 28779 22015
rect 28721 21975 28779 21981
rect 29270 21972 29276 22024
rect 29328 22012 29334 22024
rect 29917 22015 29975 22021
rect 29917 22012 29929 22015
rect 29328 21984 29929 22012
rect 29328 21972 29334 21984
rect 29917 21981 29929 21984
rect 29963 21981 29975 22015
rect 31018 22012 31024 22024
rect 30979 21984 31024 22012
rect 29917 21975 29975 21981
rect 31018 21972 31024 21984
rect 31076 21972 31082 22024
rect 37458 22012 37464 22024
rect 37419 21984 37464 22012
rect 37458 21972 37464 21984
rect 37516 21972 37522 22024
rect 37734 22012 37740 22024
rect 37695 21984 37740 22012
rect 37734 21972 37740 21984
rect 37792 21972 37798 22024
rect 29730 21944 29736 21956
rect 22152 21916 22197 21944
rect 22848 21916 29736 21944
rect 22152 21904 22158 21916
rect 29730 21904 29736 21916
rect 29788 21904 29794 21956
rect 8294 21876 8300 21888
rect 8255 21848 8300 21876
rect 8294 21836 8300 21848
rect 8352 21836 8358 21888
rect 9950 21836 9956 21888
rect 10008 21876 10014 21888
rect 10781 21879 10839 21885
rect 10781 21876 10793 21879
rect 10008 21848 10793 21876
rect 10008 21836 10014 21848
rect 10781 21845 10793 21848
rect 10827 21876 10839 21879
rect 12158 21876 12164 21888
rect 10827 21848 12164 21876
rect 10827 21845 10839 21848
rect 10781 21839 10839 21845
rect 12158 21836 12164 21848
rect 12216 21836 12222 21888
rect 13078 21876 13084 21888
rect 13039 21848 13084 21876
rect 13078 21836 13084 21848
rect 13136 21836 13142 21888
rect 20254 21876 20260 21888
rect 20215 21848 20260 21876
rect 20254 21836 20260 21848
rect 20312 21836 20318 21888
rect 20993 21879 21051 21885
rect 20993 21845 21005 21879
rect 21039 21876 21051 21879
rect 22186 21876 22192 21888
rect 21039 21848 22192 21876
rect 21039 21845 21051 21848
rect 20993 21839 21051 21845
rect 22186 21836 22192 21848
rect 22244 21836 22250 21888
rect 28074 21876 28080 21888
rect 28035 21848 28080 21876
rect 28074 21836 28080 21848
rect 28132 21836 28138 21888
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 7098 21672 7104 21684
rect 7059 21644 7104 21672
rect 7098 21632 7104 21644
rect 7156 21632 7162 21684
rect 8662 21672 8668 21684
rect 8623 21644 8668 21672
rect 8662 21632 8668 21644
rect 8720 21632 8726 21684
rect 10870 21672 10876 21684
rect 9600 21644 10272 21672
rect 10831 21644 10876 21672
rect 9600 21548 9628 21644
rect 9858 21604 9864 21616
rect 9819 21576 9864 21604
rect 9858 21564 9864 21576
rect 9916 21564 9922 21616
rect 10244 21604 10272 21644
rect 10870 21632 10876 21644
rect 10928 21632 10934 21684
rect 11882 21632 11888 21684
rect 11940 21672 11946 21684
rect 12069 21675 12127 21681
rect 12069 21672 12081 21675
rect 11940 21644 12081 21672
rect 11940 21632 11946 21644
rect 12069 21641 12081 21644
rect 12115 21641 12127 21675
rect 12069 21635 12127 21641
rect 12158 21632 12164 21684
rect 12216 21672 12222 21684
rect 13909 21675 13967 21681
rect 13909 21672 13921 21675
rect 12216 21644 13921 21672
rect 12216 21632 12222 21644
rect 13909 21641 13921 21644
rect 13955 21641 13967 21675
rect 13909 21635 13967 21641
rect 16206 21632 16212 21684
rect 16264 21672 16270 21684
rect 16264 21644 20760 21672
rect 16264 21632 16270 21644
rect 15930 21604 15936 21616
rect 10244 21576 15936 21604
rect 15930 21564 15936 21576
rect 15988 21564 15994 21616
rect 17954 21604 17960 21616
rect 17915 21576 17960 21604
rect 17954 21564 17960 21576
rect 18012 21564 18018 21616
rect 19889 21607 19947 21613
rect 19889 21573 19901 21607
rect 19935 21604 19947 21607
rect 20070 21604 20076 21616
rect 19935 21576 20076 21604
rect 19935 21573 19947 21576
rect 19889 21567 19947 21573
rect 20070 21564 20076 21576
rect 20128 21564 20134 21616
rect 20441 21607 20499 21613
rect 20441 21573 20453 21607
rect 20487 21604 20499 21607
rect 20622 21604 20628 21616
rect 20487 21576 20628 21604
rect 20487 21573 20499 21576
rect 20441 21567 20499 21573
rect 20622 21564 20628 21576
rect 20680 21564 20686 21616
rect 7006 21496 7012 21548
rect 7064 21536 7070 21548
rect 7285 21539 7343 21545
rect 7285 21536 7297 21539
rect 7064 21508 7297 21536
rect 7064 21496 7070 21508
rect 7285 21505 7297 21508
rect 7331 21505 7343 21539
rect 7285 21499 7343 21505
rect 8849 21539 8907 21545
rect 8849 21505 8861 21539
rect 8895 21536 8907 21539
rect 9582 21536 9588 21548
rect 8895 21508 9588 21536
rect 8895 21505 8907 21508
rect 8849 21499 8907 21505
rect 9582 21496 9588 21508
rect 9640 21496 9646 21548
rect 11054 21536 11060 21548
rect 11015 21508 11060 21536
rect 11054 21496 11060 21508
rect 11112 21496 11118 21548
rect 12250 21536 12256 21548
rect 12211 21508 12256 21536
rect 12250 21496 12256 21508
rect 12308 21496 12314 21548
rect 15102 21496 15108 21548
rect 15160 21536 15166 21548
rect 17586 21536 17592 21548
rect 15160 21508 17592 21536
rect 15160 21496 15166 21508
rect 17586 21496 17592 21508
rect 17644 21496 17650 21548
rect 7926 21468 7932 21480
rect 7887 21440 7932 21468
rect 7926 21428 7932 21440
rect 7984 21428 7990 21480
rect 9769 21471 9827 21477
rect 9769 21437 9781 21471
rect 9815 21468 9827 21471
rect 11146 21468 11152 21480
rect 9815 21440 11152 21468
rect 9815 21437 9827 21440
rect 9769 21431 9827 21437
rect 11146 21428 11152 21440
rect 11204 21428 11210 21480
rect 13265 21471 13323 21477
rect 13265 21437 13277 21471
rect 13311 21437 13323 21471
rect 13446 21468 13452 21480
rect 13407 21440 13452 21468
rect 13265 21431 13323 21437
rect 8662 21360 8668 21412
rect 8720 21400 8726 21412
rect 10321 21403 10379 21409
rect 10321 21400 10333 21403
rect 8720 21372 10333 21400
rect 8720 21360 8726 21372
rect 10321 21369 10333 21372
rect 10367 21369 10379 21403
rect 10321 21363 10379 21369
rect 13280 21332 13308 21431
rect 13446 21428 13452 21440
rect 13504 21428 13510 21480
rect 17862 21468 17868 21480
rect 17823 21440 17868 21468
rect 17862 21428 17868 21440
rect 17920 21428 17926 21480
rect 18141 21471 18199 21477
rect 18141 21437 18153 21471
rect 18187 21437 18199 21471
rect 19794 21468 19800 21480
rect 19755 21440 19800 21468
rect 18141 21431 18199 21437
rect 15102 21360 15108 21412
rect 15160 21400 15166 21412
rect 18156 21400 18184 21431
rect 19794 21428 19800 21440
rect 19852 21428 19858 21480
rect 15160 21372 18184 21400
rect 15160 21360 15166 21372
rect 19794 21332 19800 21344
rect 13280 21304 19800 21332
rect 19794 21292 19800 21304
rect 19852 21292 19858 21344
rect 20346 21292 20352 21344
rect 20404 21332 20410 21344
rect 20530 21332 20536 21344
rect 20404 21304 20536 21332
rect 20404 21292 20410 21304
rect 20530 21292 20536 21304
rect 20588 21292 20594 21344
rect 20732 21332 20760 21644
rect 22002 21632 22008 21684
rect 22060 21672 22066 21684
rect 28721 21675 28779 21681
rect 28721 21672 28733 21675
rect 22060 21644 28733 21672
rect 22060 21632 22066 21644
rect 28721 21641 28733 21644
rect 28767 21672 28779 21675
rect 28994 21672 29000 21684
rect 28767 21644 29000 21672
rect 28767 21641 28779 21644
rect 28721 21635 28779 21641
rect 28994 21632 29000 21644
rect 29052 21632 29058 21684
rect 29270 21672 29276 21684
rect 29231 21644 29276 21672
rect 29270 21632 29276 21644
rect 29328 21632 29334 21684
rect 29825 21675 29883 21681
rect 29825 21641 29837 21675
rect 29871 21672 29883 21675
rect 31018 21672 31024 21684
rect 29871 21644 31024 21672
rect 29871 21641 29883 21644
rect 29825 21635 29883 21641
rect 31018 21632 31024 21644
rect 31076 21632 31082 21684
rect 22186 21604 22192 21616
rect 22147 21576 22192 21604
rect 22186 21564 22192 21576
rect 22244 21564 22250 21616
rect 28074 21536 28080 21548
rect 28035 21508 28080 21536
rect 28074 21496 28080 21508
rect 28132 21496 28138 21548
rect 29178 21536 29184 21548
rect 29139 21508 29184 21536
rect 29178 21496 29184 21508
rect 29236 21536 29242 21548
rect 30009 21539 30067 21545
rect 30009 21536 30021 21539
rect 29236 21508 30021 21536
rect 29236 21496 29242 21508
rect 30009 21505 30021 21508
rect 30055 21505 30067 21539
rect 30009 21499 30067 21505
rect 22094 21428 22100 21480
rect 22152 21468 22158 21480
rect 22373 21471 22431 21477
rect 22152 21440 22197 21468
rect 22152 21428 22158 21440
rect 22373 21437 22385 21471
rect 22419 21437 22431 21471
rect 28258 21468 28264 21480
rect 28219 21440 28264 21468
rect 22373 21431 22431 21437
rect 21818 21360 21824 21412
rect 21876 21400 21882 21412
rect 22388 21400 22416 21431
rect 28258 21428 28264 21440
rect 28316 21428 28322 21480
rect 21876 21372 22416 21400
rect 21876 21360 21882 21372
rect 25682 21332 25688 21344
rect 20732 21304 25688 21332
rect 25682 21292 25688 21304
rect 25740 21292 25746 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 4985 21131 5043 21137
rect 4985 21097 4997 21131
rect 5031 21128 5043 21131
rect 5994 21128 6000 21140
rect 5031 21100 6000 21128
rect 5031 21097 5043 21100
rect 4985 21091 5043 21097
rect 5994 21088 6000 21100
rect 6052 21088 6058 21140
rect 7006 21128 7012 21140
rect 6967 21100 7012 21128
rect 7006 21088 7012 21100
rect 7064 21088 7070 21140
rect 9214 21128 9220 21140
rect 9175 21100 9220 21128
rect 9214 21088 9220 21100
rect 9272 21088 9278 21140
rect 9858 21128 9864 21140
rect 9819 21100 9864 21128
rect 9858 21088 9864 21100
rect 9916 21088 9922 21140
rect 13081 21131 13139 21137
rect 13081 21097 13093 21131
rect 13127 21128 13139 21131
rect 16942 21128 16948 21140
rect 13127 21100 16948 21128
rect 13127 21097 13139 21100
rect 13081 21091 13139 21097
rect 16942 21088 16948 21100
rect 17000 21088 17006 21140
rect 17862 21088 17868 21140
rect 17920 21128 17926 21140
rect 23474 21128 23480 21140
rect 17920 21100 23480 21128
rect 17920 21088 17926 21100
rect 23474 21088 23480 21100
rect 23532 21088 23538 21140
rect 28258 21128 28264 21140
rect 28219 21100 28264 21128
rect 28258 21088 28264 21100
rect 28316 21088 28322 21140
rect 15657 21063 15715 21069
rect 15657 21060 15669 21063
rect 12406 21032 15669 21060
rect 7926 20992 7932 21004
rect 7887 20964 7932 20992
rect 7926 20952 7932 20964
rect 7984 20952 7990 21004
rect 12406 20992 12434 21032
rect 15657 21029 15669 21032
rect 15703 21029 15715 21063
rect 15657 21023 15715 21029
rect 17586 21020 17592 21072
rect 17644 21060 17650 21072
rect 17957 21063 18015 21069
rect 17957 21060 17969 21063
rect 17644 21032 17969 21060
rect 17644 21020 17650 21032
rect 17957 21029 17969 21032
rect 18003 21029 18015 21063
rect 17957 21023 18015 21029
rect 27617 21063 27675 21069
rect 27617 21029 27629 21063
rect 27663 21029 27675 21063
rect 27617 21023 27675 21029
rect 9140 20964 12434 20992
rect 15105 20995 15163 21001
rect 1762 20924 1768 20936
rect 1723 20896 1768 20924
rect 1762 20884 1768 20896
rect 1820 20884 1826 20936
rect 3786 20884 3792 20936
rect 3844 20924 3850 20936
rect 4893 20927 4951 20933
rect 4893 20924 4905 20927
rect 3844 20896 4905 20924
rect 3844 20884 3850 20896
rect 4893 20893 4905 20896
rect 4939 20893 4951 20927
rect 4893 20887 4951 20893
rect 7193 20927 7251 20933
rect 7193 20893 7205 20927
rect 7239 20924 7251 20927
rect 7650 20924 7656 20936
rect 7239 20896 7656 20924
rect 7239 20893 7251 20896
rect 7193 20887 7251 20893
rect 7650 20884 7656 20896
rect 7708 20884 7714 20936
rect 9140 20933 9168 20964
rect 15105 20961 15117 20995
rect 15151 20992 15163 20995
rect 15151 20964 18644 20992
rect 15151 20961 15163 20964
rect 15105 20955 15163 20961
rect 8573 20927 8631 20933
rect 8573 20893 8585 20927
rect 8619 20924 8631 20927
rect 9125 20927 9183 20933
rect 9125 20924 9137 20927
rect 8619 20896 9137 20924
rect 8619 20893 8631 20896
rect 8573 20887 8631 20893
rect 9125 20893 9137 20896
rect 9171 20893 9183 20927
rect 10042 20924 10048 20936
rect 10003 20896 10048 20924
rect 9125 20887 9183 20893
rect 10042 20884 10048 20896
rect 10100 20884 10106 20936
rect 12434 20884 12440 20936
rect 12492 20924 12498 20936
rect 12986 20924 12992 20936
rect 12492 20896 12992 20924
rect 12492 20884 12498 20896
rect 12986 20884 12992 20896
rect 13044 20884 13050 20936
rect 14550 20924 14556 20936
rect 14511 20896 14556 20924
rect 14550 20884 14556 20896
rect 14608 20924 14614 20936
rect 14918 20924 14924 20936
rect 14608 20896 14924 20924
rect 14608 20884 14614 20896
rect 14918 20884 14924 20896
rect 14976 20884 14982 20936
rect 8021 20859 8079 20865
rect 8021 20825 8033 20859
rect 8067 20856 8079 20859
rect 8294 20856 8300 20868
rect 8067 20828 8300 20856
rect 8067 20825 8079 20828
rect 8021 20819 8079 20825
rect 8294 20816 8300 20828
rect 8352 20816 8358 20868
rect 15102 20856 15108 20868
rect 12406 20828 15108 20856
rect 1581 20791 1639 20797
rect 1581 20757 1593 20791
rect 1627 20788 1639 20791
rect 5350 20788 5356 20800
rect 1627 20760 5356 20788
rect 1627 20757 1639 20760
rect 1581 20751 1639 20757
rect 5350 20748 5356 20760
rect 5408 20748 5414 20800
rect 8110 20748 8116 20800
rect 8168 20788 8174 20800
rect 12406 20788 12434 20828
rect 15102 20816 15108 20828
rect 15160 20816 15166 20868
rect 15194 20816 15200 20868
rect 15252 20856 15258 20868
rect 17402 20856 17408 20868
rect 15252 20828 15297 20856
rect 17363 20828 17408 20856
rect 15252 20816 15258 20828
rect 17402 20816 17408 20828
rect 17460 20816 17466 20868
rect 17497 20859 17555 20865
rect 17497 20825 17509 20859
rect 17543 20825 17555 20859
rect 18616 20856 18644 20964
rect 20622 20952 20628 21004
rect 20680 20992 20686 21004
rect 27632 20992 27660 21023
rect 20680 20964 26280 20992
rect 27632 20964 28488 20992
rect 20680 20952 20686 20964
rect 19426 20924 19432 20936
rect 19387 20896 19432 20924
rect 19426 20884 19432 20896
rect 19484 20884 19490 20936
rect 20254 20884 20260 20936
rect 20312 20924 20318 20936
rect 20809 20927 20867 20933
rect 20809 20924 20821 20927
rect 20312 20896 20821 20924
rect 20312 20884 20318 20896
rect 20809 20893 20821 20896
rect 20855 20893 20867 20927
rect 25590 20924 25596 20936
rect 25551 20896 25596 20924
rect 20809 20887 20867 20893
rect 25590 20884 25596 20896
rect 25648 20884 25654 20936
rect 26252 20924 26280 20964
rect 27798 20924 27804 20936
rect 26252 20896 27804 20924
rect 27798 20884 27804 20896
rect 27856 20884 27862 20936
rect 28460 20933 28488 20964
rect 28445 20927 28503 20933
rect 28445 20893 28457 20927
rect 28491 20893 28503 20927
rect 29730 20924 29736 20936
rect 29691 20896 29736 20924
rect 28445 20887 28503 20893
rect 29730 20884 29736 20896
rect 29788 20884 29794 20936
rect 30374 20924 30380 20936
rect 30335 20896 30380 20924
rect 30374 20884 30380 20896
rect 30432 20884 30438 20936
rect 38286 20924 38292 20936
rect 38247 20896 38292 20924
rect 38286 20884 38292 20896
rect 38344 20884 38350 20936
rect 24762 20856 24768 20868
rect 18616 20828 24768 20856
rect 17497 20819 17555 20825
rect 8168 20760 12434 20788
rect 14369 20791 14427 20797
rect 8168 20748 8174 20760
rect 14369 20757 14381 20791
rect 14415 20788 14427 20791
rect 14642 20788 14648 20800
rect 14415 20760 14648 20788
rect 14415 20757 14427 20760
rect 14369 20751 14427 20757
rect 14642 20748 14648 20760
rect 14700 20748 14706 20800
rect 17512 20788 17540 20819
rect 24762 20816 24768 20828
rect 24820 20816 24826 20868
rect 19521 20791 19579 20797
rect 19521 20788 19533 20791
rect 17512 20760 19533 20788
rect 19521 20757 19533 20760
rect 19567 20757 19579 20791
rect 19521 20751 19579 20757
rect 19794 20748 19800 20800
rect 19852 20788 19858 20800
rect 20254 20788 20260 20800
rect 19852 20760 20260 20788
rect 19852 20748 19858 20760
rect 20254 20748 20260 20760
rect 20312 20748 20318 20800
rect 20346 20748 20352 20800
rect 20404 20788 20410 20800
rect 20625 20791 20683 20797
rect 20625 20788 20637 20791
rect 20404 20760 20637 20788
rect 20404 20748 20410 20760
rect 20625 20757 20637 20760
rect 20671 20757 20683 20791
rect 25406 20788 25412 20800
rect 25367 20760 25412 20788
rect 20625 20751 20683 20757
rect 25406 20748 25412 20760
rect 25464 20748 25470 20800
rect 28994 20748 29000 20800
rect 29052 20788 29058 20800
rect 29825 20791 29883 20797
rect 29825 20788 29837 20791
rect 29052 20760 29837 20788
rect 29052 20748 29058 20760
rect 29825 20757 29837 20760
rect 29871 20757 29883 20791
rect 29825 20751 29883 20757
rect 30469 20791 30527 20797
rect 30469 20757 30481 20791
rect 30515 20788 30527 20791
rect 31478 20788 31484 20800
rect 30515 20760 31484 20788
rect 30515 20757 30527 20760
rect 30469 20751 30527 20757
rect 31478 20748 31484 20760
rect 31536 20748 31542 20800
rect 34514 20748 34520 20800
rect 34572 20788 34578 20800
rect 38105 20791 38163 20797
rect 38105 20788 38117 20791
rect 34572 20760 38117 20788
rect 34572 20748 34578 20760
rect 38105 20757 38117 20760
rect 38151 20757 38163 20791
rect 38105 20751 38163 20757
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 5718 20544 5724 20596
rect 5776 20584 5782 20596
rect 5905 20587 5963 20593
rect 5905 20584 5917 20587
rect 5776 20556 5917 20584
rect 5776 20544 5782 20556
rect 5905 20553 5917 20556
rect 5951 20553 5963 20587
rect 5905 20547 5963 20553
rect 10965 20587 11023 20593
rect 10965 20553 10977 20587
rect 11011 20584 11023 20587
rect 11054 20584 11060 20596
rect 11011 20556 11060 20584
rect 11011 20553 11023 20556
rect 10965 20547 11023 20553
rect 11054 20544 11060 20556
rect 11112 20544 11118 20596
rect 19426 20544 19432 20596
rect 19484 20584 19490 20596
rect 21266 20584 21272 20596
rect 19484 20556 21272 20584
rect 19484 20544 19490 20556
rect 21266 20544 21272 20556
rect 21324 20544 21330 20596
rect 24949 20587 25007 20593
rect 24949 20553 24961 20587
rect 24995 20584 25007 20587
rect 25590 20584 25596 20596
rect 24995 20556 25596 20584
rect 24995 20553 25007 20556
rect 24949 20547 25007 20553
rect 25590 20544 25596 20556
rect 25648 20544 25654 20596
rect 30466 20584 30472 20596
rect 29104 20556 30472 20584
rect 8110 20516 8116 20528
rect 8071 20488 8116 20516
rect 8110 20476 8116 20488
rect 8168 20476 8174 20528
rect 8205 20519 8263 20525
rect 8205 20485 8217 20519
rect 8251 20516 8263 20519
rect 9766 20516 9772 20528
rect 8251 20488 9772 20516
rect 8251 20485 8263 20488
rect 8205 20479 8263 20485
rect 9766 20476 9772 20488
rect 9824 20476 9830 20528
rect 20438 20476 20444 20528
rect 20496 20516 20502 20528
rect 20806 20516 20812 20528
rect 20496 20488 20812 20516
rect 20496 20476 20502 20488
rect 20806 20476 20812 20488
rect 20864 20476 20870 20528
rect 23569 20519 23627 20525
rect 23569 20485 23581 20519
rect 23615 20516 23627 20519
rect 25406 20516 25412 20528
rect 23615 20488 25412 20516
rect 23615 20485 23627 20488
rect 23569 20479 23627 20485
rect 25406 20476 25412 20488
rect 25464 20476 25470 20528
rect 25608 20488 27384 20516
rect 2777 20451 2835 20457
rect 2777 20417 2789 20451
rect 2823 20448 2835 20451
rect 3234 20448 3240 20460
rect 2823 20420 3240 20448
rect 2823 20417 2835 20420
rect 2777 20411 2835 20417
rect 3234 20408 3240 20420
rect 3292 20408 3298 20460
rect 5810 20448 5816 20460
rect 5771 20420 5816 20448
rect 5810 20408 5816 20420
rect 5868 20408 5874 20460
rect 6549 20451 6607 20457
rect 6549 20417 6561 20451
rect 6595 20448 6607 20451
rect 7650 20448 7656 20460
rect 6595 20420 7656 20448
rect 6595 20417 6607 20420
rect 6549 20411 6607 20417
rect 7650 20408 7656 20420
rect 7708 20408 7714 20460
rect 11149 20451 11207 20457
rect 11149 20417 11161 20451
rect 11195 20448 11207 20451
rect 12342 20448 12348 20460
rect 11195 20420 12348 20448
rect 11195 20417 11207 20420
rect 11149 20411 11207 20417
rect 2961 20383 3019 20389
rect 2961 20349 2973 20383
rect 3007 20380 3019 20383
rect 4614 20380 4620 20392
rect 3007 20352 4620 20380
rect 3007 20349 3019 20352
rect 2961 20343 3019 20349
rect 4614 20340 4620 20352
rect 4672 20340 4678 20392
rect 5626 20340 5632 20392
rect 5684 20380 5690 20392
rect 11164 20380 11192 20411
rect 12342 20408 12348 20420
rect 12400 20408 12406 20460
rect 12713 20451 12771 20457
rect 12713 20417 12725 20451
rect 12759 20448 12771 20451
rect 13078 20448 13084 20460
rect 12759 20420 13084 20448
rect 12759 20417 12771 20420
rect 12713 20411 12771 20417
rect 13078 20408 13084 20420
rect 13136 20408 13142 20460
rect 14642 20448 14648 20460
rect 14603 20420 14648 20448
rect 14642 20408 14648 20420
rect 14700 20408 14706 20460
rect 15657 20451 15715 20457
rect 15657 20417 15669 20451
rect 15703 20448 15715 20451
rect 25130 20448 25136 20460
rect 15703 20420 22094 20448
rect 25091 20420 25136 20448
rect 15703 20417 15715 20420
rect 15657 20411 15715 20417
rect 5684 20352 11192 20380
rect 11885 20383 11943 20389
rect 5684 20340 5690 20352
rect 11885 20349 11897 20383
rect 11931 20380 11943 20383
rect 12529 20383 12587 20389
rect 12529 20380 12541 20383
rect 11931 20352 12541 20380
rect 11931 20349 11943 20352
rect 11885 20343 11943 20349
rect 12529 20349 12541 20352
rect 12575 20349 12587 20383
rect 15838 20380 15844 20392
rect 15799 20352 15844 20380
rect 12529 20343 12587 20349
rect 15838 20340 15844 20352
rect 15896 20340 15902 20392
rect 16482 20340 16488 20392
rect 16540 20380 16546 20392
rect 20809 20383 20867 20389
rect 20809 20380 20821 20383
rect 16540 20352 20821 20380
rect 16540 20340 16546 20352
rect 20809 20349 20821 20352
rect 20855 20349 20867 20383
rect 20809 20343 20867 20349
rect 20993 20383 21051 20389
rect 20993 20349 21005 20383
rect 21039 20380 21051 20383
rect 21358 20380 21364 20392
rect 21039 20352 21364 20380
rect 21039 20349 21051 20352
rect 20993 20343 21051 20349
rect 21358 20340 21364 20352
rect 21416 20340 21422 20392
rect 8662 20312 8668 20324
rect 8623 20284 8668 20312
rect 8662 20272 8668 20284
rect 8720 20272 8726 20324
rect 11146 20272 11152 20324
rect 11204 20312 11210 20324
rect 13173 20315 13231 20321
rect 13173 20312 13185 20315
rect 11204 20284 13185 20312
rect 11204 20272 11210 20284
rect 13173 20281 13185 20284
rect 13219 20312 13231 20315
rect 16025 20315 16083 20321
rect 16025 20312 16037 20315
rect 13219 20284 16037 20312
rect 13219 20281 13231 20284
rect 13173 20275 13231 20281
rect 16025 20281 16037 20284
rect 16071 20281 16083 20315
rect 22066 20312 22094 20420
rect 25130 20408 25136 20420
rect 25188 20408 25194 20460
rect 23474 20380 23480 20392
rect 23435 20352 23480 20380
rect 23474 20340 23480 20352
rect 23532 20340 23538 20392
rect 25608 20380 25636 20488
rect 25682 20408 25688 20460
rect 25740 20448 25746 20460
rect 27356 20457 27384 20488
rect 25869 20451 25927 20457
rect 25869 20448 25881 20451
rect 25740 20420 25881 20448
rect 25740 20408 25746 20420
rect 25869 20417 25881 20420
rect 25915 20417 25927 20451
rect 25869 20411 25927 20417
rect 26513 20451 26571 20457
rect 26513 20417 26525 20451
rect 26559 20417 26571 20451
rect 26513 20411 26571 20417
rect 27341 20451 27399 20457
rect 27341 20417 27353 20451
rect 27387 20448 27399 20451
rect 28166 20448 28172 20460
rect 27387 20420 28172 20448
rect 27387 20417 27399 20420
rect 27341 20411 27399 20417
rect 26528 20380 26556 20411
rect 28166 20408 28172 20420
rect 28224 20408 28230 20460
rect 28261 20451 28319 20457
rect 28261 20417 28273 20451
rect 28307 20448 28319 20451
rect 28994 20448 29000 20460
rect 28307 20420 29000 20448
rect 28307 20417 28319 20420
rect 28261 20411 28319 20417
rect 28994 20408 29000 20420
rect 29052 20408 29058 20460
rect 23860 20352 25636 20380
rect 25700 20352 26556 20380
rect 28077 20383 28135 20389
rect 22066 20284 22692 20312
rect 16025 20275 16083 20281
rect 3421 20247 3479 20253
rect 3421 20213 3433 20247
rect 3467 20244 3479 20247
rect 5074 20244 5080 20256
rect 3467 20216 5080 20244
rect 3467 20213 3479 20216
rect 3421 20207 3479 20213
rect 5074 20204 5080 20216
rect 5132 20204 5138 20256
rect 5166 20204 5172 20256
rect 5224 20244 5230 20256
rect 6641 20247 6699 20253
rect 6641 20244 6653 20247
rect 5224 20216 6653 20244
rect 5224 20204 5230 20216
rect 6641 20213 6653 20216
rect 6687 20213 6699 20247
rect 6641 20207 6699 20213
rect 9306 20204 9312 20256
rect 9364 20244 9370 20256
rect 14366 20244 14372 20256
rect 9364 20216 14372 20244
rect 9364 20204 9370 20216
rect 14366 20204 14372 20216
rect 14424 20204 14430 20256
rect 14461 20247 14519 20253
rect 14461 20213 14473 20247
rect 14507 20244 14519 20247
rect 15378 20244 15384 20256
rect 14507 20216 15384 20244
rect 14507 20213 14519 20216
rect 14461 20207 14519 20213
rect 15378 20204 15384 20216
rect 15436 20204 15442 20256
rect 21174 20244 21180 20256
rect 21135 20216 21180 20244
rect 21174 20204 21180 20216
rect 21232 20244 21238 20256
rect 22094 20244 22100 20256
rect 21232 20216 22100 20244
rect 21232 20204 21238 20216
rect 22094 20204 22100 20216
rect 22152 20204 22158 20256
rect 22664 20244 22692 20284
rect 22738 20272 22744 20324
rect 22796 20312 22802 20324
rect 23860 20312 23888 20352
rect 24026 20312 24032 20324
rect 22796 20284 23888 20312
rect 23987 20284 24032 20312
rect 22796 20272 22802 20284
rect 24026 20272 24032 20284
rect 24084 20272 24090 20324
rect 25700 20321 25728 20352
rect 28077 20349 28089 20383
rect 28123 20380 28135 20383
rect 29104 20380 29132 20556
rect 30466 20544 30472 20556
rect 30524 20544 30530 20596
rect 29362 20516 29368 20528
rect 29323 20488 29368 20516
rect 29362 20476 29368 20488
rect 29420 20476 29426 20528
rect 28123 20352 29132 20380
rect 29273 20383 29331 20389
rect 28123 20349 28135 20352
rect 28077 20343 28135 20349
rect 29273 20349 29285 20383
rect 29319 20380 29331 20383
rect 30742 20380 30748 20392
rect 29319 20352 30748 20380
rect 29319 20349 29331 20352
rect 29273 20343 29331 20349
rect 25685 20315 25743 20321
rect 25685 20281 25697 20315
rect 25731 20281 25743 20315
rect 28092 20312 28120 20343
rect 30742 20340 30748 20352
rect 30800 20340 30806 20392
rect 29822 20312 29828 20324
rect 25685 20275 25743 20281
rect 25792 20284 28120 20312
rect 29783 20284 29828 20312
rect 25792 20244 25820 20284
rect 29822 20272 29828 20284
rect 29880 20272 29886 20324
rect 22664 20216 25820 20244
rect 25866 20204 25872 20256
rect 25924 20244 25930 20256
rect 26329 20247 26387 20253
rect 26329 20244 26341 20247
rect 25924 20216 26341 20244
rect 25924 20204 25930 20216
rect 26329 20213 26341 20216
rect 26375 20213 26387 20247
rect 26329 20207 26387 20213
rect 27157 20247 27215 20253
rect 27157 20213 27169 20247
rect 27203 20244 27215 20247
rect 27338 20244 27344 20256
rect 27203 20216 27344 20244
rect 27203 20213 27215 20216
rect 27157 20207 27215 20213
rect 27338 20204 27344 20216
rect 27396 20204 27402 20256
rect 28721 20247 28779 20253
rect 28721 20213 28733 20247
rect 28767 20244 28779 20247
rect 30098 20244 30104 20256
rect 28767 20216 30104 20244
rect 28767 20213 28779 20216
rect 28721 20207 28779 20213
rect 30098 20204 30104 20216
rect 30156 20204 30162 20256
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 9769 20043 9827 20049
rect 9769 20009 9781 20043
rect 9815 20040 9827 20043
rect 10042 20040 10048 20052
rect 9815 20012 10048 20040
rect 9815 20009 9827 20012
rect 9769 20003 9827 20009
rect 10042 20000 10048 20012
rect 10100 20000 10106 20052
rect 12069 20043 12127 20049
rect 12069 20009 12081 20043
rect 12115 20040 12127 20043
rect 12250 20040 12256 20052
rect 12115 20012 12256 20040
rect 12115 20009 12127 20012
rect 12069 20003 12127 20009
rect 12250 20000 12256 20012
rect 12308 20000 12314 20052
rect 12805 20043 12863 20049
rect 12805 20009 12817 20043
rect 12851 20040 12863 20043
rect 13446 20040 13452 20052
rect 12851 20012 13452 20040
rect 12851 20009 12863 20012
rect 12805 20003 12863 20009
rect 13446 20000 13452 20012
rect 13504 20000 13510 20052
rect 15194 20000 15200 20052
rect 15252 20040 15258 20052
rect 15749 20043 15807 20049
rect 15749 20040 15761 20043
rect 15252 20012 15761 20040
rect 15252 20000 15258 20012
rect 15749 20009 15761 20012
rect 15795 20009 15807 20043
rect 15749 20003 15807 20009
rect 15930 20000 15936 20052
rect 15988 20040 15994 20052
rect 20070 20040 20076 20052
rect 15988 20012 20076 20040
rect 15988 20000 15994 20012
rect 20070 20000 20076 20012
rect 20128 20000 20134 20052
rect 21358 20040 21364 20052
rect 21319 20012 21364 20040
rect 21358 20000 21364 20012
rect 21416 20000 21422 20052
rect 28537 20043 28595 20049
rect 28537 20009 28549 20043
rect 28583 20040 28595 20043
rect 29362 20040 29368 20052
rect 28583 20012 29368 20040
rect 28583 20009 28595 20012
rect 28537 20003 28595 20009
rect 29362 20000 29368 20012
rect 29420 20000 29426 20052
rect 30742 20040 30748 20052
rect 30703 20012 30748 20040
rect 30742 20000 30748 20012
rect 30800 20000 30806 20052
rect 6086 19932 6092 19984
rect 6144 19972 6150 19984
rect 14090 19972 14096 19984
rect 6144 19944 14096 19972
rect 6144 19932 6150 19944
rect 14090 19932 14096 19944
rect 14148 19932 14154 19984
rect 14921 19975 14979 19981
rect 14921 19941 14933 19975
rect 14967 19972 14979 19975
rect 16574 19972 16580 19984
rect 14967 19944 16580 19972
rect 14967 19941 14979 19944
rect 14921 19935 14979 19941
rect 16574 19932 16580 19944
rect 16632 19932 16638 19984
rect 20162 19932 20168 19984
rect 20220 19972 20226 19984
rect 20220 19944 22876 19972
rect 20220 19932 20226 19944
rect 5074 19904 5080 19916
rect 5035 19876 5080 19904
rect 5074 19864 5080 19876
rect 5132 19864 5138 19916
rect 5721 19907 5779 19913
rect 5721 19873 5733 19907
rect 5767 19904 5779 19907
rect 7282 19904 7288 19916
rect 5767 19876 7288 19904
rect 5767 19873 5779 19876
rect 5721 19867 5779 19873
rect 7282 19864 7288 19876
rect 7340 19864 7346 19916
rect 11149 19907 11207 19913
rect 11149 19873 11161 19907
rect 11195 19904 11207 19907
rect 11974 19904 11980 19916
rect 11195 19876 11980 19904
rect 11195 19873 11207 19876
rect 11149 19867 11207 19873
rect 11974 19864 11980 19876
rect 12032 19864 12038 19916
rect 15010 19864 15016 19916
rect 15068 19904 15074 19916
rect 15068 19876 16528 19904
rect 15068 19864 15074 19876
rect 6181 19839 6239 19845
rect 6181 19805 6193 19839
rect 6227 19836 6239 19839
rect 9306 19836 9312 19848
rect 6227 19808 9312 19836
rect 6227 19805 6239 19808
rect 6181 19799 6239 19805
rect 9306 19796 9312 19808
rect 9364 19796 9370 19848
rect 9950 19836 9956 19848
rect 9911 19808 9956 19836
rect 9950 19796 9956 19808
rect 10008 19796 10014 19848
rect 12066 19796 12072 19848
rect 12124 19836 12130 19848
rect 12253 19839 12311 19845
rect 12253 19836 12265 19839
rect 12124 19808 12265 19836
rect 12124 19796 12130 19808
rect 12253 19805 12265 19808
rect 12299 19805 12311 19839
rect 12253 19799 12311 19805
rect 12342 19796 12348 19848
rect 12400 19836 12406 19848
rect 12713 19839 12771 19845
rect 12713 19836 12725 19839
rect 12400 19808 12725 19836
rect 12400 19796 12406 19808
rect 12713 19805 12725 19808
rect 12759 19805 12771 19839
rect 12713 19799 12771 19805
rect 14277 19839 14335 19845
rect 14277 19805 14289 19839
rect 14323 19805 14335 19839
rect 15102 19836 15108 19848
rect 15063 19808 15108 19836
rect 14277 19799 14335 19805
rect 5166 19728 5172 19780
rect 5224 19768 5230 19780
rect 10502 19768 10508 19780
rect 5224 19740 5269 19768
rect 10463 19740 10508 19768
rect 5224 19728 5230 19740
rect 10502 19728 10508 19740
rect 10560 19728 10566 19780
rect 10597 19771 10655 19777
rect 10597 19737 10609 19771
rect 10643 19768 10655 19771
rect 12158 19768 12164 19780
rect 10643 19740 12164 19768
rect 10643 19737 10655 19740
rect 10597 19731 10655 19737
rect 12158 19728 12164 19740
rect 12216 19728 12222 19780
rect 6273 19703 6331 19709
rect 6273 19669 6285 19703
rect 6319 19700 6331 19703
rect 7282 19700 7288 19712
rect 6319 19672 7288 19700
rect 6319 19669 6331 19672
rect 6273 19663 6331 19669
rect 7282 19660 7288 19672
rect 7340 19660 7346 19712
rect 14292 19700 14320 19799
rect 15102 19796 15108 19808
rect 15160 19796 15166 19848
rect 15657 19839 15715 19845
rect 15657 19805 15669 19839
rect 15703 19836 15715 19839
rect 15930 19836 15936 19848
rect 15703 19808 15936 19836
rect 15703 19805 15715 19808
rect 15657 19799 15715 19805
rect 15930 19796 15936 19808
rect 15988 19796 15994 19848
rect 16500 19845 16528 19876
rect 16758 19864 16764 19916
rect 16816 19904 16822 19916
rect 17129 19907 17187 19913
rect 17129 19904 17141 19907
rect 16816 19876 17141 19904
rect 16816 19864 16822 19876
rect 17129 19873 17141 19876
rect 17175 19904 17187 19907
rect 18322 19904 18328 19916
rect 17175 19876 18328 19904
rect 17175 19873 17187 19876
rect 17129 19867 17187 19873
rect 18322 19864 18328 19876
rect 18380 19864 18386 19916
rect 18874 19864 18880 19916
rect 18932 19904 18938 19916
rect 22738 19904 22744 19916
rect 18932 19876 22744 19904
rect 18932 19864 18938 19876
rect 22738 19864 22744 19876
rect 22796 19864 22802 19916
rect 22848 19913 22876 19944
rect 24762 19932 24768 19984
rect 24820 19972 24826 19984
rect 27433 19975 27491 19981
rect 27433 19972 27445 19975
rect 24820 19944 27445 19972
rect 24820 19932 24826 19944
rect 27433 19941 27445 19944
rect 27479 19972 27491 19975
rect 29822 19972 29828 19984
rect 27479 19944 29828 19972
rect 27479 19941 27491 19944
rect 27433 19935 27491 19941
rect 29822 19932 29828 19944
rect 29880 19932 29886 19984
rect 22833 19907 22891 19913
rect 22833 19873 22845 19907
rect 22879 19873 22891 19907
rect 26326 19904 26332 19916
rect 26287 19876 26332 19904
rect 22833 19867 22891 19873
rect 26326 19864 26332 19876
rect 26384 19864 26390 19916
rect 26881 19907 26939 19913
rect 26881 19873 26893 19907
rect 26927 19904 26939 19907
rect 27706 19904 27712 19916
rect 26927 19876 27712 19904
rect 26927 19873 26939 19876
rect 26881 19867 26939 19873
rect 27706 19864 27712 19876
rect 27764 19864 27770 19916
rect 30466 19904 30472 19916
rect 29564 19876 30472 19904
rect 16485 19839 16543 19845
rect 16485 19805 16497 19839
rect 16531 19805 16543 19839
rect 16485 19799 16543 19805
rect 19334 19796 19340 19848
rect 19392 19836 19398 19848
rect 20622 19836 20628 19848
rect 19392 19808 20628 19836
rect 19392 19796 19398 19808
rect 20622 19796 20628 19808
rect 20680 19836 20686 19848
rect 21269 19839 21327 19845
rect 21269 19836 21281 19839
rect 20680 19808 21281 19836
rect 20680 19796 20686 19808
rect 21269 19805 21281 19808
rect 21315 19805 21327 19839
rect 21269 19799 21327 19805
rect 28166 19796 28172 19848
rect 28224 19836 28230 19848
rect 28445 19839 28503 19845
rect 28445 19836 28457 19839
rect 28224 19808 28457 19836
rect 28224 19796 28230 19808
rect 28445 19805 28457 19808
rect 28491 19805 28503 19839
rect 28445 19799 28503 19805
rect 14369 19771 14427 19777
rect 14369 19737 14381 19771
rect 14415 19768 14427 19771
rect 16942 19768 16948 19780
rect 14415 19740 16948 19768
rect 14415 19737 14427 19740
rect 14369 19731 14427 19737
rect 16942 19728 16948 19740
rect 17000 19728 17006 19780
rect 17218 19728 17224 19780
rect 17276 19768 17282 19780
rect 17276 19740 17321 19768
rect 17276 19728 17282 19740
rect 17586 19728 17592 19780
rect 17644 19768 17650 19780
rect 17773 19771 17831 19777
rect 17773 19768 17785 19771
rect 17644 19740 17785 19768
rect 17644 19728 17650 19740
rect 17773 19737 17785 19740
rect 17819 19737 17831 19771
rect 17773 19731 17831 19737
rect 22557 19771 22615 19777
rect 22557 19737 22569 19771
rect 22603 19737 22615 19771
rect 22557 19731 22615 19737
rect 15654 19700 15660 19712
rect 14292 19672 15660 19700
rect 15654 19660 15660 19672
rect 15712 19660 15718 19712
rect 16301 19703 16359 19709
rect 16301 19669 16313 19703
rect 16347 19700 16359 19703
rect 19426 19700 19432 19712
rect 16347 19672 19432 19700
rect 16347 19669 16359 19672
rect 16301 19663 16359 19669
rect 19426 19660 19432 19672
rect 19484 19660 19490 19712
rect 22572 19700 22600 19731
rect 22646 19728 22652 19780
rect 22704 19768 22710 19780
rect 25682 19768 25688 19780
rect 22704 19740 22749 19768
rect 25643 19740 25688 19768
rect 22704 19728 22710 19740
rect 25682 19728 25688 19740
rect 25740 19728 25746 19780
rect 25777 19771 25835 19777
rect 25777 19737 25789 19771
rect 25823 19768 25835 19771
rect 25866 19768 25872 19780
rect 25823 19740 25872 19768
rect 25823 19737 25835 19740
rect 25777 19731 25835 19737
rect 25866 19728 25872 19740
rect 25924 19728 25930 19780
rect 26973 19771 27031 19777
rect 26973 19737 26985 19771
rect 27019 19768 27031 19771
rect 27154 19768 27160 19780
rect 27019 19740 27160 19768
rect 27019 19737 27031 19740
rect 26973 19731 27031 19737
rect 27154 19728 27160 19740
rect 27212 19728 27218 19780
rect 29564 19700 29592 19876
rect 30466 19864 30472 19876
rect 30524 19864 30530 19916
rect 34514 19904 34520 19916
rect 30668 19876 34520 19904
rect 29730 19796 29736 19848
rect 29788 19836 29794 19848
rect 30668 19845 30696 19876
rect 34514 19864 34520 19876
rect 34572 19864 34578 19916
rect 30193 19839 30251 19845
rect 30193 19836 30205 19839
rect 29788 19808 30205 19836
rect 29788 19796 29794 19808
rect 30193 19805 30205 19808
rect 30239 19805 30251 19839
rect 30193 19799 30251 19805
rect 30653 19839 30711 19845
rect 30653 19805 30665 19839
rect 30699 19805 30711 19839
rect 30653 19799 30711 19805
rect 31481 19839 31539 19845
rect 31481 19805 31493 19839
rect 31527 19805 31539 19839
rect 31481 19799 31539 19805
rect 31496 19768 31524 19799
rect 30024 19740 31524 19768
rect 30024 19709 30052 19740
rect 22572 19672 29592 19700
rect 30009 19703 30067 19709
rect 30009 19669 30021 19703
rect 30055 19669 30067 19703
rect 31294 19700 31300 19712
rect 31255 19672 31300 19700
rect 30009 19663 30067 19669
rect 31294 19660 31300 19672
rect 31352 19660 31358 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 4893 19499 4951 19505
rect 4893 19465 4905 19499
rect 4939 19496 4951 19499
rect 5074 19496 5080 19508
rect 4939 19468 5080 19496
rect 4939 19465 4951 19468
rect 4893 19459 4951 19465
rect 5074 19456 5080 19468
rect 5132 19456 5138 19508
rect 9766 19496 9772 19508
rect 9727 19468 9772 19496
rect 9766 19456 9772 19468
rect 9824 19456 9830 19508
rect 10965 19499 11023 19505
rect 10965 19465 10977 19499
rect 11011 19465 11023 19499
rect 10965 19459 11023 19465
rect 11793 19499 11851 19505
rect 11793 19465 11805 19499
rect 11839 19496 11851 19499
rect 12894 19496 12900 19508
rect 11839 19468 12900 19496
rect 11839 19465 11851 19468
rect 11793 19459 11851 19465
rect 6822 19428 6828 19440
rect 1596 19400 6828 19428
rect 1596 19369 1624 19400
rect 6822 19388 6828 19400
rect 6880 19388 6886 19440
rect 10980 19428 11008 19459
rect 12894 19456 12900 19468
rect 12952 19456 12958 19508
rect 17129 19499 17187 19505
rect 17129 19465 17141 19499
rect 17175 19496 17187 19499
rect 17218 19496 17224 19508
rect 17175 19468 17224 19496
rect 17175 19465 17187 19468
rect 17129 19459 17187 19465
rect 17218 19456 17224 19468
rect 17276 19456 17282 19508
rect 17586 19456 17592 19508
rect 17644 19496 17650 19508
rect 19245 19499 19303 19505
rect 17644 19468 18552 19496
rect 17644 19456 17650 19468
rect 10980 19400 12020 19428
rect 1581 19363 1639 19369
rect 1581 19329 1593 19363
rect 1627 19329 1639 19363
rect 1581 19323 1639 19329
rect 3418 19320 3424 19372
rect 3476 19360 3482 19372
rect 4249 19363 4307 19369
rect 4249 19360 4261 19363
rect 3476 19332 4261 19360
rect 3476 19320 3482 19332
rect 4249 19329 4261 19332
rect 4295 19329 4307 19363
rect 4249 19323 4307 19329
rect 5442 19320 5448 19372
rect 5500 19360 5506 19372
rect 5537 19363 5595 19369
rect 5537 19360 5549 19363
rect 5500 19332 5549 19360
rect 5500 19320 5506 19332
rect 5537 19329 5549 19332
rect 5583 19329 5595 19363
rect 5537 19323 5595 19329
rect 9677 19363 9735 19369
rect 9677 19329 9689 19363
rect 9723 19360 9735 19363
rect 9950 19360 9956 19372
rect 9723 19332 9956 19360
rect 9723 19329 9735 19332
rect 9677 19323 9735 19329
rect 9950 19320 9956 19332
rect 10008 19360 10014 19372
rect 10686 19360 10692 19372
rect 10008 19332 10692 19360
rect 10008 19320 10014 19332
rect 10686 19320 10692 19332
rect 10744 19320 10750 19372
rect 11149 19363 11207 19369
rect 11149 19329 11161 19363
rect 11195 19360 11207 19363
rect 11514 19360 11520 19372
rect 11195 19332 11520 19360
rect 11195 19329 11207 19332
rect 11149 19323 11207 19329
rect 11514 19320 11520 19332
rect 11572 19320 11578 19372
rect 11992 19369 12020 19400
rect 13630 19388 13636 19440
rect 13688 19428 13694 19440
rect 14185 19431 14243 19437
rect 14185 19428 14197 19431
rect 13688 19400 14197 19428
rect 13688 19388 13694 19400
rect 14185 19397 14197 19400
rect 14231 19397 14243 19431
rect 16482 19428 16488 19440
rect 14185 19391 14243 19397
rect 15212 19400 16488 19428
rect 15212 19372 15240 19400
rect 16482 19388 16488 19400
rect 16540 19388 16546 19440
rect 17954 19428 17960 19440
rect 17915 19400 17960 19428
rect 17954 19388 17960 19400
rect 18012 19388 18018 19440
rect 18524 19437 18552 19468
rect 19245 19465 19257 19499
rect 19291 19496 19303 19499
rect 20714 19496 20720 19508
rect 19291 19468 20720 19496
rect 19291 19465 19303 19468
rect 19245 19459 19303 19465
rect 20714 19456 20720 19468
rect 20772 19456 20778 19508
rect 20809 19499 20867 19505
rect 20809 19465 20821 19499
rect 20855 19496 20867 19499
rect 21174 19496 21180 19508
rect 20855 19468 21180 19496
rect 20855 19465 20867 19468
rect 20809 19459 20867 19465
rect 21174 19456 21180 19468
rect 21232 19456 21238 19508
rect 22097 19499 22155 19505
rect 22097 19465 22109 19499
rect 22143 19496 22155 19499
rect 22646 19496 22652 19508
rect 22143 19468 22652 19496
rect 22143 19465 22155 19468
rect 22097 19459 22155 19465
rect 22646 19456 22652 19468
rect 22704 19456 22710 19508
rect 27154 19496 27160 19508
rect 27115 19468 27160 19496
rect 27154 19456 27160 19468
rect 27212 19456 27218 19508
rect 18509 19431 18567 19437
rect 18509 19397 18521 19431
rect 18555 19397 18567 19431
rect 18509 19391 18567 19397
rect 25682 19388 25688 19440
rect 25740 19428 25746 19440
rect 32582 19428 32588 19440
rect 25740 19400 32588 19428
rect 25740 19388 25746 19400
rect 32582 19388 32588 19400
rect 32640 19388 32646 19440
rect 11977 19363 12035 19369
rect 11977 19329 11989 19363
rect 12023 19329 12035 19363
rect 15194 19360 15200 19372
rect 15155 19332 15200 19360
rect 11977 19323 12035 19329
rect 15194 19320 15200 19332
rect 15252 19320 15258 19372
rect 15841 19363 15899 19369
rect 15841 19329 15853 19363
rect 15887 19360 15899 19363
rect 17034 19360 17040 19372
rect 15887 19332 17040 19360
rect 15887 19329 15899 19332
rect 15841 19323 15899 19329
rect 17034 19320 17040 19332
rect 17092 19320 17098 19372
rect 17310 19360 17316 19372
rect 17271 19332 17316 19360
rect 17310 19320 17316 19332
rect 17368 19320 17374 19372
rect 19426 19360 19432 19372
rect 19387 19332 19432 19360
rect 19426 19320 19432 19332
rect 19484 19320 19490 19372
rect 20530 19320 20536 19372
rect 20588 19360 20594 19372
rect 22005 19363 22063 19369
rect 22005 19360 22017 19363
rect 20588 19332 22017 19360
rect 20588 19320 20594 19332
rect 22005 19329 22017 19332
rect 22051 19329 22063 19363
rect 22005 19323 22063 19329
rect 22094 19320 22100 19372
rect 22152 19360 22158 19372
rect 25130 19360 25136 19372
rect 22152 19332 25136 19360
rect 22152 19320 22158 19332
rect 25130 19320 25136 19332
rect 25188 19320 25194 19372
rect 27338 19360 27344 19372
rect 27299 19332 27344 19360
rect 27338 19320 27344 19332
rect 27396 19320 27402 19372
rect 30098 19320 30104 19372
rect 30156 19360 30162 19372
rect 30469 19363 30527 19369
rect 30469 19360 30481 19363
rect 30156 19332 30481 19360
rect 30156 19320 30162 19332
rect 30469 19329 30481 19332
rect 30515 19329 30527 19363
rect 30469 19323 30527 19329
rect 4433 19295 4491 19301
rect 4433 19261 4445 19295
rect 4479 19292 4491 19295
rect 14090 19292 14096 19304
rect 4479 19264 5396 19292
rect 14051 19264 14096 19292
rect 4479 19261 4491 19264
rect 4433 19255 4491 19261
rect 5368 19233 5396 19264
rect 14090 19252 14096 19264
rect 14148 19252 14154 19304
rect 15378 19292 15384 19304
rect 15339 19264 15384 19292
rect 15378 19252 15384 19264
rect 15436 19252 15442 19304
rect 17865 19295 17923 19301
rect 17865 19261 17877 19295
rect 17911 19292 17923 19295
rect 19242 19292 19248 19304
rect 17911 19264 19248 19292
rect 17911 19261 17923 19264
rect 17865 19255 17923 19261
rect 19242 19252 19248 19264
rect 19300 19252 19306 19304
rect 20162 19292 20168 19304
rect 20123 19264 20168 19292
rect 20162 19252 20168 19264
rect 20220 19252 20226 19304
rect 20346 19292 20352 19304
rect 20307 19264 20352 19292
rect 20346 19252 20352 19264
rect 20404 19252 20410 19304
rect 29822 19292 29828 19304
rect 29783 19264 29828 19292
rect 29822 19252 29828 19264
rect 29880 19252 29886 19304
rect 30009 19295 30067 19301
rect 30009 19261 30021 19295
rect 30055 19292 30067 19295
rect 31294 19292 31300 19304
rect 30055 19264 31300 19292
rect 30055 19261 30067 19264
rect 30009 19255 30067 19261
rect 31294 19252 31300 19264
rect 31352 19252 31358 19304
rect 5353 19227 5411 19233
rect 5353 19193 5365 19227
rect 5399 19193 5411 19227
rect 5353 19187 5411 19193
rect 14645 19227 14703 19233
rect 14645 19193 14657 19227
rect 14691 19224 14703 19227
rect 32674 19224 32680 19236
rect 14691 19196 32680 19224
rect 14691 19193 14703 19196
rect 14645 19187 14703 19193
rect 32674 19184 32680 19196
rect 32732 19184 32738 19236
rect 1762 19156 1768 19168
rect 1723 19128 1768 19156
rect 1762 19116 1768 19128
rect 1820 19116 1826 19168
rect 5810 19116 5816 19168
rect 5868 19156 5874 19168
rect 14182 19156 14188 19168
rect 5868 19128 14188 19156
rect 5868 19116 5874 19128
rect 14182 19116 14188 19128
rect 14240 19156 14246 19168
rect 14826 19156 14832 19168
rect 14240 19128 14832 19156
rect 14240 19116 14246 19128
rect 14826 19116 14832 19128
rect 14884 19116 14890 19168
rect 18782 19116 18788 19168
rect 18840 19156 18846 19168
rect 22094 19156 22100 19168
rect 18840 19128 22100 19156
rect 18840 19116 18846 19128
rect 22094 19116 22100 19128
rect 22152 19116 22158 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 4525 18955 4583 18961
rect 4525 18921 4537 18955
rect 4571 18952 4583 18955
rect 4614 18952 4620 18964
rect 4571 18924 4620 18952
rect 4571 18921 4583 18924
rect 4525 18915 4583 18921
rect 4614 18912 4620 18924
rect 4672 18912 4678 18964
rect 5169 18955 5227 18961
rect 5169 18921 5181 18955
rect 5215 18952 5227 18955
rect 14182 18952 14188 18964
rect 5215 18924 14188 18952
rect 5215 18921 5227 18924
rect 5169 18915 5227 18921
rect 14182 18912 14188 18924
rect 14240 18912 14246 18964
rect 14277 18955 14335 18961
rect 14277 18921 14289 18955
rect 14323 18952 14335 18955
rect 15102 18952 15108 18964
rect 14323 18924 15108 18952
rect 14323 18921 14335 18924
rect 14277 18915 14335 18921
rect 15102 18912 15108 18924
rect 15160 18912 15166 18964
rect 15838 18912 15844 18964
rect 15896 18952 15902 18964
rect 16117 18955 16175 18961
rect 16117 18952 16129 18955
rect 15896 18924 16129 18952
rect 15896 18912 15902 18924
rect 16117 18921 16129 18924
rect 16163 18921 16175 18955
rect 16117 18915 16175 18921
rect 16390 18912 16396 18964
rect 16448 18952 16454 18964
rect 20162 18952 20168 18964
rect 16448 18924 20168 18952
rect 16448 18912 16454 18924
rect 20162 18912 20168 18924
rect 20220 18912 20226 18964
rect 22370 18952 22376 18964
rect 22331 18924 22376 18952
rect 22370 18912 22376 18924
rect 22428 18912 22434 18964
rect 4982 18844 4988 18896
rect 5040 18884 5046 18896
rect 5040 18856 8708 18884
rect 5040 18844 5046 18856
rect 5626 18816 5632 18828
rect 4448 18788 5632 18816
rect 4448 18757 4476 18788
rect 5626 18776 5632 18788
rect 5684 18776 5690 18828
rect 5813 18819 5871 18825
rect 5813 18785 5825 18819
rect 5859 18816 5871 18819
rect 5902 18816 5908 18828
rect 5859 18788 5908 18816
rect 5859 18785 5871 18788
rect 5813 18779 5871 18785
rect 5902 18776 5908 18788
rect 5960 18776 5966 18828
rect 6086 18816 6092 18828
rect 6047 18788 6092 18816
rect 6086 18776 6092 18788
rect 6144 18776 6150 18828
rect 8680 18816 8708 18856
rect 9398 18844 9404 18896
rect 9456 18884 9462 18896
rect 23566 18884 23572 18896
rect 9456 18856 23572 18884
rect 9456 18844 9462 18856
rect 23566 18844 23572 18856
rect 23624 18844 23630 18896
rect 30558 18884 30564 18896
rect 24596 18856 30564 18884
rect 16850 18816 16856 18828
rect 8680 18788 16856 18816
rect 16850 18776 16856 18788
rect 16908 18776 16914 18828
rect 17034 18776 17040 18828
rect 17092 18816 17098 18828
rect 17221 18819 17279 18825
rect 17221 18816 17233 18819
rect 17092 18788 17233 18816
rect 17092 18776 17098 18788
rect 17221 18785 17233 18788
rect 17267 18785 17279 18819
rect 17221 18779 17279 18785
rect 18233 18819 18291 18825
rect 18233 18785 18245 18819
rect 18279 18816 18291 18819
rect 18506 18816 18512 18828
rect 18279 18788 18512 18816
rect 18279 18785 18291 18788
rect 18233 18779 18291 18785
rect 18506 18776 18512 18788
rect 18564 18776 18570 18828
rect 24596 18825 24624 18856
rect 30558 18844 30564 18856
rect 30616 18844 30622 18896
rect 24581 18819 24639 18825
rect 24581 18816 24593 18819
rect 22066 18788 24593 18816
rect 4433 18751 4491 18757
rect 4433 18717 4445 18751
rect 4479 18717 4491 18751
rect 5074 18748 5080 18760
rect 5035 18720 5080 18748
rect 4433 18711 4491 18717
rect 5074 18708 5080 18720
rect 5132 18708 5138 18760
rect 6914 18748 6920 18760
rect 6875 18720 6920 18748
rect 6914 18708 6920 18720
rect 6972 18708 6978 18760
rect 7098 18748 7104 18760
rect 7059 18720 7104 18748
rect 7098 18708 7104 18720
rect 7156 18708 7162 18760
rect 8018 18748 8024 18760
rect 7979 18720 8024 18748
rect 8018 18708 8024 18720
rect 8076 18708 8082 18760
rect 11057 18751 11115 18757
rect 11057 18717 11069 18751
rect 11103 18748 11115 18751
rect 11514 18748 11520 18760
rect 11103 18720 11520 18748
rect 11103 18717 11115 18720
rect 11057 18711 11115 18717
rect 11514 18708 11520 18720
rect 11572 18708 11578 18760
rect 14461 18751 14519 18757
rect 14461 18717 14473 18751
rect 14507 18748 14519 18751
rect 14642 18748 14648 18760
rect 14507 18720 14648 18748
rect 14507 18717 14519 18720
rect 14461 18711 14519 18717
rect 14642 18708 14648 18720
rect 14700 18708 14706 18760
rect 14826 18708 14832 18760
rect 14884 18748 14890 18760
rect 16025 18751 16083 18757
rect 16025 18748 16037 18751
rect 14884 18720 16037 18748
rect 14884 18708 14890 18720
rect 16025 18717 16037 18720
rect 16071 18717 16083 18751
rect 16025 18711 16083 18717
rect 20625 18751 20683 18757
rect 20625 18717 20637 18751
rect 20671 18748 20683 18751
rect 20806 18748 20812 18760
rect 20671 18720 20812 18748
rect 20671 18717 20683 18720
rect 20625 18711 20683 18717
rect 20806 18708 20812 18720
rect 20864 18708 20870 18760
rect 21542 18748 21548 18760
rect 21503 18720 21548 18748
rect 21542 18708 21548 18720
rect 21600 18708 21606 18760
rect 22066 18692 22094 18788
rect 24581 18785 24593 18788
rect 24627 18785 24639 18819
rect 24581 18779 24639 18785
rect 29822 18776 29828 18828
rect 29880 18816 29886 18828
rect 29917 18819 29975 18825
rect 29917 18816 29929 18819
rect 29880 18788 29929 18816
rect 29880 18776 29886 18788
rect 29917 18785 29929 18788
rect 29963 18785 29975 18819
rect 29917 18779 29975 18785
rect 22278 18748 22284 18760
rect 22239 18720 22284 18748
rect 22278 18708 22284 18720
rect 22336 18708 22342 18760
rect 24762 18748 24768 18760
rect 24723 18720 24768 18748
rect 24762 18708 24768 18720
rect 24820 18708 24826 18760
rect 28261 18751 28319 18757
rect 28261 18717 28273 18751
rect 28307 18748 28319 18751
rect 28442 18748 28448 18760
rect 28307 18720 28448 18748
rect 28307 18717 28319 18720
rect 28261 18711 28319 18717
rect 28442 18708 28448 18720
rect 28500 18708 28506 18760
rect 4798 18640 4804 18692
rect 4856 18680 4862 18692
rect 5905 18683 5963 18689
rect 5905 18680 5917 18683
rect 4856 18652 5917 18680
rect 4856 18640 4862 18652
rect 5905 18649 5917 18652
rect 5951 18649 5963 18683
rect 8113 18683 8171 18689
rect 8113 18680 8125 18683
rect 5905 18643 5963 18649
rect 6564 18652 8125 18680
rect 5166 18572 5172 18624
rect 5224 18612 5230 18624
rect 6564 18612 6592 18652
rect 8113 18649 8125 18652
rect 8159 18649 8171 18683
rect 11974 18680 11980 18692
rect 11936 18652 11980 18680
rect 8113 18643 8171 18649
rect 11974 18640 11980 18652
rect 12032 18640 12038 18692
rect 12069 18683 12127 18689
rect 12069 18649 12081 18683
rect 12115 18649 12127 18683
rect 12069 18643 12127 18649
rect 12621 18683 12679 18689
rect 12621 18649 12633 18683
rect 12667 18680 12679 18683
rect 12710 18680 12716 18692
rect 12667 18652 12716 18680
rect 12667 18649 12679 18652
rect 12621 18643 12679 18649
rect 7558 18612 7564 18624
rect 5224 18584 6592 18612
rect 7519 18584 7564 18612
rect 5224 18572 5230 18584
rect 7558 18572 7564 18584
rect 7616 18572 7622 18624
rect 9214 18612 9220 18624
rect 9175 18584 9220 18612
rect 9214 18572 9220 18584
rect 9272 18572 9278 18624
rect 11149 18615 11207 18621
rect 11149 18581 11161 18615
rect 11195 18612 11207 18615
rect 12084 18612 12112 18643
rect 12710 18640 12716 18652
rect 12768 18640 12774 18692
rect 14182 18640 14188 18692
rect 14240 18680 14246 18692
rect 16390 18680 16396 18692
rect 14240 18652 16396 18680
rect 14240 18640 14246 18652
rect 16390 18640 16396 18652
rect 16448 18640 16454 18692
rect 16942 18640 16948 18692
rect 17000 18680 17006 18692
rect 17313 18683 17371 18689
rect 17313 18680 17325 18683
rect 17000 18652 17325 18680
rect 17000 18640 17006 18652
rect 17313 18649 17325 18652
rect 17359 18649 17371 18683
rect 17313 18643 17371 18649
rect 19242 18640 19248 18692
rect 19300 18680 19306 18692
rect 22002 18680 22008 18692
rect 19300 18652 22008 18680
rect 19300 18640 19306 18652
rect 22002 18640 22008 18652
rect 22060 18652 22094 18692
rect 22060 18640 22066 18652
rect 11195 18584 12112 18612
rect 11195 18581 11207 18584
rect 11149 18575 11207 18581
rect 19426 18572 19432 18624
rect 19484 18612 19490 18624
rect 20717 18615 20775 18621
rect 20717 18612 20729 18615
rect 19484 18584 20729 18612
rect 19484 18572 19490 18584
rect 20717 18581 20729 18584
rect 20763 18581 20775 18615
rect 21358 18612 21364 18624
rect 21319 18584 21364 18612
rect 20717 18575 20775 18581
rect 21358 18572 21364 18584
rect 21416 18572 21422 18624
rect 24578 18572 24584 18624
rect 24636 18612 24642 18624
rect 25225 18615 25283 18621
rect 25225 18612 25237 18615
rect 24636 18584 25237 18612
rect 24636 18572 24642 18584
rect 25225 18581 25237 18584
rect 25271 18581 25283 18615
rect 28074 18612 28080 18624
rect 28035 18584 28080 18612
rect 25225 18575 25283 18581
rect 28074 18572 28080 18584
rect 28132 18572 28138 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 1581 18411 1639 18417
rect 1581 18377 1593 18411
rect 1627 18408 1639 18411
rect 3786 18408 3792 18420
rect 1627 18380 3792 18408
rect 1627 18377 1639 18380
rect 1581 18371 1639 18377
rect 3786 18368 3792 18380
rect 3844 18368 3850 18420
rect 5537 18411 5595 18417
rect 5537 18377 5549 18411
rect 5583 18408 5595 18411
rect 6914 18408 6920 18420
rect 5583 18380 6920 18408
rect 5583 18377 5595 18380
rect 5537 18371 5595 18377
rect 6914 18368 6920 18380
rect 6972 18368 6978 18420
rect 12158 18408 12164 18420
rect 12119 18380 12164 18408
rect 12158 18368 12164 18380
rect 12216 18368 12222 18420
rect 17221 18411 17279 18417
rect 12636 18380 16804 18408
rect 7374 18300 7380 18352
rect 7432 18340 7438 18352
rect 8481 18343 8539 18349
rect 8481 18340 8493 18343
rect 7432 18312 8493 18340
rect 7432 18300 7438 18312
rect 8481 18309 8493 18312
rect 8527 18309 8539 18343
rect 9398 18340 9404 18352
rect 9359 18312 9404 18340
rect 8481 18303 8539 18309
rect 9398 18300 9404 18312
rect 9456 18300 9462 18352
rect 10226 18300 10232 18352
rect 10284 18340 10290 18352
rect 12636 18340 12664 18380
rect 12802 18340 12808 18352
rect 10284 18312 12664 18340
rect 12763 18312 12808 18340
rect 10284 18300 10290 18312
rect 12802 18300 12808 18312
rect 12860 18300 12866 18352
rect 12894 18300 12900 18352
rect 12952 18340 12958 18352
rect 14182 18340 14188 18352
rect 12952 18312 12997 18340
rect 14143 18312 14188 18340
rect 12952 18300 12958 18312
rect 14182 18300 14188 18312
rect 14240 18300 14246 18352
rect 1762 18272 1768 18284
rect 1723 18244 1768 18272
rect 1762 18232 1768 18244
rect 1820 18232 1826 18284
rect 5350 18272 5356 18284
rect 5311 18244 5356 18272
rect 5350 18232 5356 18244
rect 5408 18232 5414 18284
rect 7282 18272 7288 18284
rect 7243 18244 7288 18272
rect 7282 18232 7288 18244
rect 7340 18232 7346 18284
rect 10042 18272 10048 18284
rect 10003 18244 10048 18272
rect 10042 18232 10048 18244
rect 10100 18232 10106 18284
rect 12066 18272 12072 18284
rect 12027 18244 12072 18272
rect 12066 18232 12072 18244
rect 12124 18232 12130 18284
rect 16776 18272 16804 18380
rect 17221 18377 17233 18411
rect 17267 18408 17279 18411
rect 17310 18408 17316 18420
rect 17267 18380 17316 18408
rect 17267 18377 17279 18380
rect 17221 18371 17279 18377
rect 17310 18368 17316 18380
rect 17368 18368 17374 18420
rect 20806 18408 20812 18420
rect 18432 18380 20812 18408
rect 16850 18300 16856 18352
rect 16908 18340 16914 18352
rect 17957 18343 18015 18349
rect 17957 18340 17969 18343
rect 16908 18312 17969 18340
rect 16908 18300 16914 18312
rect 17957 18309 17969 18312
rect 18003 18309 18015 18343
rect 17957 18303 18015 18309
rect 17402 18272 17408 18284
rect 16776 18244 17408 18272
rect 17402 18232 17408 18244
rect 17460 18232 17466 18284
rect 17865 18275 17923 18281
rect 17865 18241 17877 18275
rect 17911 18272 17923 18275
rect 18432 18272 18460 18380
rect 20806 18368 20812 18380
rect 20864 18368 20870 18420
rect 23937 18411 23995 18417
rect 23937 18377 23949 18411
rect 23983 18408 23995 18411
rect 24762 18408 24768 18420
rect 23983 18380 24768 18408
rect 23983 18377 23995 18380
rect 23937 18371 23995 18377
rect 24762 18368 24768 18380
rect 24820 18368 24826 18420
rect 28442 18408 28448 18420
rect 28403 18380 28448 18408
rect 28442 18368 28448 18380
rect 28500 18368 28506 18420
rect 18690 18340 18696 18352
rect 18651 18312 18696 18340
rect 18690 18300 18696 18312
rect 18748 18300 18754 18352
rect 21177 18343 21235 18349
rect 21177 18309 21189 18343
rect 21223 18340 21235 18343
rect 24578 18340 24584 18352
rect 21223 18312 24584 18340
rect 21223 18309 21235 18312
rect 21177 18303 21235 18309
rect 24578 18300 24584 18312
rect 24636 18300 24642 18352
rect 24673 18343 24731 18349
rect 24673 18309 24685 18343
rect 24719 18340 24731 18343
rect 25777 18343 25835 18349
rect 25777 18340 25789 18343
rect 24719 18312 25789 18340
rect 24719 18309 24731 18312
rect 24673 18303 24731 18309
rect 25777 18309 25789 18312
rect 25823 18309 25835 18343
rect 25777 18303 25835 18309
rect 17911 18244 18460 18272
rect 17911 18241 17923 18244
rect 17865 18235 17923 18241
rect 20162 18232 20168 18284
rect 20220 18272 20226 18284
rect 20533 18275 20591 18281
rect 20533 18272 20545 18275
rect 20220 18244 20545 18272
rect 20220 18232 20226 18244
rect 20533 18241 20545 18244
rect 20579 18241 20591 18275
rect 20533 18235 20591 18241
rect 20717 18275 20775 18281
rect 20717 18241 20729 18275
rect 20763 18272 20775 18275
rect 21358 18272 21364 18284
rect 20763 18244 21364 18272
rect 20763 18241 20775 18244
rect 20717 18235 20775 18241
rect 21358 18232 21364 18244
rect 21416 18232 21422 18284
rect 22002 18272 22008 18284
rect 21963 18244 22008 18272
rect 22002 18232 22008 18244
rect 22060 18232 22066 18284
rect 23845 18275 23903 18281
rect 23845 18241 23857 18275
rect 23891 18241 23903 18275
rect 25682 18272 25688 18284
rect 25643 18244 25688 18272
rect 23845 18235 23903 18241
rect 7558 18164 7564 18216
rect 7616 18204 7622 18216
rect 8389 18207 8447 18213
rect 8389 18204 8401 18207
rect 7616 18176 8401 18204
rect 7616 18164 7622 18176
rect 8389 18173 8401 18176
rect 8435 18204 8447 18207
rect 11054 18204 11060 18216
rect 8435 18176 11060 18204
rect 8435 18173 8447 18176
rect 8389 18167 8447 18173
rect 11054 18164 11060 18176
rect 11112 18164 11118 18216
rect 12802 18164 12808 18216
rect 12860 18204 12866 18216
rect 13081 18207 13139 18213
rect 13081 18204 13093 18207
rect 12860 18176 13093 18204
rect 12860 18164 12866 18176
rect 13081 18173 13093 18176
rect 13127 18173 13139 18207
rect 13081 18167 13139 18173
rect 14093 18207 14151 18213
rect 14093 18173 14105 18207
rect 14139 18173 14151 18207
rect 14093 18167 14151 18173
rect 6822 18096 6828 18148
rect 6880 18136 6886 18148
rect 7101 18139 7159 18145
rect 7101 18136 7113 18139
rect 6880 18108 7113 18136
rect 6880 18096 6886 18108
rect 7101 18105 7113 18108
rect 7147 18105 7159 18139
rect 7101 18099 7159 18105
rect 9861 18071 9919 18077
rect 9861 18037 9873 18071
rect 9907 18068 9919 18071
rect 11974 18068 11980 18080
rect 9907 18040 11980 18068
rect 9907 18037 9919 18040
rect 9861 18031 9919 18037
rect 11974 18028 11980 18040
rect 12032 18028 12038 18080
rect 14108 18068 14136 18167
rect 14366 18164 14372 18216
rect 14424 18204 14430 18216
rect 14737 18207 14795 18213
rect 14737 18204 14749 18207
rect 14424 18176 14749 18204
rect 14424 18164 14430 18176
rect 14737 18173 14749 18176
rect 14783 18204 14795 18207
rect 14826 18204 14832 18216
rect 14783 18176 14832 18204
rect 14783 18173 14795 18176
rect 14737 18167 14795 18173
rect 14826 18164 14832 18176
rect 14884 18164 14890 18216
rect 18598 18204 18604 18216
rect 18559 18176 18604 18204
rect 18598 18164 18604 18176
rect 18656 18164 18662 18216
rect 18877 18207 18935 18213
rect 18877 18173 18889 18207
rect 18923 18173 18935 18207
rect 22186 18204 22192 18216
rect 22147 18176 22192 18204
rect 18877 18167 18935 18173
rect 15838 18096 15844 18148
rect 15896 18136 15902 18148
rect 18892 18136 18920 18167
rect 22186 18164 22192 18176
rect 22244 18164 22250 18216
rect 23860 18204 23888 18235
rect 25682 18232 25688 18244
rect 25740 18232 25746 18284
rect 27341 18275 27399 18281
rect 27341 18241 27353 18275
rect 27387 18272 27399 18275
rect 27706 18272 27712 18284
rect 27387 18244 27712 18272
rect 27387 18241 27399 18244
rect 27341 18235 27399 18241
rect 27706 18232 27712 18244
rect 27764 18232 27770 18284
rect 28629 18275 28687 18281
rect 28629 18241 28641 18275
rect 28675 18241 28687 18275
rect 31202 18272 31208 18284
rect 31163 18244 31208 18272
rect 28629 18235 28687 18241
rect 24854 18204 24860 18216
rect 23860 18176 24860 18204
rect 24854 18164 24860 18176
rect 24912 18164 24918 18216
rect 25225 18207 25283 18213
rect 25225 18173 25237 18207
rect 25271 18204 25283 18207
rect 25958 18204 25964 18216
rect 25271 18176 25964 18204
rect 25271 18173 25283 18176
rect 25225 18167 25283 18173
rect 25958 18164 25964 18176
rect 26016 18164 26022 18216
rect 27522 18204 27528 18216
rect 27483 18176 27528 18204
rect 27522 18164 27528 18176
rect 27580 18164 27586 18216
rect 27614 18164 27620 18216
rect 27672 18204 27678 18216
rect 28644 18204 28672 18235
rect 31202 18232 31208 18244
rect 31260 18232 31266 18284
rect 29086 18204 29092 18216
rect 27672 18176 28672 18204
rect 29047 18176 29092 18204
rect 27672 18164 27678 18176
rect 29086 18164 29092 18176
rect 29144 18164 29150 18216
rect 24394 18136 24400 18148
rect 15896 18108 24400 18136
rect 15896 18096 15902 18108
rect 24394 18096 24400 18108
rect 24452 18096 24458 18148
rect 17126 18068 17132 18080
rect 14108 18040 17132 18068
rect 17126 18028 17132 18040
rect 17184 18068 17190 18080
rect 22373 18071 22431 18077
rect 22373 18068 22385 18071
rect 17184 18040 22385 18068
rect 17184 18028 17190 18040
rect 22373 18037 22385 18040
rect 22419 18037 22431 18071
rect 22373 18031 22431 18037
rect 27985 18071 28043 18077
rect 27985 18037 27997 18071
rect 28031 18068 28043 18071
rect 28258 18068 28264 18080
rect 28031 18040 28264 18068
rect 28031 18037 28043 18040
rect 27985 18031 28043 18037
rect 28258 18028 28264 18040
rect 28316 18028 28322 18080
rect 31018 18068 31024 18080
rect 30979 18040 31024 18068
rect 31018 18028 31024 18040
rect 31076 18028 31082 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 5442 17864 5448 17876
rect 5403 17836 5448 17864
rect 5442 17824 5448 17836
rect 5500 17824 5506 17876
rect 8389 17867 8447 17873
rect 8389 17833 8401 17867
rect 8435 17864 8447 17867
rect 10042 17864 10048 17876
rect 8435 17836 10048 17864
rect 8435 17833 8447 17836
rect 8389 17827 8447 17833
rect 10042 17824 10048 17836
rect 10100 17824 10106 17876
rect 11054 17864 11060 17876
rect 11015 17836 11060 17864
rect 11054 17824 11060 17836
rect 11112 17824 11118 17876
rect 13630 17864 13636 17876
rect 13591 17836 13636 17864
rect 13630 17824 13636 17836
rect 13688 17824 13694 17876
rect 14182 17824 14188 17876
rect 14240 17864 14246 17876
rect 14369 17867 14427 17873
rect 14369 17864 14381 17867
rect 14240 17836 14381 17864
rect 14240 17824 14246 17836
rect 14369 17833 14381 17836
rect 14415 17833 14427 17867
rect 14369 17827 14427 17833
rect 17037 17867 17095 17873
rect 17037 17833 17049 17867
rect 17083 17864 17095 17867
rect 17126 17864 17132 17876
rect 17083 17836 17132 17864
rect 17083 17833 17095 17836
rect 17037 17827 17095 17833
rect 17126 17824 17132 17836
rect 17184 17824 17190 17876
rect 21542 17824 21548 17876
rect 21600 17864 21606 17876
rect 21821 17867 21879 17873
rect 21821 17864 21833 17867
rect 21600 17836 21833 17864
rect 21600 17824 21606 17836
rect 21821 17833 21833 17836
rect 21867 17833 21879 17867
rect 21821 17827 21879 17833
rect 22186 17824 22192 17876
rect 22244 17864 22250 17876
rect 22557 17867 22615 17873
rect 22557 17864 22569 17867
rect 22244 17836 22569 17864
rect 22244 17824 22250 17836
rect 22557 17833 22569 17836
rect 22603 17833 22615 17867
rect 22557 17827 22615 17833
rect 26881 17867 26939 17873
rect 26881 17833 26893 17867
rect 26927 17864 26939 17867
rect 27522 17864 27528 17876
rect 26927 17836 27528 17864
rect 26927 17833 26939 17836
rect 26881 17827 26939 17833
rect 27522 17824 27528 17836
rect 27580 17824 27586 17876
rect 2133 17799 2191 17805
rect 2133 17765 2145 17799
rect 2179 17765 2191 17799
rect 2133 17759 2191 17765
rect 6917 17799 6975 17805
rect 6917 17765 6929 17799
rect 6963 17765 6975 17799
rect 6917 17759 6975 17765
rect 7653 17799 7711 17805
rect 7653 17765 7665 17799
rect 7699 17796 7711 17799
rect 8294 17796 8300 17808
rect 7699 17768 8300 17796
rect 7699 17765 7711 17768
rect 7653 17759 7711 17765
rect 2148 17728 2176 17759
rect 4157 17731 4215 17737
rect 4157 17728 4169 17731
rect 2148 17700 4169 17728
rect 4157 17697 4169 17700
rect 4203 17697 4215 17731
rect 6932 17728 6960 17759
rect 8294 17756 8300 17768
rect 8352 17756 8358 17808
rect 10410 17796 10416 17808
rect 8588 17768 10416 17796
rect 6932 17700 7880 17728
rect 4157 17691 4215 17697
rect 2314 17660 2320 17672
rect 2275 17632 2320 17660
rect 2314 17620 2320 17632
rect 2372 17620 2378 17672
rect 3237 17663 3295 17669
rect 3237 17629 3249 17663
rect 3283 17660 3295 17663
rect 3973 17663 4031 17669
rect 3973 17660 3985 17663
rect 3283 17632 3985 17660
rect 3283 17629 3295 17632
rect 3237 17623 3295 17629
rect 3973 17629 3985 17632
rect 4019 17629 4031 17663
rect 5626 17660 5632 17672
rect 5539 17632 5632 17660
rect 3973 17623 4031 17629
rect 5626 17620 5632 17632
rect 5684 17660 5690 17672
rect 5902 17660 5908 17672
rect 5684 17632 5908 17660
rect 5684 17620 5690 17632
rect 5902 17620 5908 17632
rect 5960 17620 5966 17672
rect 6270 17660 6276 17672
rect 6231 17632 6276 17660
rect 6270 17620 6276 17632
rect 6328 17620 6334 17672
rect 7101 17663 7159 17669
rect 7101 17629 7113 17663
rect 7147 17660 7159 17663
rect 7742 17660 7748 17672
rect 7147 17632 7748 17660
rect 7147 17629 7159 17632
rect 7101 17623 7159 17629
rect 7742 17620 7748 17632
rect 7800 17620 7806 17672
rect 7852 17669 7880 17700
rect 7837 17663 7895 17669
rect 7837 17629 7849 17663
rect 7883 17629 7895 17663
rect 7837 17623 7895 17629
rect 7926 17620 7932 17672
rect 7984 17660 7990 17672
rect 8588 17669 8616 17768
rect 10410 17756 10416 17768
rect 10468 17756 10474 17808
rect 10502 17756 10508 17808
rect 10560 17796 10566 17808
rect 24118 17796 24124 17808
rect 10560 17768 24124 17796
rect 10560 17756 10566 17768
rect 24118 17756 24124 17768
rect 24176 17756 24182 17808
rect 28258 17756 28264 17808
rect 28316 17796 28322 17808
rect 28353 17799 28411 17805
rect 28353 17796 28365 17799
rect 28316 17768 28365 17796
rect 28316 17756 28322 17768
rect 28353 17765 28365 17768
rect 28399 17765 28411 17799
rect 28353 17759 28411 17765
rect 9214 17728 9220 17740
rect 9175 17700 9220 17728
rect 9214 17688 9220 17700
rect 9272 17688 9278 17740
rect 10689 17731 10747 17737
rect 10689 17697 10701 17731
rect 10735 17728 10747 17731
rect 11054 17728 11060 17740
rect 10735 17700 11060 17728
rect 10735 17697 10747 17700
rect 10689 17691 10747 17697
rect 11054 17688 11060 17700
rect 11112 17728 11118 17740
rect 11330 17728 11336 17740
rect 11112 17700 11336 17728
rect 11112 17688 11118 17700
rect 11330 17688 11336 17700
rect 11388 17688 11394 17740
rect 11885 17731 11943 17737
rect 11885 17697 11897 17731
rect 11931 17728 11943 17731
rect 12618 17728 12624 17740
rect 11931 17700 12624 17728
rect 11931 17697 11943 17700
rect 11885 17691 11943 17697
rect 12618 17688 12624 17700
rect 12676 17688 12682 17740
rect 16390 17728 16396 17740
rect 16351 17700 16396 17728
rect 16390 17688 16396 17700
rect 16448 17688 16454 17740
rect 16574 17728 16580 17740
rect 16535 17700 16580 17728
rect 16574 17688 16580 17700
rect 16632 17688 16638 17740
rect 18598 17688 18604 17740
rect 18656 17728 18662 17740
rect 18693 17731 18751 17737
rect 18693 17728 18705 17731
rect 18656 17700 18705 17728
rect 18656 17688 18662 17700
rect 18693 17697 18705 17700
rect 18739 17697 18751 17731
rect 20073 17731 20131 17737
rect 20073 17728 20085 17731
rect 18693 17691 18751 17697
rect 18800 17700 20085 17728
rect 8573 17663 8631 17669
rect 8573 17660 8585 17663
rect 7984 17632 8585 17660
rect 7984 17620 7990 17632
rect 8573 17629 8585 17632
rect 8619 17629 8631 17663
rect 10870 17660 10876 17672
rect 10831 17632 10876 17660
rect 8573 17623 8631 17629
rect 10870 17620 10876 17632
rect 10928 17620 10934 17672
rect 13541 17663 13599 17669
rect 13541 17629 13553 17663
rect 13587 17629 13599 17663
rect 13541 17623 13599 17629
rect 8294 17552 8300 17604
rect 8352 17592 8358 17604
rect 9309 17595 9367 17601
rect 9309 17592 9321 17595
rect 8352 17564 9321 17592
rect 8352 17552 8358 17564
rect 9309 17561 9321 17564
rect 9355 17561 9367 17595
rect 9858 17592 9864 17604
rect 9819 17564 9864 17592
rect 9309 17555 9367 17561
rect 9858 17552 9864 17564
rect 9916 17552 9922 17604
rect 11974 17592 11980 17604
rect 11935 17564 11980 17592
rect 11974 17552 11980 17564
rect 12032 17552 12038 17604
rect 12526 17592 12532 17604
rect 12487 17564 12532 17592
rect 12526 17552 12532 17564
rect 12584 17552 12590 17604
rect 4614 17524 4620 17536
rect 4575 17496 4620 17524
rect 4614 17484 4620 17496
rect 4672 17484 4678 17536
rect 5442 17484 5448 17536
rect 5500 17524 5506 17536
rect 6089 17527 6147 17533
rect 6089 17524 6101 17527
rect 5500 17496 6101 17524
rect 5500 17484 5506 17496
rect 6089 17493 6101 17496
rect 6135 17493 6147 17527
rect 6089 17487 6147 17493
rect 11790 17484 11796 17536
rect 11848 17524 11854 17536
rect 13556 17524 13584 17623
rect 13814 17620 13820 17672
rect 13872 17660 13878 17672
rect 14277 17663 14335 17669
rect 14277 17660 14289 17663
rect 13872 17632 14289 17660
rect 13872 17620 13878 17632
rect 14277 17629 14289 17632
rect 14323 17660 14335 17663
rect 15010 17660 15016 17672
rect 14323 17632 15016 17660
rect 14323 17629 14335 17632
rect 14277 17623 14335 17629
rect 15010 17620 15016 17632
rect 15068 17620 15074 17672
rect 16666 17620 16672 17672
rect 16724 17660 16730 17672
rect 18800 17660 18828 17700
rect 20073 17697 20085 17700
rect 20119 17728 20131 17731
rect 24854 17728 24860 17740
rect 20119 17700 20484 17728
rect 20119 17697 20131 17700
rect 20073 17691 20131 17697
rect 16724 17632 18828 17660
rect 16724 17620 16730 17632
rect 19797 17595 19855 17601
rect 19797 17561 19809 17595
rect 19843 17561 19855 17595
rect 19797 17555 19855 17561
rect 19889 17595 19947 17601
rect 19889 17561 19901 17595
rect 19935 17592 19947 17595
rect 19978 17592 19984 17604
rect 19935 17564 19984 17592
rect 19935 17561 19947 17564
rect 19889 17555 19947 17561
rect 11848 17496 13584 17524
rect 11848 17484 11854 17496
rect 14642 17484 14648 17536
rect 14700 17524 14706 17536
rect 19242 17524 19248 17536
rect 14700 17496 19248 17524
rect 14700 17484 14706 17496
rect 19242 17484 19248 17496
rect 19300 17484 19306 17536
rect 19812 17524 19840 17555
rect 19978 17552 19984 17564
rect 20036 17552 20042 17604
rect 20456 17592 20484 17700
rect 22020 17700 24860 17728
rect 22020 17669 22048 17700
rect 24854 17688 24860 17700
rect 24912 17688 24918 17740
rect 28074 17688 28080 17740
rect 28132 17728 28138 17740
rect 28169 17731 28227 17737
rect 28169 17728 28181 17731
rect 28132 17700 28181 17728
rect 28132 17688 28138 17700
rect 28169 17697 28181 17700
rect 28215 17697 28227 17731
rect 28169 17691 28227 17697
rect 22005 17663 22063 17669
rect 22005 17629 22017 17663
rect 22051 17629 22063 17663
rect 22462 17660 22468 17672
rect 22375 17632 22468 17660
rect 22005 17623 22063 17629
rect 22462 17620 22468 17632
rect 22520 17660 22526 17672
rect 26789 17663 26847 17669
rect 22520 17632 26740 17660
rect 22520 17620 22526 17632
rect 24210 17592 24216 17604
rect 20456 17564 24216 17592
rect 24210 17552 24216 17564
rect 24268 17552 24274 17604
rect 26712 17592 26740 17632
rect 26789 17629 26801 17663
rect 26835 17660 26847 17663
rect 27614 17660 27620 17672
rect 26835 17632 27620 17660
rect 26835 17629 26847 17632
rect 26789 17623 26847 17629
rect 27614 17620 27620 17632
rect 27672 17620 27678 17672
rect 27985 17663 28043 17669
rect 27985 17629 27997 17663
rect 28031 17660 28043 17663
rect 29086 17660 29092 17672
rect 28031 17632 29092 17660
rect 28031 17629 28043 17632
rect 27985 17623 28043 17629
rect 29086 17620 29092 17632
rect 29144 17620 29150 17672
rect 31018 17660 31024 17672
rect 30979 17632 31024 17660
rect 31018 17620 31024 17632
rect 31076 17620 31082 17672
rect 31202 17592 31208 17604
rect 26712 17564 31208 17592
rect 31202 17552 31208 17564
rect 31260 17552 31266 17604
rect 23474 17524 23480 17536
rect 19812 17496 23480 17524
rect 23474 17484 23480 17496
rect 23532 17524 23538 17536
rect 25866 17524 25872 17536
rect 23532 17496 25872 17524
rect 23532 17484 23538 17496
rect 25866 17484 25872 17496
rect 25924 17484 25930 17536
rect 30374 17484 30380 17536
rect 30432 17524 30438 17536
rect 30837 17527 30895 17533
rect 30837 17524 30849 17527
rect 30432 17496 30849 17524
rect 30432 17484 30438 17496
rect 30837 17493 30849 17496
rect 30883 17493 30895 17527
rect 30837 17487 30895 17493
rect 31941 17527 31999 17533
rect 31941 17493 31953 17527
rect 31987 17524 31999 17527
rect 32398 17524 32404 17536
rect 31987 17496 32404 17524
rect 31987 17493 31999 17496
rect 31941 17487 31999 17493
rect 32398 17484 32404 17496
rect 32456 17484 32462 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 3234 17280 3240 17332
rect 3292 17320 3298 17332
rect 5905 17323 5963 17329
rect 3292 17292 5856 17320
rect 3292 17280 3298 17292
rect 3053 17255 3111 17261
rect 3053 17221 3065 17255
rect 3099 17252 3111 17255
rect 4614 17252 4620 17264
rect 3099 17224 4620 17252
rect 3099 17221 3111 17224
rect 3053 17215 3111 17221
rect 4614 17212 4620 17224
rect 4672 17212 4678 17264
rect 5828 17252 5856 17292
rect 5905 17289 5917 17323
rect 5951 17320 5963 17323
rect 7098 17320 7104 17332
rect 5951 17292 7104 17320
rect 5951 17289 5963 17292
rect 5905 17283 5963 17289
rect 7098 17280 7104 17292
rect 7156 17280 7162 17332
rect 7653 17323 7711 17329
rect 7653 17289 7665 17323
rect 7699 17320 7711 17323
rect 10870 17320 10876 17332
rect 7699 17292 10876 17320
rect 7699 17289 7711 17292
rect 7653 17283 7711 17289
rect 10870 17280 10876 17292
rect 10928 17280 10934 17332
rect 17034 17280 17040 17332
rect 17092 17320 17098 17332
rect 17497 17323 17555 17329
rect 17497 17320 17509 17323
rect 17092 17292 17509 17320
rect 17092 17280 17098 17292
rect 17497 17289 17509 17292
rect 17543 17289 17555 17323
rect 17497 17283 17555 17289
rect 18509 17323 18567 17329
rect 18509 17289 18521 17323
rect 18555 17320 18567 17323
rect 18690 17320 18696 17332
rect 18555 17292 18696 17320
rect 18555 17289 18567 17292
rect 18509 17283 18567 17289
rect 18690 17280 18696 17292
rect 18748 17280 18754 17332
rect 19242 17280 19248 17332
rect 19300 17320 19306 17332
rect 20346 17320 20352 17332
rect 19300 17292 20352 17320
rect 19300 17280 19306 17292
rect 20346 17280 20352 17292
rect 20404 17280 20410 17332
rect 21450 17320 21456 17332
rect 20548 17292 21456 17320
rect 8294 17252 8300 17264
rect 5828 17224 8300 17252
rect 8294 17212 8300 17224
rect 8352 17212 8358 17264
rect 8757 17255 8815 17261
rect 8757 17221 8769 17255
rect 8803 17252 8815 17255
rect 9030 17252 9036 17264
rect 8803 17224 9036 17252
rect 8803 17221 8815 17224
rect 8757 17215 8815 17221
rect 9030 17212 9036 17224
rect 9088 17212 9094 17264
rect 12618 17252 12624 17264
rect 12176 17224 12624 17252
rect 3878 17184 3884 17196
rect 3839 17156 3884 17184
rect 3878 17144 3884 17156
rect 3936 17144 3942 17196
rect 4706 17184 4712 17196
rect 4667 17156 4712 17184
rect 4706 17144 4712 17156
rect 4764 17144 4770 17196
rect 5350 17184 5356 17196
rect 5311 17156 5356 17184
rect 5350 17144 5356 17156
rect 5408 17144 5414 17196
rect 5813 17187 5871 17193
rect 5813 17153 5825 17187
rect 5859 17184 5871 17187
rect 5994 17184 6000 17196
rect 5859 17156 6000 17184
rect 5859 17153 5871 17156
rect 5813 17147 5871 17153
rect 5994 17144 6000 17156
rect 6052 17184 6058 17196
rect 7193 17187 7251 17193
rect 7193 17184 7205 17187
rect 6052 17156 7205 17184
rect 6052 17144 6058 17156
rect 7193 17153 7205 17156
rect 7239 17153 7251 17187
rect 7193 17147 7251 17153
rect 7837 17187 7895 17193
rect 7837 17153 7849 17187
rect 7883 17153 7895 17187
rect 7837 17147 7895 17153
rect 2038 17076 2044 17128
rect 2096 17116 2102 17128
rect 2409 17119 2467 17125
rect 2409 17116 2421 17119
rect 2096 17088 2421 17116
rect 2096 17076 2102 17088
rect 2409 17085 2421 17088
rect 2455 17085 2467 17119
rect 2409 17079 2467 17085
rect 2593 17119 2651 17125
rect 2593 17085 2605 17119
rect 2639 17116 2651 17119
rect 3326 17116 3332 17128
rect 2639 17088 3332 17116
rect 2639 17085 2651 17088
rect 2593 17079 2651 17085
rect 3326 17076 3332 17088
rect 3384 17076 3390 17128
rect 3973 17119 4031 17125
rect 3973 17085 3985 17119
rect 4019 17116 4031 17119
rect 7852 17116 7880 17147
rect 8386 17144 8392 17196
rect 8444 17184 8450 17196
rect 10321 17187 10379 17193
rect 10321 17184 10333 17187
rect 8444 17156 8524 17184
rect 8444 17144 8450 17156
rect 4019 17088 6960 17116
rect 4019 17085 4031 17088
rect 3973 17079 4031 17085
rect 4525 17051 4583 17057
rect 4525 17017 4537 17051
rect 4571 17048 4583 17051
rect 6546 17048 6552 17060
rect 4571 17020 6552 17048
rect 4571 17017 4583 17020
rect 4525 17011 4583 17017
rect 6546 17008 6552 17020
rect 6604 17008 6610 17060
rect 5169 16983 5227 16989
rect 5169 16949 5181 16983
rect 5215 16980 5227 16983
rect 6822 16980 6828 16992
rect 5215 16952 6828 16980
rect 5215 16949 5227 16952
rect 5169 16943 5227 16949
rect 6822 16940 6828 16952
rect 6880 16940 6886 16992
rect 6932 16980 6960 17088
rect 7024 17088 7880 17116
rect 8496 17116 8524 17156
rect 9324 17156 10333 17184
rect 8665 17119 8723 17125
rect 8665 17116 8677 17119
rect 8496 17088 8677 17116
rect 7024 17057 7052 17088
rect 8665 17085 8677 17088
rect 8711 17085 8723 17119
rect 9324 17116 9352 17156
rect 10321 17153 10333 17156
rect 10367 17184 10379 17187
rect 12176 17184 12204 17224
rect 12618 17212 12624 17224
rect 12676 17212 12682 17264
rect 14826 17212 14832 17264
rect 14884 17252 14890 17264
rect 17862 17252 17868 17264
rect 14884 17224 17868 17252
rect 14884 17212 14890 17224
rect 17862 17212 17868 17224
rect 17920 17212 17926 17264
rect 12342 17184 12348 17196
rect 10367 17156 12204 17184
rect 12303 17156 12348 17184
rect 10367 17153 10379 17156
rect 10321 17147 10379 17153
rect 12342 17144 12348 17156
rect 12400 17144 12406 17196
rect 12986 17184 12992 17196
rect 12947 17156 12992 17184
rect 12986 17144 12992 17156
rect 13044 17144 13050 17196
rect 14550 17144 14556 17196
rect 14608 17184 14614 17196
rect 16117 17187 16175 17193
rect 16117 17184 16129 17187
rect 14608 17156 16129 17184
rect 14608 17144 14614 17156
rect 16117 17153 16129 17156
rect 16163 17153 16175 17187
rect 16117 17147 16175 17153
rect 16209 17187 16267 17193
rect 16209 17153 16221 17187
rect 16255 17184 16267 17187
rect 17037 17187 17095 17193
rect 17037 17184 17049 17187
rect 16255 17156 17049 17184
rect 16255 17153 16267 17156
rect 16209 17147 16267 17153
rect 17037 17153 17049 17156
rect 17083 17153 17095 17187
rect 18690 17184 18696 17196
rect 18651 17156 18696 17184
rect 17037 17147 17095 17153
rect 18690 17144 18696 17156
rect 18748 17144 18754 17196
rect 8665 17079 8723 17085
rect 9140 17088 9352 17116
rect 7009 17051 7067 17057
rect 7009 17017 7021 17051
rect 7055 17017 7067 17051
rect 7009 17011 7067 17017
rect 8018 17008 8024 17060
rect 8076 17048 8082 17060
rect 9140 17048 9168 17088
rect 9858 17076 9864 17128
rect 9916 17116 9922 17128
rect 16853 17119 16911 17125
rect 9916 17088 16804 17116
rect 9916 17076 9922 17088
rect 8076 17020 9168 17048
rect 9217 17051 9275 17057
rect 8076 17008 8082 17020
rect 9217 17017 9229 17051
rect 9263 17048 9275 17051
rect 16666 17048 16672 17060
rect 9263 17020 16672 17048
rect 9263 17017 9275 17020
rect 9217 17011 9275 17017
rect 16666 17008 16672 17020
rect 16724 17008 16730 17060
rect 8294 16980 8300 16992
rect 6932 16952 8300 16980
rect 8294 16940 8300 16952
rect 8352 16940 8358 16992
rect 8386 16940 8392 16992
rect 8444 16980 8450 16992
rect 10226 16980 10232 16992
rect 8444 16952 10232 16980
rect 8444 16940 8450 16952
rect 10226 16940 10232 16952
rect 10284 16940 10290 16992
rect 10413 16983 10471 16989
rect 10413 16949 10425 16983
rect 10459 16980 10471 16983
rect 10870 16980 10876 16992
rect 10459 16952 10876 16980
rect 10459 16949 10471 16952
rect 10413 16943 10471 16949
rect 10870 16940 10876 16952
rect 10928 16940 10934 16992
rect 11882 16940 11888 16992
rect 11940 16980 11946 16992
rect 12161 16983 12219 16989
rect 12161 16980 12173 16983
rect 11940 16952 12173 16980
rect 11940 16940 11946 16952
rect 12161 16949 12173 16952
rect 12207 16949 12219 16983
rect 12161 16943 12219 16949
rect 12805 16983 12863 16989
rect 12805 16949 12817 16983
rect 12851 16980 12863 16983
rect 15102 16980 15108 16992
rect 12851 16952 15108 16980
rect 12851 16949 12863 16952
rect 12805 16943 12863 16949
rect 15102 16940 15108 16952
rect 15160 16940 15166 16992
rect 16776 16980 16804 17088
rect 16853 17085 16865 17119
rect 16899 17116 16911 17119
rect 20548 17116 20576 17292
rect 21450 17280 21456 17292
rect 21508 17280 21514 17332
rect 23566 17280 23572 17332
rect 23624 17320 23630 17332
rect 25130 17320 25136 17332
rect 23624 17292 25136 17320
rect 23624 17280 23630 17292
rect 25130 17280 25136 17292
rect 25188 17280 25194 17332
rect 25685 17323 25743 17329
rect 25685 17289 25697 17323
rect 25731 17320 25743 17323
rect 25731 17292 27384 17320
rect 25731 17289 25743 17292
rect 25685 17283 25743 17289
rect 20714 17212 20720 17264
rect 20772 17252 20778 17264
rect 20809 17255 20867 17261
rect 20809 17252 20821 17255
rect 20772 17224 20821 17252
rect 20772 17212 20778 17224
rect 20809 17221 20821 17224
rect 20855 17221 20867 17255
rect 20809 17215 20867 17221
rect 21358 17212 21364 17264
rect 21416 17252 21422 17264
rect 23293 17255 23351 17261
rect 23293 17252 23305 17255
rect 21416 17224 23305 17252
rect 21416 17212 21422 17224
rect 23293 17221 23305 17224
rect 23339 17221 23351 17255
rect 23293 17215 23351 17221
rect 23385 17255 23443 17261
rect 23385 17221 23397 17255
rect 23431 17252 23443 17255
rect 23658 17252 23664 17264
rect 23431 17224 23664 17252
rect 23431 17221 23443 17224
rect 23385 17215 23443 17221
rect 23658 17212 23664 17224
rect 23716 17212 23722 17264
rect 27246 17252 27252 17264
rect 27207 17224 27252 17252
rect 27246 17212 27252 17224
rect 27304 17212 27310 17264
rect 27356 17261 27384 17292
rect 27341 17255 27399 17261
rect 27341 17221 27353 17255
rect 27387 17221 27399 17255
rect 32398 17252 32404 17264
rect 32359 17224 32404 17252
rect 27341 17215 27399 17221
rect 32398 17212 32404 17224
rect 32456 17212 32462 17264
rect 32490 17212 32496 17264
rect 32548 17252 32554 17264
rect 32548 17224 32593 17252
rect 32548 17212 32554 17224
rect 25593 17187 25651 17193
rect 25593 17153 25605 17187
rect 25639 17153 25651 17187
rect 38286 17184 38292 17196
rect 38247 17156 38292 17184
rect 25593 17147 25651 17153
rect 16899 17088 20576 17116
rect 20717 17119 20775 17125
rect 16899 17085 16911 17088
rect 16853 17079 16911 17085
rect 20717 17085 20729 17119
rect 20763 17116 20775 17119
rect 25608 17116 25636 17147
rect 38286 17144 38292 17156
rect 38344 17144 38350 17196
rect 27890 17116 27896 17128
rect 20763 17088 22048 17116
rect 25608 17088 27896 17116
rect 20763 17085 20775 17088
rect 20717 17079 20775 17085
rect 17862 17008 17868 17060
rect 17920 17048 17926 17060
rect 21269 17051 21327 17057
rect 21269 17048 21281 17051
rect 17920 17020 21281 17048
rect 17920 17008 17926 17020
rect 21269 17017 21281 17020
rect 21315 17017 21327 17051
rect 22020 17048 22048 17088
rect 27890 17076 27896 17088
rect 27948 17076 27954 17128
rect 30190 17116 30196 17128
rect 30151 17088 30196 17116
rect 30190 17076 30196 17088
rect 30248 17076 30254 17128
rect 32214 17076 32220 17128
rect 32272 17116 32278 17128
rect 32582 17116 32588 17128
rect 32272 17088 32588 17116
rect 32272 17076 32278 17088
rect 32582 17076 32588 17088
rect 32640 17116 32646 17128
rect 32677 17119 32735 17125
rect 32677 17116 32689 17119
rect 32640 17088 32689 17116
rect 32640 17076 32646 17088
rect 32677 17085 32689 17088
rect 32723 17085 32735 17119
rect 32677 17079 32735 17085
rect 23842 17048 23848 17060
rect 22020 17020 23704 17048
rect 23803 17020 23848 17048
rect 21269 17011 21327 17017
rect 21358 16980 21364 16992
rect 16776 16952 21364 16980
rect 21358 16940 21364 16952
rect 21416 16940 21422 16992
rect 21450 16940 21456 16992
rect 21508 16980 21514 16992
rect 22830 16980 22836 16992
rect 21508 16952 22836 16980
rect 21508 16940 21514 16952
rect 22830 16940 22836 16952
rect 22888 16940 22894 16992
rect 23676 16980 23704 17020
rect 23842 17008 23848 17020
rect 23900 17008 23906 17060
rect 27801 17051 27859 17057
rect 27801 17017 27813 17051
rect 27847 17048 27859 17051
rect 31110 17048 31116 17060
rect 27847 17020 31116 17048
rect 27847 17017 27859 17020
rect 27801 17011 27859 17017
rect 31110 17008 31116 17020
rect 31168 17008 31174 17060
rect 30558 16980 30564 16992
rect 23676 16952 30564 16980
rect 30558 16940 30564 16952
rect 30616 16940 30622 16992
rect 35894 16940 35900 16992
rect 35952 16980 35958 16992
rect 38105 16983 38163 16989
rect 38105 16980 38117 16983
rect 35952 16952 38117 16980
rect 35952 16940 35958 16952
rect 38105 16949 38117 16952
rect 38151 16949 38163 16983
rect 38105 16943 38163 16949
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 2314 16776 2320 16788
rect 2275 16748 2320 16776
rect 2314 16736 2320 16748
rect 2372 16736 2378 16788
rect 4706 16776 4712 16788
rect 4667 16748 4712 16776
rect 4706 16736 4712 16748
rect 4764 16736 4770 16788
rect 5350 16776 5356 16788
rect 5311 16748 5356 16776
rect 5350 16736 5356 16748
rect 5408 16736 5414 16788
rect 5626 16736 5632 16788
rect 5684 16776 5690 16788
rect 5684 16748 8616 16776
rect 5684 16736 5690 16748
rect 7926 16708 7932 16720
rect 3804 16680 7932 16708
rect 2501 16575 2559 16581
rect 2501 16541 2513 16575
rect 2547 16572 2559 16575
rect 3234 16572 3240 16584
rect 2547 16544 3240 16572
rect 2547 16541 2559 16544
rect 2501 16535 2559 16541
rect 3234 16532 3240 16544
rect 3292 16532 3298 16584
rect 3326 16532 3332 16584
rect 3384 16572 3390 16584
rect 3804 16572 3832 16680
rect 7926 16668 7932 16680
rect 7984 16668 7990 16720
rect 3878 16600 3884 16652
rect 3936 16640 3942 16652
rect 8018 16640 8024 16652
rect 3936 16612 8024 16640
rect 3936 16600 3942 16612
rect 4065 16575 4123 16581
rect 4065 16572 4077 16575
rect 3384 16544 3429 16572
rect 3804 16544 4077 16572
rect 3384 16532 3390 16544
rect 4065 16541 4077 16544
rect 4111 16541 4123 16575
rect 4890 16572 4896 16584
rect 4851 16544 4896 16572
rect 4065 16535 4123 16541
rect 4890 16532 4896 16544
rect 4948 16532 4954 16584
rect 5537 16575 5595 16581
rect 5537 16541 5549 16575
rect 5583 16572 5595 16575
rect 6362 16572 6368 16584
rect 5583 16544 6368 16572
rect 5583 16541 5595 16544
rect 5537 16535 5595 16541
rect 6362 16532 6368 16544
rect 6420 16532 6426 16584
rect 6564 16581 6592 16612
rect 8018 16600 8024 16612
rect 8076 16600 8082 16652
rect 8588 16640 8616 16748
rect 9030 16736 9036 16788
rect 9088 16776 9094 16788
rect 9217 16779 9275 16785
rect 9217 16776 9229 16779
rect 9088 16748 9229 16776
rect 9088 16736 9094 16748
rect 9217 16745 9229 16748
rect 9263 16745 9275 16779
rect 9217 16739 9275 16745
rect 12069 16779 12127 16785
rect 12069 16745 12081 16779
rect 12115 16776 12127 16779
rect 12342 16776 12348 16788
rect 12115 16748 12348 16776
rect 12115 16745 12127 16748
rect 12069 16739 12127 16745
rect 12342 16736 12348 16748
rect 12400 16736 12406 16788
rect 12618 16736 12624 16788
rect 12676 16776 12682 16788
rect 18509 16779 18567 16785
rect 12676 16748 14780 16776
rect 12676 16736 12682 16748
rect 12986 16708 12992 16720
rect 9140 16680 12992 16708
rect 9140 16640 9168 16680
rect 12986 16668 12992 16680
rect 13044 16668 13050 16720
rect 14366 16668 14372 16720
rect 14424 16708 14430 16720
rect 14642 16708 14648 16720
rect 14424 16680 14648 16708
rect 14424 16668 14430 16680
rect 14642 16668 14648 16680
rect 14700 16668 14706 16720
rect 14752 16708 14780 16748
rect 18509 16745 18521 16779
rect 18555 16776 18567 16779
rect 18690 16776 18696 16788
rect 18555 16748 18696 16776
rect 18555 16745 18567 16748
rect 18509 16739 18567 16745
rect 18690 16736 18696 16748
rect 18748 16736 18754 16788
rect 20346 16736 20352 16788
rect 20404 16776 20410 16788
rect 22462 16776 22468 16788
rect 20404 16748 22468 16776
rect 20404 16736 20410 16748
rect 22462 16736 22468 16748
rect 22520 16736 22526 16788
rect 23658 16776 23664 16788
rect 23619 16748 23664 16776
rect 23658 16736 23664 16748
rect 23716 16736 23722 16788
rect 30558 16776 30564 16788
rect 30519 16748 30564 16776
rect 30558 16736 30564 16748
rect 30616 16736 30622 16788
rect 32401 16779 32459 16785
rect 32401 16745 32413 16779
rect 32447 16776 32459 16779
rect 32490 16776 32496 16788
rect 32447 16748 32496 16776
rect 32447 16745 32459 16748
rect 32401 16739 32459 16745
rect 32490 16736 32496 16748
rect 32548 16736 32554 16788
rect 20714 16708 20720 16720
rect 14752 16680 20720 16708
rect 20714 16668 20720 16680
rect 20772 16668 20778 16720
rect 8588 16612 9168 16640
rect 6549 16575 6607 16581
rect 6549 16541 6561 16575
rect 6595 16541 6607 16575
rect 7190 16572 7196 16584
rect 7151 16544 7196 16572
rect 6549 16535 6607 16541
rect 7190 16532 7196 16544
rect 7248 16532 7254 16584
rect 7285 16575 7343 16581
rect 7285 16541 7297 16575
rect 7331 16572 7343 16575
rect 7374 16572 7380 16584
rect 7331 16544 7380 16572
rect 7331 16541 7343 16544
rect 7285 16535 7343 16541
rect 7374 16532 7380 16544
rect 7432 16532 7438 16584
rect 9140 16581 9168 16612
rect 16022 16600 16028 16652
rect 16080 16640 16086 16652
rect 30190 16640 30196 16652
rect 16080 16612 19334 16640
rect 30151 16612 30196 16640
rect 16080 16600 16086 16612
rect 9125 16575 9183 16581
rect 9125 16541 9137 16575
rect 9171 16541 9183 16575
rect 12250 16572 12256 16584
rect 12211 16544 12256 16572
rect 9125 16535 9183 16541
rect 12250 16532 12256 16544
rect 12308 16532 12314 16584
rect 17865 16575 17923 16581
rect 17865 16541 17877 16575
rect 17911 16541 17923 16575
rect 17865 16535 17923 16541
rect 8110 16464 8116 16516
rect 8168 16504 8174 16516
rect 14550 16504 14556 16516
rect 8168 16476 14556 16504
rect 8168 16464 8174 16476
rect 14550 16464 14556 16476
rect 14608 16464 14614 16516
rect 4157 16439 4215 16445
rect 4157 16405 4169 16439
rect 4203 16436 4215 16439
rect 4706 16436 4712 16448
rect 4203 16408 4712 16436
rect 4203 16405 4215 16408
rect 4157 16399 4215 16405
rect 4706 16396 4712 16408
rect 4764 16396 4770 16448
rect 6641 16439 6699 16445
rect 6641 16405 6653 16439
rect 6687 16436 6699 16439
rect 9398 16436 9404 16448
rect 6687 16408 9404 16436
rect 6687 16405 6699 16408
rect 6641 16399 6699 16405
rect 9398 16396 9404 16408
rect 9456 16396 9462 16448
rect 9490 16396 9496 16448
rect 9548 16436 9554 16448
rect 15654 16436 15660 16448
rect 9548 16408 15660 16436
rect 9548 16396 9554 16408
rect 15654 16396 15660 16408
rect 15712 16396 15718 16448
rect 17402 16396 17408 16448
rect 17460 16436 17466 16448
rect 17880 16436 17908 16535
rect 17954 16532 17960 16584
rect 18012 16572 18018 16584
rect 18690 16572 18696 16584
rect 18012 16544 18057 16572
rect 18651 16544 18696 16572
rect 18012 16532 18018 16544
rect 18690 16532 18696 16544
rect 18748 16532 18754 16584
rect 19306 16572 19334 16612
rect 30190 16600 30196 16612
rect 30248 16600 30254 16652
rect 30374 16640 30380 16652
rect 30335 16612 30380 16640
rect 30374 16600 30380 16612
rect 30432 16600 30438 16652
rect 20622 16572 20628 16584
rect 19306 16544 20628 16572
rect 20622 16532 20628 16544
rect 20680 16532 20686 16584
rect 23290 16532 23296 16584
rect 23348 16572 23354 16584
rect 23845 16575 23903 16581
rect 23845 16572 23857 16575
rect 23348 16544 23857 16572
rect 23348 16532 23354 16544
rect 23845 16541 23857 16544
rect 23891 16541 23903 16575
rect 23845 16535 23903 16541
rect 25961 16575 26019 16581
rect 25961 16541 25973 16575
rect 26007 16541 26019 16575
rect 25961 16535 26019 16541
rect 32585 16575 32643 16581
rect 32585 16541 32597 16575
rect 32631 16572 32643 16575
rect 33226 16572 33232 16584
rect 32631 16544 33088 16572
rect 33187 16544 33232 16572
rect 32631 16541 32643 16544
rect 32585 16535 32643 16541
rect 18046 16464 18052 16516
rect 18104 16504 18110 16516
rect 21358 16504 21364 16516
rect 18104 16476 21364 16504
rect 18104 16464 18110 16476
rect 21358 16464 21364 16476
rect 21416 16464 21422 16516
rect 25682 16504 25688 16516
rect 22066 16476 25688 16504
rect 17460 16408 17908 16436
rect 17460 16396 17466 16408
rect 17954 16396 17960 16448
rect 18012 16436 18018 16448
rect 18414 16436 18420 16448
rect 18012 16408 18420 16436
rect 18012 16396 18018 16408
rect 18414 16396 18420 16408
rect 18472 16396 18478 16448
rect 20898 16396 20904 16448
rect 20956 16436 20962 16448
rect 22066 16436 22094 16476
rect 25682 16464 25688 16476
rect 25740 16504 25746 16516
rect 25976 16504 26004 16535
rect 25740 16476 26004 16504
rect 25740 16464 25746 16476
rect 20956 16408 22094 16436
rect 25777 16439 25835 16445
rect 20956 16396 20962 16408
rect 25777 16405 25789 16439
rect 25823 16436 25835 16439
rect 27338 16436 27344 16448
rect 25823 16408 27344 16436
rect 25823 16405 25835 16408
rect 25777 16399 25835 16405
rect 27338 16396 27344 16408
rect 27396 16396 27402 16448
rect 33060 16445 33088 16544
rect 33226 16532 33232 16544
rect 33284 16532 33290 16584
rect 33045 16439 33103 16445
rect 33045 16405 33057 16439
rect 33091 16405 33103 16439
rect 33045 16399 33103 16405
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 4798 16232 4804 16244
rect 4759 16204 4804 16232
rect 4798 16192 4804 16204
rect 4856 16192 4862 16244
rect 5537 16235 5595 16241
rect 5537 16201 5549 16235
rect 5583 16232 5595 16235
rect 6270 16232 6276 16244
rect 5583 16204 6276 16232
rect 5583 16201 5595 16204
rect 5537 16195 5595 16201
rect 6270 16192 6276 16204
rect 6328 16192 6334 16244
rect 8570 16192 8576 16244
rect 8628 16232 8634 16244
rect 8628 16204 11284 16232
rect 8628 16192 8634 16204
rect 8662 16164 8668 16176
rect 2792 16136 8668 16164
rect 1578 16096 1584 16108
rect 1539 16068 1584 16096
rect 1578 16056 1584 16068
rect 1636 16056 1642 16108
rect 2792 16105 2820 16136
rect 8662 16124 8668 16136
rect 8720 16124 8726 16176
rect 10502 16164 10508 16176
rect 10463 16136 10508 16164
rect 10502 16124 10508 16136
rect 10560 16124 10566 16176
rect 10597 16167 10655 16173
rect 10597 16133 10609 16167
rect 10643 16164 10655 16167
rect 11146 16164 11152 16176
rect 10643 16136 11152 16164
rect 10643 16133 10655 16136
rect 10597 16127 10655 16133
rect 11146 16124 11152 16136
rect 11204 16124 11210 16176
rect 2777 16099 2835 16105
rect 2777 16065 2789 16099
rect 2823 16065 2835 16099
rect 2777 16059 2835 16065
rect 4709 16099 4767 16105
rect 4709 16065 4721 16099
rect 4755 16096 4767 16099
rect 5718 16096 5724 16108
rect 4755 16068 5724 16096
rect 4755 16065 4767 16068
rect 4709 16059 4767 16065
rect 5718 16056 5724 16068
rect 5776 16056 5782 16108
rect 6362 16056 6368 16108
rect 6420 16096 6426 16108
rect 10318 16096 10324 16108
rect 6420 16068 10324 16096
rect 6420 16056 6426 16068
rect 10318 16056 10324 16068
rect 10376 16056 10382 16108
rect 11256 16096 11284 16204
rect 11330 16192 11336 16244
rect 11388 16232 11394 16244
rect 11388 16204 20116 16232
rect 11388 16192 11394 16204
rect 12618 16124 12624 16176
rect 12676 16164 12682 16176
rect 18690 16164 18696 16176
rect 12676 16136 18696 16164
rect 12676 16124 12682 16136
rect 18690 16124 18696 16136
rect 18748 16124 18754 16176
rect 17954 16096 17960 16108
rect 11256 16068 17960 16096
rect 17954 16056 17960 16068
rect 18012 16056 18018 16108
rect 19794 16056 19800 16108
rect 19852 16056 19858 16108
rect 20088 16096 20116 16204
rect 20162 16192 20168 16244
rect 20220 16232 20226 16244
rect 23290 16232 23296 16244
rect 20220 16204 20265 16232
rect 23251 16204 23296 16232
rect 20220 16192 20226 16204
rect 23290 16192 23296 16204
rect 23348 16192 23354 16244
rect 27157 16235 27215 16241
rect 27157 16232 27169 16235
rect 25608 16204 27169 16232
rect 22278 16124 22284 16176
rect 22336 16164 22342 16176
rect 25608 16173 25636 16204
rect 27157 16201 27169 16204
rect 27203 16201 27215 16235
rect 27157 16195 27215 16201
rect 30558 16192 30564 16244
rect 30616 16232 30622 16244
rect 30837 16235 30895 16241
rect 30837 16232 30849 16235
rect 30616 16204 30849 16232
rect 30616 16192 30622 16204
rect 30837 16201 30849 16204
rect 30883 16201 30895 16235
rect 30837 16195 30895 16201
rect 25593 16167 25651 16173
rect 22336 16136 24164 16164
rect 22336 16124 22342 16136
rect 20438 16096 20444 16108
rect 20088 16068 20444 16096
rect 20438 16056 20444 16068
rect 20496 16056 20502 16108
rect 20714 16056 20720 16108
rect 20772 16096 20778 16108
rect 20901 16099 20959 16105
rect 20901 16096 20913 16099
rect 20772 16068 20913 16096
rect 20772 16056 20778 16068
rect 20901 16065 20913 16068
rect 20947 16096 20959 16099
rect 21174 16096 21180 16108
rect 20947 16068 21180 16096
rect 20947 16065 20959 16068
rect 20901 16059 20959 16065
rect 21174 16056 21180 16068
rect 21232 16056 21238 16108
rect 22465 16099 22523 16105
rect 22465 16065 22477 16099
rect 22511 16065 22523 16099
rect 22465 16059 22523 16065
rect 23477 16099 23535 16105
rect 23477 16065 23489 16099
rect 23523 16096 23535 16099
rect 23566 16096 23572 16108
rect 23523 16068 23572 16096
rect 23523 16065 23535 16068
rect 23477 16059 23535 16065
rect 7374 15988 7380 16040
rect 7432 16028 7438 16040
rect 10781 16031 10839 16037
rect 10781 16028 10793 16031
rect 7432 16000 10793 16028
rect 7432 15988 7438 16000
rect 10781 15997 10793 16000
rect 10827 15997 10839 16031
rect 10781 15991 10839 15997
rect 10962 15988 10968 16040
rect 11020 16028 11026 16040
rect 17586 16028 17592 16040
rect 11020 16000 17592 16028
rect 11020 15988 11026 16000
rect 17586 15988 17592 16000
rect 17644 15988 17650 16040
rect 17862 15988 17868 16040
rect 17920 16028 17926 16040
rect 18417 16031 18475 16037
rect 18417 16028 18429 16031
rect 17920 16000 18429 16028
rect 17920 15988 17926 16000
rect 18417 15997 18429 16000
rect 18463 15997 18475 16031
rect 18690 16028 18696 16040
rect 18417 15991 18475 15997
rect 18524 16000 18696 16028
rect 6270 15920 6276 15972
rect 6328 15960 6334 15972
rect 9490 15960 9496 15972
rect 6328 15932 9496 15960
rect 6328 15920 6334 15932
rect 9490 15920 9496 15932
rect 9548 15920 9554 15972
rect 12434 15960 12440 15972
rect 9600 15932 12440 15960
rect 1762 15892 1768 15904
rect 1723 15864 1768 15892
rect 1762 15852 1768 15864
rect 1820 15852 1826 15904
rect 2866 15892 2872 15904
rect 2827 15864 2872 15892
rect 2866 15852 2872 15864
rect 2924 15852 2930 15904
rect 6730 15852 6736 15904
rect 6788 15892 6794 15904
rect 9600 15892 9628 15932
rect 12434 15920 12440 15932
rect 12492 15920 12498 15972
rect 17954 15920 17960 15972
rect 18012 15960 18018 15972
rect 18524 15960 18552 16000
rect 18690 15988 18696 16000
rect 18748 15988 18754 16040
rect 18782 15988 18788 16040
rect 18840 16028 18846 16040
rect 22480 16028 22508 16059
rect 23566 16056 23572 16068
rect 23624 16056 23630 16108
rect 24136 16105 24164 16136
rect 25593 16133 25605 16167
rect 25639 16133 25651 16167
rect 28534 16164 28540 16176
rect 28495 16136 28540 16164
rect 25593 16127 25651 16133
rect 28534 16124 28540 16136
rect 28592 16124 28598 16176
rect 24121 16099 24179 16105
rect 24121 16065 24133 16099
rect 24167 16065 24179 16099
rect 27338 16096 27344 16108
rect 27299 16068 27344 16096
rect 24121 16059 24179 16065
rect 27338 16056 27344 16068
rect 27396 16056 27402 16108
rect 29733 16099 29791 16105
rect 29733 16096 29745 16099
rect 29380 16068 29745 16096
rect 23934 16028 23940 16040
rect 18840 16000 19748 16028
rect 22480 16000 23940 16028
rect 18840 15988 18846 16000
rect 18012 15932 18552 15960
rect 19720 15960 19748 16000
rect 23934 15988 23940 16000
rect 23992 15988 23998 16040
rect 25498 16028 25504 16040
rect 25459 16000 25504 16028
rect 25498 15988 25504 16000
rect 25556 15988 25562 16040
rect 25958 16028 25964 16040
rect 25919 16000 25964 16028
rect 25958 15988 25964 16000
rect 26016 15988 26022 16040
rect 28445 16031 28503 16037
rect 28445 15997 28457 16031
rect 28491 16028 28503 16031
rect 28626 16028 28632 16040
rect 28491 16000 28632 16028
rect 28491 15997 28503 16000
rect 28445 15991 28503 15997
rect 28626 15988 28632 16000
rect 28684 15988 28690 16040
rect 29089 16031 29147 16037
rect 29089 15997 29101 16031
rect 29135 16028 29147 16031
rect 29270 16028 29276 16040
rect 29135 16000 29276 16028
rect 29135 15997 29147 16000
rect 29089 15991 29147 15997
rect 29270 15988 29276 16000
rect 29328 15988 29334 16040
rect 25774 15960 25780 15972
rect 19720 15932 25780 15960
rect 18012 15920 18018 15932
rect 25774 15920 25780 15932
rect 25832 15920 25838 15972
rect 6788 15864 9628 15892
rect 6788 15852 6794 15864
rect 10502 15852 10508 15904
rect 10560 15892 10566 15904
rect 19242 15892 19248 15904
rect 10560 15864 19248 15892
rect 10560 15852 10566 15864
rect 19242 15852 19248 15864
rect 19300 15852 19306 15904
rect 20622 15852 20628 15904
rect 20680 15892 20686 15904
rect 20993 15895 21051 15901
rect 20993 15892 21005 15895
rect 20680 15864 21005 15892
rect 20680 15852 20686 15864
rect 20993 15861 21005 15864
rect 21039 15861 21051 15895
rect 22554 15892 22560 15904
rect 22515 15864 22560 15892
rect 20993 15855 21051 15861
rect 22554 15852 22560 15864
rect 22612 15852 22618 15904
rect 23937 15895 23995 15901
rect 23937 15861 23949 15895
rect 23983 15892 23995 15895
rect 29380 15892 29408 16068
rect 29733 16065 29745 16068
rect 29779 16065 29791 16099
rect 31478 16096 31484 16108
rect 31439 16068 31484 16096
rect 29733 16059 29791 16065
rect 31478 16056 31484 16068
rect 31536 16056 31542 16108
rect 38013 16099 38071 16105
rect 38013 16096 38025 16099
rect 35866 16068 38025 16096
rect 30193 16031 30251 16037
rect 30193 15997 30205 16031
rect 30239 15997 30251 16031
rect 30374 16028 30380 16040
rect 30335 16000 30380 16028
rect 30193 15991 30251 15997
rect 30208 15960 30236 15991
rect 30374 15988 30380 16000
rect 30432 15988 30438 16040
rect 31297 15963 31355 15969
rect 30208 15932 30972 15960
rect 23983 15864 29408 15892
rect 29549 15895 29607 15901
rect 23983 15861 23995 15864
rect 23937 15855 23995 15861
rect 29549 15861 29561 15895
rect 29595 15892 29607 15895
rect 30006 15892 30012 15904
rect 29595 15864 30012 15892
rect 29595 15861 29607 15864
rect 29549 15855 29607 15861
rect 30006 15852 30012 15864
rect 30064 15852 30070 15904
rect 30944 15892 30972 15932
rect 31297 15929 31309 15963
rect 31343 15960 31355 15963
rect 35866 15960 35894 16068
rect 38013 16065 38025 16068
rect 38059 16065 38071 16099
rect 38013 16059 38071 16065
rect 31343 15932 35894 15960
rect 31343 15929 31355 15932
rect 31297 15923 31355 15929
rect 33502 15892 33508 15904
rect 30944 15864 33508 15892
rect 33502 15852 33508 15864
rect 33560 15852 33566 15904
rect 38194 15892 38200 15904
rect 38155 15864 38200 15892
rect 38194 15852 38200 15864
rect 38252 15852 38258 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 8481 15691 8539 15697
rect 8481 15657 8493 15691
rect 8527 15688 8539 15691
rect 8570 15688 8576 15700
rect 8527 15660 8576 15688
rect 8527 15657 8539 15660
rect 8481 15651 8539 15657
rect 8570 15648 8576 15660
rect 8628 15648 8634 15700
rect 8662 15648 8668 15700
rect 8720 15688 8726 15700
rect 11330 15688 11336 15700
rect 8720 15660 11336 15688
rect 8720 15648 8726 15660
rect 11330 15648 11336 15660
rect 11388 15648 11394 15700
rect 18509 15691 18567 15697
rect 12728 15660 18460 15688
rect 6270 15620 6276 15632
rect 6231 15592 6276 15620
rect 6270 15580 6276 15592
rect 6328 15580 6334 15632
rect 10778 15580 10784 15632
rect 10836 15620 10842 15632
rect 10873 15623 10931 15629
rect 10873 15620 10885 15623
rect 10836 15592 10885 15620
rect 10836 15580 10842 15592
rect 10873 15589 10885 15592
rect 10919 15589 10931 15623
rect 10873 15583 10931 15589
rect 4525 15555 4583 15561
rect 4525 15521 4537 15555
rect 4571 15552 4583 15555
rect 6722 15555 6780 15561
rect 6722 15552 6734 15555
rect 4571 15524 6734 15552
rect 4571 15521 4583 15524
rect 4525 15515 4583 15521
rect 6722 15521 6734 15524
rect 6768 15552 6780 15555
rect 8754 15552 8760 15564
rect 6768 15524 8760 15552
rect 6768 15521 6780 15524
rect 6722 15515 6780 15521
rect 8754 15512 8760 15524
rect 8812 15552 8818 15564
rect 9125 15555 9183 15561
rect 9125 15552 9137 15555
rect 8812 15524 9137 15552
rect 8812 15512 8818 15524
rect 9125 15521 9137 15524
rect 9171 15552 9183 15555
rect 11333 15555 11391 15561
rect 11333 15552 11345 15555
rect 9171 15524 11345 15552
rect 9171 15521 9183 15524
rect 9125 15515 9183 15521
rect 11333 15521 11345 15524
rect 11379 15552 11391 15555
rect 12158 15552 12164 15564
rect 11379 15524 12164 15552
rect 11379 15521 11391 15524
rect 11333 15515 11391 15521
rect 12158 15512 12164 15524
rect 12216 15512 12222 15564
rect 8110 15444 8116 15496
rect 8168 15444 8174 15496
rect 10502 15444 10508 15496
rect 10560 15444 10566 15496
rect 12728 15470 12756 15660
rect 18432 15620 18460 15660
rect 18509 15657 18521 15691
rect 18555 15688 18567 15691
rect 19978 15688 19984 15700
rect 18555 15660 19984 15688
rect 18555 15657 18567 15660
rect 18509 15651 18567 15657
rect 19978 15648 19984 15660
rect 20036 15648 20042 15700
rect 20438 15648 20444 15700
rect 20496 15688 20502 15700
rect 22649 15691 22707 15697
rect 22649 15688 22661 15691
rect 20496 15660 22661 15688
rect 20496 15648 20502 15660
rect 22649 15657 22661 15660
rect 22695 15657 22707 15691
rect 22649 15651 22707 15657
rect 22738 15648 22744 15700
rect 22796 15688 22802 15700
rect 22796 15660 28948 15688
rect 22796 15648 22802 15660
rect 20806 15620 20812 15632
rect 18432 15592 20812 15620
rect 20806 15580 20812 15592
rect 20864 15580 20870 15632
rect 23658 15580 23664 15632
rect 23716 15620 23722 15632
rect 25501 15623 25559 15629
rect 25501 15620 25513 15623
rect 23716 15592 25513 15620
rect 23716 15580 23722 15592
rect 25501 15589 25513 15592
rect 25547 15589 25559 15623
rect 25501 15583 25559 15589
rect 28813 15623 28871 15629
rect 28813 15589 28825 15623
rect 28859 15589 28871 15623
rect 28920 15620 28948 15660
rect 30374 15648 30380 15700
rect 30432 15688 30438 15700
rect 31481 15691 31539 15697
rect 31481 15688 31493 15691
rect 30432 15660 31493 15688
rect 30432 15648 30438 15660
rect 31481 15657 31493 15660
rect 31527 15657 31539 15691
rect 33502 15688 33508 15700
rect 33463 15660 33508 15688
rect 31481 15651 31539 15657
rect 33502 15648 33508 15660
rect 33560 15648 33566 15700
rect 30469 15623 30527 15629
rect 30469 15620 30481 15623
rect 28920 15592 30481 15620
rect 28813 15583 28871 15589
rect 30469 15589 30481 15592
rect 30515 15589 30527 15623
rect 30469 15583 30527 15589
rect 13357 15555 13415 15561
rect 13357 15521 13369 15555
rect 13403 15552 13415 15555
rect 14458 15552 14464 15564
rect 13403 15524 14464 15552
rect 13403 15521 13415 15524
rect 13357 15515 13415 15521
rect 14458 15512 14464 15524
rect 14516 15512 14522 15564
rect 15289 15555 15347 15561
rect 15289 15521 15301 15555
rect 15335 15552 15347 15555
rect 17862 15552 17868 15564
rect 15335 15524 17868 15552
rect 15335 15521 15347 15524
rect 15289 15515 15347 15521
rect 17862 15512 17868 15524
rect 17920 15512 17926 15564
rect 21269 15555 21327 15561
rect 21269 15552 21281 15555
rect 18616 15524 21281 15552
rect 18616 15484 18644 15524
rect 21269 15521 21281 15524
rect 21315 15521 21327 15555
rect 23842 15552 23848 15564
rect 23803 15524 23848 15552
rect 21269 15515 21327 15521
rect 23842 15512 23848 15524
rect 23900 15512 23906 15564
rect 16698 15456 18644 15484
rect 18690 15444 18696 15496
rect 18748 15484 18754 15496
rect 20349 15487 20407 15493
rect 18748 15456 18793 15484
rect 18748 15444 18754 15456
rect 20349 15453 20361 15487
rect 20395 15484 20407 15487
rect 20714 15484 20720 15496
rect 20395 15456 20720 15484
rect 20395 15453 20407 15456
rect 20349 15447 20407 15453
rect 20714 15444 20720 15456
rect 20772 15444 20778 15496
rect 21177 15487 21235 15493
rect 21177 15453 21189 15487
rect 21223 15484 21235 15487
rect 21821 15487 21879 15493
rect 21821 15484 21833 15487
rect 21223 15456 21833 15484
rect 21223 15453 21235 15456
rect 21177 15447 21235 15453
rect 21821 15453 21833 15456
rect 21867 15484 21879 15487
rect 22462 15484 22468 15496
rect 21867 15456 22468 15484
rect 21867 15453 21879 15456
rect 21821 15447 21879 15453
rect 22462 15444 22468 15456
rect 22520 15484 22526 15496
rect 22557 15487 22615 15493
rect 22557 15484 22569 15487
rect 22520 15456 22569 15484
rect 22520 15444 22526 15456
rect 22557 15453 22569 15456
rect 22603 15453 22615 15487
rect 25038 15484 25044 15496
rect 24999 15456 25044 15484
rect 22557 15447 22615 15453
rect 25038 15444 25044 15456
rect 25096 15444 25102 15496
rect 25685 15487 25743 15493
rect 25685 15453 25697 15487
rect 25731 15453 25743 15487
rect 27522 15484 27528 15496
rect 27483 15456 27528 15484
rect 25685 15447 25743 15453
rect 4801 15419 4859 15425
rect 4801 15385 4813 15419
rect 4847 15385 4859 15419
rect 6026 15388 6684 15416
rect 4801 15379 4859 15385
rect 4816 15348 4844 15379
rect 5534 15348 5540 15360
rect 4816 15320 5540 15348
rect 5534 15308 5540 15320
rect 5592 15348 5598 15360
rect 6454 15348 6460 15360
rect 5592 15320 6460 15348
rect 5592 15308 5598 15320
rect 6454 15308 6460 15320
rect 6512 15308 6518 15360
rect 6656 15348 6684 15388
rect 6730 15376 6736 15428
rect 6788 15416 6794 15428
rect 7009 15419 7067 15425
rect 7009 15416 7021 15419
rect 6788 15388 7021 15416
rect 6788 15376 6794 15388
rect 7009 15385 7021 15388
rect 7055 15385 7067 15419
rect 7009 15379 7067 15385
rect 9401 15419 9459 15425
rect 9401 15385 9413 15419
rect 9447 15385 9459 15419
rect 9401 15379 9459 15385
rect 8662 15348 8668 15360
rect 6656 15320 8668 15348
rect 8662 15308 8668 15320
rect 8720 15308 8726 15360
rect 9416 15348 9444 15379
rect 11514 15376 11520 15428
rect 11572 15416 11578 15428
rect 11609 15419 11667 15425
rect 11609 15416 11621 15419
rect 11572 15388 11621 15416
rect 11572 15376 11578 15388
rect 11609 15385 11621 15388
rect 11655 15385 11667 15419
rect 11609 15379 11667 15385
rect 15565 15419 15623 15425
rect 15565 15385 15577 15419
rect 15611 15416 15623 15419
rect 15654 15416 15660 15428
rect 15611 15388 15660 15416
rect 15611 15385 15623 15388
rect 15565 15379 15623 15385
rect 15654 15376 15660 15388
rect 15712 15376 15718 15428
rect 17126 15376 17132 15428
rect 17184 15416 17190 15428
rect 17313 15419 17371 15425
rect 17313 15416 17325 15419
rect 17184 15388 17325 15416
rect 17184 15376 17190 15388
rect 17313 15385 17325 15388
rect 17359 15416 17371 15419
rect 19334 15416 19340 15428
rect 17359 15388 19340 15416
rect 17359 15385 17371 15388
rect 17313 15379 17371 15385
rect 19334 15376 19340 15388
rect 19392 15376 19398 15428
rect 20732 15416 20760 15444
rect 22002 15416 22008 15428
rect 20732 15388 22008 15416
rect 22002 15376 22008 15388
rect 22060 15376 22066 15428
rect 23385 15419 23443 15425
rect 23385 15385 23397 15419
rect 23431 15385 23443 15419
rect 23385 15379 23443 15385
rect 15010 15348 15016 15360
rect 9416 15320 15016 15348
rect 15010 15308 15016 15320
rect 15068 15308 15074 15360
rect 15102 15308 15108 15360
rect 15160 15348 15166 15360
rect 18690 15348 18696 15360
rect 15160 15320 18696 15348
rect 15160 15308 15166 15320
rect 18690 15308 18696 15320
rect 18748 15308 18754 15360
rect 20438 15348 20444 15360
rect 20399 15320 20444 15348
rect 20438 15308 20444 15320
rect 20496 15308 20502 15360
rect 21910 15348 21916 15360
rect 21871 15320 21916 15348
rect 21910 15308 21916 15320
rect 21968 15308 21974 15360
rect 23400 15348 23428 15379
rect 23474 15376 23480 15428
rect 23532 15416 23538 15428
rect 25700 15416 25728 15447
rect 27522 15444 27528 15456
rect 27580 15444 27586 15496
rect 28353 15487 28411 15493
rect 28353 15453 28365 15487
rect 28399 15484 28411 15487
rect 28828 15484 28856 15583
rect 29917 15555 29975 15561
rect 29917 15521 29929 15555
rect 29963 15552 29975 15555
rect 31018 15552 31024 15564
rect 29963 15524 31024 15552
rect 29963 15521 29975 15524
rect 29917 15515 29975 15521
rect 31018 15512 31024 15524
rect 31076 15512 31082 15564
rect 35894 15552 35900 15564
rect 32784 15524 35900 15552
rect 28399 15456 28856 15484
rect 28997 15487 29055 15493
rect 28399 15453 28411 15456
rect 28353 15447 28411 15453
rect 28997 15453 29009 15487
rect 29043 15453 29055 15487
rect 28997 15447 29055 15453
rect 23532 15388 23577 15416
rect 24872 15388 25728 15416
rect 23532 15376 23538 15388
rect 23750 15348 23756 15360
rect 23400 15320 23756 15348
rect 23750 15308 23756 15320
rect 23808 15308 23814 15360
rect 24872 15357 24900 15388
rect 25774 15376 25780 15428
rect 25832 15416 25838 15428
rect 26510 15416 26516 15428
rect 25832 15388 26516 15416
rect 25832 15376 25838 15388
rect 26510 15376 26516 15388
rect 26568 15416 26574 15428
rect 29012 15416 29040 15447
rect 31202 15444 31208 15496
rect 31260 15484 31266 15496
rect 32784 15493 32812 15524
rect 35894 15512 35900 15524
rect 35952 15512 35958 15564
rect 31389 15487 31447 15493
rect 31389 15484 31401 15487
rect 31260 15456 31401 15484
rect 31260 15444 31266 15456
rect 31389 15453 31401 15456
rect 31435 15453 31447 15487
rect 31389 15447 31447 15453
rect 32769 15487 32827 15493
rect 32769 15453 32781 15487
rect 32815 15453 32827 15487
rect 32769 15447 32827 15453
rect 33413 15487 33471 15493
rect 33413 15453 33425 15487
rect 33459 15484 33471 15487
rect 34606 15484 34612 15496
rect 33459 15456 34612 15484
rect 33459 15453 33471 15456
rect 33413 15447 33471 15453
rect 34606 15444 34612 15456
rect 34664 15444 34670 15496
rect 26568 15388 29040 15416
rect 26568 15376 26574 15388
rect 30006 15376 30012 15428
rect 30064 15416 30070 15428
rect 30064 15388 30109 15416
rect 30064 15376 30070 15388
rect 24857 15351 24915 15357
rect 24857 15317 24869 15351
rect 24903 15317 24915 15351
rect 27338 15348 27344 15360
rect 27299 15320 27344 15348
rect 24857 15311 24915 15317
rect 27338 15308 27344 15320
rect 27396 15308 27402 15360
rect 27430 15308 27436 15360
rect 27488 15348 27494 15360
rect 28169 15351 28227 15357
rect 28169 15348 28181 15351
rect 27488 15320 28181 15348
rect 27488 15308 27494 15320
rect 28169 15317 28181 15320
rect 28215 15317 28227 15351
rect 32858 15348 32864 15360
rect 32819 15320 32864 15348
rect 28169 15311 28227 15317
rect 32858 15308 32864 15320
rect 32916 15308 32922 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 13354 15144 13360 15156
rect 3896 15116 13360 15144
rect 3896 15085 3924 15116
rect 13354 15104 13360 15116
rect 13412 15104 13418 15156
rect 13909 15147 13967 15153
rect 13909 15113 13921 15147
rect 13955 15144 13967 15147
rect 15562 15144 15568 15156
rect 13955 15116 15568 15144
rect 13955 15113 13967 15116
rect 13909 15107 13967 15113
rect 15562 15104 15568 15116
rect 15620 15144 15626 15156
rect 16482 15144 16488 15156
rect 15620 15116 16488 15144
rect 15620 15104 15626 15116
rect 16482 15104 16488 15116
rect 16540 15104 16546 15156
rect 18690 15104 18696 15156
rect 18748 15144 18754 15156
rect 20622 15144 20628 15156
rect 18748 15116 20628 15144
rect 18748 15104 18754 15116
rect 20622 15104 20628 15116
rect 20680 15104 20686 15156
rect 20714 15104 20720 15156
rect 20772 15144 20778 15156
rect 23017 15147 23075 15153
rect 23017 15144 23029 15147
rect 20772 15116 23029 15144
rect 20772 15104 20778 15116
rect 23017 15113 23029 15116
rect 23063 15113 23075 15147
rect 23017 15107 23075 15113
rect 23474 15104 23480 15156
rect 23532 15144 23538 15156
rect 23661 15147 23719 15153
rect 23661 15144 23673 15147
rect 23532 15116 23673 15144
rect 23532 15104 23538 15116
rect 23661 15113 23673 15116
rect 23707 15113 23719 15147
rect 23661 15107 23719 15113
rect 26053 15147 26111 15153
rect 26053 15113 26065 15147
rect 26099 15113 26111 15147
rect 29273 15147 29331 15153
rect 29273 15144 29285 15147
rect 26053 15107 26111 15113
rect 28276 15116 29285 15144
rect 3881 15079 3939 15085
rect 3881 15045 3893 15079
rect 3927 15045 3939 15079
rect 3881 15039 3939 15045
rect 8570 15036 8576 15088
rect 8628 15076 8634 15088
rect 9033 15079 9091 15085
rect 9033 15076 9045 15079
rect 8628 15048 9045 15076
rect 8628 15036 8634 15048
rect 9033 15045 9045 15048
rect 9079 15045 9091 15079
rect 10962 15076 10968 15088
rect 10258 15048 10968 15076
rect 9033 15039 9091 15045
rect 10962 15036 10968 15048
rect 11020 15036 11026 15088
rect 17586 15076 17592 15088
rect 15962 15048 17592 15076
rect 17586 15036 17592 15048
rect 17644 15036 17650 15088
rect 20438 15076 20444 15088
rect 19642 15048 20444 15076
rect 20438 15036 20444 15048
rect 20496 15036 20502 15088
rect 26068 15076 26096 15107
rect 26068 15048 27384 15076
rect 1762 15008 1768 15020
rect 1723 14980 1768 15008
rect 1762 14968 1768 14980
rect 1820 14968 1826 15020
rect 4982 14968 4988 15020
rect 5040 14968 5046 15020
rect 8754 15008 8760 15020
rect 8715 14980 8760 15008
rect 8754 14968 8760 14980
rect 8812 14968 8818 15020
rect 12158 15008 12164 15020
rect 12119 14980 12164 15008
rect 12158 14968 12164 14980
rect 12216 14968 12222 15020
rect 14458 15008 14464 15020
rect 3510 14900 3516 14952
rect 3568 14940 3574 14952
rect 3605 14943 3663 14949
rect 3605 14940 3617 14943
rect 3568 14912 3617 14940
rect 3568 14900 3574 14912
rect 3605 14909 3617 14912
rect 3651 14909 3663 14943
rect 5350 14940 5356 14952
rect 5311 14912 5356 14940
rect 3605 14903 3663 14909
rect 5350 14900 5356 14912
rect 5408 14900 5414 14952
rect 12434 14940 12440 14952
rect 12395 14912 12440 14940
rect 12434 14900 12440 14912
rect 12492 14900 12498 14952
rect 13556 14872 13584 14994
rect 14419 14980 14464 15008
rect 14458 14968 14464 14980
rect 14516 14968 14522 15020
rect 17862 14968 17868 15020
rect 17920 15008 17926 15020
rect 18141 15011 18199 15017
rect 18141 15008 18153 15011
rect 17920 14980 18153 15008
rect 17920 14968 17926 14980
rect 18141 14977 18153 14980
rect 18187 14977 18199 15011
rect 18141 14971 18199 14977
rect 21818 14968 21824 15020
rect 21876 15008 21882 15020
rect 22281 15011 22339 15017
rect 22281 15008 22293 15011
rect 21876 14980 22293 15008
rect 21876 14968 21882 14980
rect 22281 14977 22293 14980
rect 22327 14977 22339 15011
rect 22281 14971 22339 14977
rect 22462 14968 22468 15020
rect 22520 15008 22526 15020
rect 22925 15011 22983 15017
rect 22925 15008 22937 15011
rect 22520 14980 22937 15008
rect 22520 14968 22526 14980
rect 22925 14977 22937 14980
rect 22971 14977 22983 15011
rect 22925 14971 22983 14977
rect 23474 14968 23480 15020
rect 23532 15008 23538 15020
rect 23569 15011 23627 15017
rect 23569 15008 23581 15011
rect 23532 14980 23581 15008
rect 23532 14968 23538 14980
rect 23569 14977 23581 14980
rect 23615 14977 23627 15011
rect 23569 14971 23627 14977
rect 24854 14968 24860 15020
rect 24912 15008 24918 15020
rect 27356 15017 27384 15048
rect 27982 15036 27988 15088
rect 28040 15076 28046 15088
rect 28276 15085 28304 15116
rect 29273 15113 29285 15116
rect 29319 15113 29331 15147
rect 29273 15107 29331 15113
rect 28169 15079 28227 15085
rect 28169 15076 28181 15079
rect 28040 15048 28181 15076
rect 28040 15036 28046 15048
rect 28169 15045 28181 15048
rect 28215 15045 28227 15079
rect 28169 15039 28227 15045
rect 28261 15079 28319 15085
rect 28261 15045 28273 15079
rect 28307 15045 28319 15079
rect 28261 15039 28319 15045
rect 26237 15011 26295 15017
rect 26237 15008 26249 15011
rect 24912 14980 26249 15008
rect 24912 14968 24918 14980
rect 26237 14977 26249 14980
rect 26283 14977 26295 15011
rect 26237 14971 26295 14977
rect 27341 15011 27399 15017
rect 27341 14977 27353 15011
rect 27387 14977 27399 15011
rect 29454 15008 29460 15020
rect 29415 14980 29460 15008
rect 27341 14971 27399 14977
rect 29454 14968 29460 14980
rect 29512 14968 29518 15020
rect 14274 14900 14280 14952
rect 14332 14940 14338 14952
rect 14737 14943 14795 14949
rect 14737 14940 14749 14943
rect 14332 14912 14749 14940
rect 14332 14900 14338 14912
rect 14737 14909 14749 14912
rect 14783 14909 14795 14943
rect 19426 14940 19432 14952
rect 14737 14903 14795 14909
rect 16132 14912 19432 14940
rect 13556 14844 14596 14872
rect 1581 14807 1639 14813
rect 1581 14773 1593 14807
rect 1627 14804 1639 14807
rect 5074 14804 5080 14816
rect 1627 14776 5080 14804
rect 1627 14773 1639 14776
rect 1581 14767 1639 14773
rect 5074 14764 5080 14776
rect 5132 14764 5138 14816
rect 5350 14764 5356 14816
rect 5408 14804 5414 14816
rect 5626 14804 5632 14816
rect 5408 14776 5632 14804
rect 5408 14764 5414 14776
rect 5626 14764 5632 14776
rect 5684 14764 5690 14816
rect 10505 14807 10563 14813
rect 10505 14773 10517 14807
rect 10551 14804 10563 14807
rect 13814 14804 13820 14816
rect 10551 14776 13820 14804
rect 10551 14773 10563 14776
rect 10505 14767 10563 14773
rect 13814 14764 13820 14776
rect 13872 14764 13878 14816
rect 14568 14804 14596 14844
rect 16132 14804 16160 14912
rect 19426 14900 19432 14912
rect 19484 14900 19490 14952
rect 20162 14940 20168 14952
rect 20123 14912 20168 14940
rect 20162 14900 20168 14912
rect 20220 14900 20226 14952
rect 28813 14943 28871 14949
rect 28813 14909 28825 14943
rect 28859 14940 28871 14943
rect 28994 14940 29000 14952
rect 28859 14912 29000 14940
rect 28859 14909 28871 14912
rect 28813 14903 28871 14909
rect 28994 14900 29000 14912
rect 29052 14900 29058 14952
rect 16206 14832 16212 14884
rect 16264 14872 16270 14884
rect 16264 14844 16309 14872
rect 16264 14832 16270 14844
rect 19518 14832 19524 14884
rect 19576 14872 19582 14884
rect 25314 14872 25320 14884
rect 19576 14844 25320 14872
rect 19576 14832 19582 14844
rect 25314 14832 25320 14844
rect 25372 14832 25378 14884
rect 14568 14776 16160 14804
rect 18138 14764 18144 14816
rect 18196 14804 18202 14816
rect 18398 14807 18456 14813
rect 18398 14804 18410 14807
rect 18196 14776 18410 14804
rect 18196 14764 18202 14776
rect 18398 14773 18410 14776
rect 18444 14773 18456 14807
rect 18398 14767 18456 14773
rect 18506 14764 18512 14816
rect 18564 14804 18570 14816
rect 22373 14807 22431 14813
rect 22373 14804 22385 14807
rect 18564 14776 22385 14804
rect 18564 14764 18570 14776
rect 22373 14773 22385 14776
rect 22419 14773 22431 14807
rect 22373 14767 22431 14773
rect 25222 14764 25228 14816
rect 25280 14804 25286 14816
rect 27157 14807 27215 14813
rect 27157 14804 27169 14807
rect 25280 14776 27169 14804
rect 25280 14764 25286 14776
rect 27157 14773 27169 14776
rect 27203 14773 27215 14807
rect 27157 14767 27215 14773
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 5626 14560 5632 14612
rect 5684 14600 5690 14612
rect 5902 14600 5908 14612
rect 5684 14572 5908 14600
rect 5684 14560 5690 14572
rect 5902 14560 5908 14572
rect 5960 14560 5966 14612
rect 11057 14603 11115 14609
rect 11057 14569 11069 14603
rect 11103 14600 11115 14603
rect 11146 14600 11152 14612
rect 11103 14572 11152 14600
rect 11103 14569 11115 14572
rect 11057 14563 11115 14569
rect 11146 14560 11152 14572
rect 11204 14560 11210 14612
rect 12434 14560 12440 14612
rect 12492 14600 12498 14612
rect 12618 14600 12624 14612
rect 12492 14572 12624 14600
rect 12492 14560 12498 14572
rect 12618 14560 12624 14572
rect 12676 14560 12682 14612
rect 13446 14560 13452 14612
rect 13504 14600 13510 14612
rect 13504 14572 17172 14600
rect 13504 14560 13510 14572
rect 17144 14532 17172 14572
rect 18138 14560 18144 14612
rect 18196 14600 18202 14612
rect 19518 14600 19524 14612
rect 18196 14572 19524 14600
rect 18196 14560 18202 14572
rect 19518 14560 19524 14572
rect 19576 14560 19582 14612
rect 19978 14560 19984 14612
rect 20036 14600 20042 14612
rect 22281 14603 22339 14609
rect 22281 14600 22293 14603
rect 20036 14572 22293 14600
rect 20036 14560 20042 14572
rect 22281 14569 22293 14572
rect 22327 14569 22339 14603
rect 22281 14563 22339 14569
rect 23477 14603 23535 14609
rect 23477 14569 23489 14603
rect 23523 14600 23535 14603
rect 23750 14600 23756 14612
rect 23523 14572 23756 14600
rect 23523 14569 23535 14572
rect 23477 14563 23535 14569
rect 23750 14560 23756 14572
rect 23808 14560 23814 14612
rect 26789 14603 26847 14609
rect 26789 14569 26801 14603
rect 26835 14600 26847 14603
rect 27522 14600 27528 14612
rect 26835 14572 27528 14600
rect 26835 14569 26847 14572
rect 26789 14563 26847 14569
rect 27522 14560 27528 14572
rect 27580 14560 27586 14612
rect 28261 14603 28319 14609
rect 28261 14569 28273 14603
rect 28307 14600 28319 14603
rect 29454 14600 29460 14612
rect 28307 14572 29460 14600
rect 28307 14569 28319 14572
rect 28261 14563 28319 14569
rect 29454 14560 29460 14572
rect 29512 14560 29518 14612
rect 34606 14560 34612 14612
rect 34664 14600 34670 14612
rect 38105 14603 38163 14609
rect 38105 14600 38117 14603
rect 34664 14572 38117 14600
rect 34664 14560 34670 14572
rect 38105 14569 38117 14572
rect 38151 14569 38163 14603
rect 38105 14563 38163 14569
rect 26418 14532 26424 14544
rect 17144 14504 26424 14532
rect 26418 14492 26424 14504
rect 26476 14532 26482 14544
rect 26476 14504 27016 14532
rect 26476 14492 26482 14504
rect 13722 14424 13728 14476
rect 13780 14464 13786 14476
rect 14458 14464 14464 14476
rect 13780 14436 14464 14464
rect 13780 14424 13786 14436
rect 14458 14424 14464 14436
rect 14516 14464 14522 14476
rect 15841 14467 15899 14473
rect 15841 14464 15853 14467
rect 14516 14436 15853 14464
rect 14516 14424 14522 14436
rect 15841 14433 15853 14436
rect 15887 14464 15899 14467
rect 17862 14464 17868 14476
rect 15887 14436 17868 14464
rect 15887 14433 15899 14436
rect 15841 14427 15899 14433
rect 17862 14424 17868 14436
rect 17920 14424 17926 14476
rect 22462 14464 22468 14476
rect 21100 14436 22468 14464
rect 1949 14399 2007 14405
rect 1949 14365 1961 14399
rect 1995 14396 2007 14399
rect 2866 14396 2872 14408
rect 1995 14368 2872 14396
rect 1995 14365 2007 14368
rect 1949 14359 2007 14365
rect 2866 14356 2872 14368
rect 2924 14356 2930 14408
rect 10318 14356 10324 14408
rect 10376 14396 10382 14408
rect 10965 14399 11023 14405
rect 10965 14396 10977 14399
rect 10376 14368 10977 14396
rect 10376 14356 10382 14368
rect 10965 14365 10977 14368
rect 11011 14365 11023 14399
rect 10965 14359 11023 14365
rect 13354 14356 13360 14408
rect 13412 14396 13418 14408
rect 15746 14396 15752 14408
rect 13412 14368 15752 14396
rect 13412 14356 13418 14368
rect 15746 14356 15752 14368
rect 15804 14356 15810 14408
rect 17494 14356 17500 14408
rect 17552 14396 17558 14408
rect 20438 14396 20444 14408
rect 17552 14368 20444 14396
rect 17552 14356 17558 14368
rect 20438 14356 20444 14368
rect 20496 14356 20502 14408
rect 21100 14405 21128 14436
rect 22462 14424 22468 14436
rect 22520 14424 22526 14476
rect 22830 14464 22836 14476
rect 22791 14436 22836 14464
rect 22830 14424 22836 14436
rect 22888 14424 22894 14476
rect 23017 14467 23075 14473
rect 23017 14433 23029 14467
rect 23063 14464 23075 14467
rect 23658 14464 23664 14476
rect 23063 14436 23664 14464
rect 23063 14433 23075 14436
rect 23017 14427 23075 14433
rect 23658 14424 23664 14436
rect 23716 14424 23722 14476
rect 21085 14399 21143 14405
rect 21085 14365 21097 14399
rect 21131 14365 21143 14399
rect 21085 14359 21143 14365
rect 21818 14356 21824 14408
rect 21876 14396 21882 14408
rect 22189 14399 22247 14405
rect 22189 14396 22201 14399
rect 21876 14368 22201 14396
rect 21876 14356 21882 14368
rect 22189 14365 22201 14368
rect 22235 14365 22247 14399
rect 22848 14396 22876 14424
rect 23198 14396 23204 14408
rect 22848 14368 23204 14396
rect 22189 14359 22247 14365
rect 23198 14356 23204 14368
rect 23256 14356 23262 14408
rect 25038 14356 25044 14408
rect 25096 14396 25102 14408
rect 25225 14399 25283 14405
rect 25225 14396 25237 14399
rect 25096 14368 25237 14396
rect 25096 14356 25102 14368
rect 25225 14365 25237 14368
rect 25271 14396 25283 14399
rect 25590 14396 25596 14408
rect 25271 14368 25596 14396
rect 25271 14365 25283 14368
rect 25225 14359 25283 14365
rect 25590 14356 25596 14368
rect 25648 14356 25654 14408
rect 26988 14405 27016 14504
rect 31297 14467 31355 14473
rect 31297 14433 31309 14467
rect 31343 14464 31355 14467
rect 32858 14464 32864 14476
rect 31343 14436 32864 14464
rect 31343 14433 31355 14436
rect 31297 14427 31355 14433
rect 32858 14424 32864 14436
rect 32916 14424 32922 14476
rect 26973 14399 27031 14405
rect 26973 14365 26985 14399
rect 27019 14365 27031 14399
rect 26973 14359 27031 14365
rect 27798 14356 27804 14408
rect 27856 14396 27862 14408
rect 28445 14399 28503 14405
rect 28445 14396 28457 14399
rect 27856 14368 28457 14396
rect 27856 14356 27862 14368
rect 28445 14365 28457 14368
rect 28491 14365 28503 14399
rect 38286 14396 38292 14408
rect 38247 14368 38292 14396
rect 28445 14359 28503 14365
rect 38286 14356 38292 14368
rect 38344 14356 38350 14408
rect 7466 14288 7472 14340
rect 7524 14328 7530 14340
rect 12250 14328 12256 14340
rect 7524 14300 12256 14328
rect 7524 14288 7530 14300
rect 12250 14288 12256 14300
rect 12308 14288 12314 14340
rect 16117 14331 16175 14337
rect 16117 14297 16129 14331
rect 16163 14297 16175 14331
rect 21910 14328 21916 14340
rect 17342 14300 21916 14328
rect 16117 14291 16175 14297
rect 1486 14220 1492 14272
rect 1544 14260 1550 14272
rect 1765 14263 1823 14269
rect 1765 14260 1777 14263
rect 1544 14232 1777 14260
rect 1544 14220 1550 14232
rect 1765 14229 1777 14232
rect 1811 14229 1823 14263
rect 16132 14260 16160 14291
rect 21910 14288 21916 14300
rect 21968 14288 21974 14340
rect 31389 14331 31447 14337
rect 31389 14297 31401 14331
rect 31435 14328 31447 14331
rect 31754 14328 31760 14340
rect 31435 14300 31760 14328
rect 31435 14297 31447 14300
rect 31389 14291 31447 14297
rect 31754 14288 31760 14300
rect 31812 14288 31818 14340
rect 31938 14328 31944 14340
rect 31899 14300 31944 14328
rect 31938 14288 31944 14300
rect 31996 14288 32002 14340
rect 17126 14260 17132 14272
rect 16132 14232 17132 14260
rect 1765 14223 1823 14229
rect 17126 14220 17132 14232
rect 17184 14220 17190 14272
rect 17586 14260 17592 14272
rect 17547 14232 17592 14260
rect 17586 14220 17592 14232
rect 17644 14220 17650 14272
rect 17770 14220 17776 14272
rect 17828 14260 17834 14272
rect 20162 14260 20168 14272
rect 17828 14232 20168 14260
rect 17828 14220 17834 14232
rect 20162 14220 20168 14232
rect 20220 14220 20226 14272
rect 20622 14220 20628 14272
rect 20680 14260 20686 14272
rect 21177 14263 21235 14269
rect 21177 14260 21189 14263
rect 20680 14232 21189 14260
rect 20680 14220 20686 14232
rect 21177 14229 21189 14232
rect 21223 14229 21235 14263
rect 21177 14223 21235 14229
rect 24026 14220 24032 14272
rect 24084 14260 24090 14272
rect 25317 14263 25375 14269
rect 25317 14260 25329 14263
rect 24084 14232 25329 14260
rect 24084 14220 24090 14232
rect 25317 14229 25329 14232
rect 25363 14229 25375 14263
rect 25317 14223 25375 14229
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 1578 14016 1584 14068
rect 1636 14056 1642 14068
rect 1765 14059 1823 14065
rect 1765 14056 1777 14059
rect 1636 14028 1777 14056
rect 1636 14016 1642 14028
rect 1765 14025 1777 14028
rect 1811 14025 1823 14059
rect 1765 14019 1823 14025
rect 2501 14059 2559 14065
rect 2501 14025 2513 14059
rect 2547 14056 2559 14059
rect 3418 14056 3424 14068
rect 2547 14028 3424 14056
rect 2547 14025 2559 14028
rect 2501 14019 2559 14025
rect 3418 14016 3424 14028
rect 3476 14016 3482 14068
rect 8754 14056 8760 14068
rect 7668 14028 8760 14056
rect 5166 13988 5172 14000
rect 5014 13960 5172 13988
rect 5166 13948 5172 13960
rect 5224 13948 5230 14000
rect 5537 13991 5595 13997
rect 5537 13957 5549 13991
rect 5583 13988 5595 13991
rect 5902 13988 5908 14000
rect 5583 13960 5908 13988
rect 5583 13957 5595 13960
rect 5537 13951 5595 13957
rect 5902 13948 5908 13960
rect 5960 13988 5966 14000
rect 6178 13988 6184 14000
rect 5960 13960 6184 13988
rect 5960 13948 5966 13960
rect 6178 13948 6184 13960
rect 6236 13948 6242 14000
rect 1946 13920 1952 13932
rect 1907 13892 1952 13920
rect 1946 13880 1952 13892
rect 2004 13880 2010 13932
rect 2406 13920 2412 13932
rect 2367 13892 2412 13920
rect 2406 13880 2412 13892
rect 2464 13880 2470 13932
rect 7668 13929 7696 14028
rect 8754 14016 8760 14028
rect 8812 14016 8818 14068
rect 20714 14056 20720 14068
rect 12406 14028 20720 14056
rect 12406 13988 12434 14028
rect 20714 14016 20720 14028
rect 20772 14016 20778 14068
rect 20806 14016 20812 14068
rect 20864 14056 20870 14068
rect 22097 14059 22155 14065
rect 22097 14056 22109 14059
rect 20864 14028 22109 14056
rect 20864 14016 20870 14028
rect 22097 14025 22109 14028
rect 22143 14025 22155 14059
rect 22097 14019 22155 14025
rect 23750 14016 23756 14068
rect 23808 14056 23814 14068
rect 24489 14059 24547 14065
rect 24489 14056 24501 14059
rect 23808 14028 24501 14056
rect 23808 14016 23814 14028
rect 24489 14025 24501 14028
rect 24535 14025 24547 14059
rect 24489 14019 24547 14025
rect 25498 14016 25504 14068
rect 25556 14056 25562 14068
rect 25685 14059 25743 14065
rect 25685 14056 25697 14059
rect 25556 14028 25697 14056
rect 25556 14016 25562 14028
rect 25685 14025 25697 14028
rect 25731 14025 25743 14059
rect 31018 14056 31024 14068
rect 30979 14028 31024 14056
rect 25685 14019 25743 14025
rect 31018 14016 31024 14028
rect 31076 14016 31082 14068
rect 13722 13988 13728 14000
rect 9154 13960 12434 13988
rect 13556 13960 13728 13988
rect 13556 13929 13584 13960
rect 13722 13948 13728 13960
rect 13780 13948 13786 14000
rect 18506 13988 18512 14000
rect 15042 13960 18512 13988
rect 18506 13948 18512 13960
rect 18564 13948 18570 14000
rect 20622 13988 20628 14000
rect 19826 13960 20628 13988
rect 20622 13948 20628 13960
rect 20680 13948 20686 14000
rect 27706 13988 27712 14000
rect 21008 13960 21496 13988
rect 7653 13923 7711 13929
rect 7653 13889 7665 13923
rect 7699 13889 7711 13923
rect 7653 13883 7711 13889
rect 13541 13923 13599 13929
rect 13541 13889 13553 13923
rect 13587 13889 13599 13923
rect 13541 13883 13599 13889
rect 15746 13880 15752 13932
rect 15804 13920 15810 13932
rect 17770 13920 17776 13932
rect 15804 13892 17776 13920
rect 15804 13880 15810 13892
rect 17770 13880 17776 13892
rect 17828 13880 17834 13932
rect 17862 13880 17868 13932
rect 17920 13920 17926 13932
rect 18325 13923 18383 13929
rect 18325 13920 18337 13923
rect 17920 13892 18337 13920
rect 17920 13880 17926 13892
rect 18325 13889 18337 13892
rect 18371 13889 18383 13923
rect 20346 13920 20352 13932
rect 20307 13892 20352 13920
rect 18325 13883 18383 13889
rect 20346 13880 20352 13892
rect 20404 13880 20410 13932
rect 20438 13880 20444 13932
rect 20496 13920 20502 13932
rect 21008 13920 21036 13960
rect 20496 13892 21036 13920
rect 21177 13923 21235 13929
rect 20496 13880 20502 13892
rect 21177 13889 21189 13923
rect 21223 13889 21235 13923
rect 21177 13883 21235 13889
rect 3510 13852 3516 13864
rect 3423 13824 3516 13852
rect 3510 13812 3516 13824
rect 3568 13812 3574 13864
rect 3786 13852 3792 13864
rect 3747 13824 3792 13852
rect 3786 13812 3792 13824
rect 3844 13812 3850 13864
rect 9677 13855 9735 13861
rect 9677 13821 9689 13855
rect 9723 13852 9735 13855
rect 13170 13852 13176 13864
rect 9723 13824 13176 13852
rect 9723 13821 9735 13824
rect 9677 13815 9735 13821
rect 13170 13812 13176 13824
rect 13228 13852 13234 13864
rect 13446 13852 13452 13864
rect 13228 13824 13452 13852
rect 13228 13812 13234 13824
rect 13446 13812 13452 13824
rect 13504 13812 13510 13864
rect 15289 13855 15347 13861
rect 13648 13824 14872 13852
rect 3528 13716 3556 13812
rect 11422 13784 11428 13796
rect 10060 13756 11428 13784
rect 3970 13716 3976 13728
rect 3528 13688 3976 13716
rect 3970 13676 3976 13688
rect 4028 13676 4034 13728
rect 7916 13719 7974 13725
rect 7916 13685 7928 13719
rect 7962 13716 7974 13719
rect 10060 13716 10088 13756
rect 11422 13744 11428 13756
rect 11480 13744 11486 13796
rect 13538 13744 13544 13796
rect 13596 13784 13602 13796
rect 13648 13784 13676 13824
rect 13596 13756 13676 13784
rect 14844 13784 14872 13824
rect 15289 13821 15301 13855
rect 15335 13852 15347 13855
rect 17954 13852 17960 13864
rect 15335 13824 17960 13852
rect 15335 13821 15347 13824
rect 15289 13815 15347 13821
rect 17954 13812 17960 13824
rect 18012 13812 18018 13864
rect 18601 13855 18659 13861
rect 18601 13852 18613 13855
rect 18432 13824 18613 13852
rect 14844 13756 15424 13784
rect 13596 13744 13602 13756
rect 7962 13688 10088 13716
rect 7962 13685 7974 13688
rect 7916 13679 7974 13685
rect 10134 13676 10140 13728
rect 10192 13716 10198 13728
rect 13630 13716 13636 13728
rect 10192 13688 13636 13716
rect 10192 13676 10198 13688
rect 13630 13676 13636 13688
rect 13688 13676 13694 13728
rect 13804 13719 13862 13725
rect 13804 13685 13816 13719
rect 13850 13716 13862 13719
rect 13998 13716 14004 13728
rect 13850 13688 14004 13716
rect 13850 13685 13862 13688
rect 13804 13679 13862 13685
rect 13998 13676 14004 13688
rect 14056 13716 14062 13728
rect 15010 13716 15016 13728
rect 14056 13688 15016 13716
rect 14056 13676 14062 13688
rect 15010 13676 15016 13688
rect 15068 13676 15074 13728
rect 15396 13716 15424 13756
rect 17586 13744 17592 13796
rect 17644 13784 17650 13796
rect 18432 13784 18460 13824
rect 18601 13821 18613 13824
rect 18647 13852 18659 13855
rect 18647 13824 19656 13852
rect 18647 13821 18659 13824
rect 18601 13815 18659 13821
rect 17644 13756 18460 13784
rect 19628 13784 19656 13824
rect 20990 13784 20996 13796
rect 19628 13756 20996 13784
rect 17644 13744 17650 13756
rect 20990 13744 20996 13756
rect 21048 13744 21054 13796
rect 19058 13716 19064 13728
rect 15396 13688 19064 13716
rect 19058 13676 19064 13688
rect 19116 13676 19122 13728
rect 21192 13716 21220 13883
rect 21358 13852 21364 13864
rect 21284 13824 21364 13852
rect 21284 13793 21312 13824
rect 21358 13812 21364 13824
rect 21416 13812 21422 13864
rect 21468 13852 21496 13960
rect 23860 13960 27712 13988
rect 21726 13880 21732 13932
rect 21784 13920 21790 13932
rect 22005 13923 22063 13929
rect 22005 13920 22017 13923
rect 21784 13892 22017 13920
rect 21784 13880 21790 13892
rect 22005 13889 22017 13892
rect 22051 13889 22063 13923
rect 22005 13883 22063 13889
rect 22649 13923 22707 13929
rect 22649 13889 22661 13923
rect 22695 13920 22707 13923
rect 22738 13920 22744 13932
rect 22695 13892 22744 13920
rect 22695 13889 22707 13892
rect 22649 13883 22707 13889
rect 22738 13880 22744 13892
rect 22796 13880 22802 13932
rect 23860 13929 23888 13960
rect 23845 13923 23903 13929
rect 23845 13889 23857 13923
rect 23891 13889 23903 13923
rect 24026 13920 24032 13932
rect 23987 13892 24032 13920
rect 23845 13883 23903 13889
rect 24026 13880 24032 13892
rect 24084 13880 24090 13932
rect 25222 13920 25228 13932
rect 25183 13892 25228 13920
rect 25222 13880 25228 13892
rect 25280 13880 25286 13932
rect 27172 13929 27200 13960
rect 27706 13948 27712 13960
rect 27764 13948 27770 14000
rect 28442 13988 28448 14000
rect 28403 13960 28448 13988
rect 28442 13948 28448 13960
rect 28500 13948 28506 14000
rect 27157 13923 27215 13929
rect 27157 13889 27169 13923
rect 27203 13889 27215 13923
rect 27338 13920 27344 13932
rect 27299 13892 27344 13920
rect 27157 13883 27215 13889
rect 27338 13880 27344 13892
rect 27396 13880 27402 13932
rect 30929 13923 30987 13929
rect 30929 13889 30941 13923
rect 30975 13920 30987 13923
rect 38102 13920 38108 13932
rect 30975 13892 38108 13920
rect 30975 13889 30987 13892
rect 30929 13883 30987 13889
rect 38102 13880 38108 13892
rect 38160 13880 38166 13932
rect 25038 13852 25044 13864
rect 21468 13824 24900 13852
rect 24999 13824 25044 13852
rect 21269 13787 21327 13793
rect 21269 13753 21281 13787
rect 21315 13753 21327 13787
rect 24872 13784 24900 13824
rect 25038 13812 25044 13824
rect 25096 13812 25102 13864
rect 27062 13852 27068 13864
rect 25148 13824 27068 13852
rect 25148 13784 25176 13824
rect 27062 13812 27068 13824
rect 27120 13812 27126 13864
rect 27801 13855 27859 13861
rect 27801 13821 27813 13855
rect 27847 13852 27859 13855
rect 28350 13852 28356 13864
rect 27847 13824 28356 13852
rect 27847 13821 27859 13824
rect 27801 13815 27859 13821
rect 28350 13812 28356 13824
rect 28408 13812 28414 13864
rect 28813 13855 28871 13861
rect 28813 13821 28825 13855
rect 28859 13852 28871 13855
rect 28994 13852 29000 13864
rect 28859 13824 29000 13852
rect 28859 13821 28871 13824
rect 28813 13815 28871 13821
rect 28994 13812 29000 13824
rect 29052 13852 29058 13864
rect 30190 13852 30196 13864
rect 29052 13824 30196 13852
rect 29052 13812 29058 13824
rect 30190 13812 30196 13824
rect 30248 13812 30254 13864
rect 24872 13756 25176 13784
rect 21269 13747 21327 13753
rect 21358 13716 21364 13728
rect 21192 13688 21364 13716
rect 21358 13676 21364 13688
rect 21416 13676 21422 13728
rect 21450 13676 21456 13728
rect 21508 13716 21514 13728
rect 22741 13719 22799 13725
rect 22741 13716 22753 13719
rect 21508 13688 22753 13716
rect 21508 13676 21514 13688
rect 22741 13685 22753 13688
rect 22787 13685 22799 13719
rect 22741 13679 22799 13685
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 4890 13472 4896 13524
rect 4948 13512 4954 13524
rect 5721 13515 5779 13521
rect 4948 13484 5672 13512
rect 4948 13472 4954 13484
rect 5644 13444 5672 13484
rect 5721 13481 5733 13515
rect 5767 13512 5779 13515
rect 6730 13512 6736 13524
rect 5767 13484 6736 13512
rect 5767 13481 5779 13484
rect 5721 13475 5779 13481
rect 6730 13472 6736 13484
rect 6788 13472 6794 13524
rect 13538 13512 13544 13524
rect 8680 13484 13544 13512
rect 8680 13444 8708 13484
rect 13538 13472 13544 13484
rect 13596 13472 13602 13524
rect 13814 13472 13820 13524
rect 13872 13512 13878 13524
rect 14550 13521 14556 13524
rect 14534 13515 14556 13521
rect 14534 13512 14546 13515
rect 13872 13484 14546 13512
rect 13872 13472 13878 13484
rect 14534 13481 14546 13484
rect 14608 13512 14614 13524
rect 14608 13484 14682 13512
rect 14534 13475 14556 13481
rect 14550 13472 14556 13475
rect 14608 13472 14614 13484
rect 15654 13472 15660 13524
rect 15712 13512 15718 13524
rect 20990 13512 20996 13524
rect 15712 13484 20996 13512
rect 15712 13472 15718 13484
rect 20990 13472 20996 13484
rect 21048 13472 21054 13524
rect 21928 13484 26648 13512
rect 5644 13416 8708 13444
rect 12710 13404 12716 13456
rect 12768 13444 12774 13456
rect 12768 13416 14412 13444
rect 12768 13404 12774 13416
rect 1949 13379 2007 13385
rect 1949 13345 1961 13379
rect 1995 13376 2007 13379
rect 3878 13376 3884 13388
rect 1995 13348 3884 13376
rect 1995 13345 2007 13348
rect 1949 13339 2007 13345
rect 3878 13336 3884 13348
rect 3936 13336 3942 13388
rect 4249 13379 4307 13385
rect 4249 13345 4261 13379
rect 4295 13376 4307 13379
rect 10134 13376 10140 13388
rect 4295 13348 10140 13376
rect 4295 13345 4307 13348
rect 4249 13339 4307 13345
rect 10134 13336 10140 13348
rect 10192 13336 10198 13388
rect 11057 13379 11115 13385
rect 11057 13345 11069 13379
rect 11103 13376 11115 13379
rect 12066 13376 12072 13388
rect 11103 13348 12072 13376
rect 11103 13345 11115 13348
rect 11057 13339 11115 13345
rect 12066 13336 12072 13348
rect 12124 13376 12130 13388
rect 13722 13376 13728 13388
rect 12124 13348 13728 13376
rect 12124 13336 12130 13348
rect 13722 13336 13728 13348
rect 13780 13376 13786 13388
rect 14277 13379 14335 13385
rect 14277 13376 14289 13379
rect 13780 13348 14289 13376
rect 13780 13336 13786 13348
rect 14277 13345 14289 13348
rect 14323 13345 14335 13379
rect 14384 13376 14412 13416
rect 15562 13404 15568 13456
rect 15620 13444 15626 13456
rect 21928 13444 21956 13484
rect 15620 13416 21956 13444
rect 15620 13404 15626 13416
rect 26234 13404 26240 13456
rect 26292 13444 26298 13456
rect 26513 13447 26571 13453
rect 26513 13444 26525 13447
rect 26292 13416 26525 13444
rect 26292 13404 26298 13416
rect 26513 13413 26525 13416
rect 26559 13413 26571 13447
rect 26620 13444 26648 13484
rect 28534 13472 28540 13524
rect 28592 13512 28598 13524
rect 28721 13515 28779 13521
rect 28721 13512 28733 13515
rect 28592 13484 28733 13512
rect 28592 13472 28598 13484
rect 28721 13481 28733 13484
rect 28767 13481 28779 13515
rect 28721 13475 28779 13481
rect 31754 13472 31760 13524
rect 31812 13512 31818 13524
rect 31941 13515 31999 13521
rect 31941 13512 31953 13515
rect 31812 13484 31953 13512
rect 31812 13472 31818 13484
rect 31941 13481 31953 13484
rect 31987 13481 31999 13515
rect 31941 13475 31999 13481
rect 29178 13444 29184 13456
rect 26620 13416 29184 13444
rect 26513 13407 26571 13413
rect 29178 13404 29184 13416
rect 29236 13404 29242 13456
rect 30466 13404 30472 13456
rect 30524 13444 30530 13456
rect 31113 13447 31171 13453
rect 31113 13444 31125 13447
rect 30524 13416 31125 13444
rect 30524 13404 30530 13416
rect 31113 13413 31125 13416
rect 31159 13444 31171 13447
rect 31202 13444 31208 13456
rect 31159 13416 31208 13444
rect 31159 13413 31171 13416
rect 31113 13407 31171 13413
rect 31202 13404 31208 13416
rect 31260 13404 31266 13456
rect 21450 13376 21456 13388
rect 14384 13348 21456 13376
rect 14277 13339 14335 13345
rect 21450 13336 21456 13348
rect 21508 13336 21514 13388
rect 21542 13336 21548 13388
rect 21600 13376 21606 13388
rect 21821 13379 21879 13385
rect 21821 13376 21833 13379
rect 21600 13348 21833 13376
rect 21600 13336 21606 13348
rect 21821 13345 21833 13348
rect 21867 13345 21879 13379
rect 21821 13339 21879 13345
rect 25038 13336 25044 13388
rect 25096 13376 25102 13388
rect 25133 13379 25191 13385
rect 25133 13376 25145 13379
rect 25096 13348 25145 13376
rect 25096 13336 25102 13348
rect 25133 13345 25145 13348
rect 25179 13345 25191 13379
rect 25133 13339 25191 13345
rect 26145 13379 26203 13385
rect 26145 13345 26157 13379
rect 26191 13376 26203 13379
rect 30561 13379 30619 13385
rect 30561 13376 30573 13379
rect 26191 13348 30573 13376
rect 26191 13345 26203 13348
rect 26145 13339 26203 13345
rect 30561 13345 30573 13348
rect 30607 13376 30619 13379
rect 31846 13376 31852 13388
rect 30607 13348 31852 13376
rect 30607 13345 30619 13348
rect 30561 13339 30619 13345
rect 31846 13336 31852 13348
rect 31904 13336 31910 13388
rect 1578 13268 1584 13320
rect 1636 13308 1642 13320
rect 1857 13311 1915 13317
rect 1857 13308 1869 13311
rect 1636 13280 1869 13308
rect 1636 13268 1642 13280
rect 1857 13277 1869 13280
rect 1903 13277 1915 13311
rect 3970 13308 3976 13320
rect 3931 13280 3976 13308
rect 1857 13271 1915 13277
rect 3970 13268 3976 13280
rect 4028 13268 4034 13320
rect 7742 13268 7748 13320
rect 7800 13308 7806 13320
rect 9122 13308 9128 13320
rect 7800 13280 9128 13308
rect 7800 13268 7806 13280
rect 9122 13268 9128 13280
rect 9180 13268 9186 13320
rect 12618 13268 12624 13320
rect 12676 13308 12682 13320
rect 14182 13308 14188 13320
rect 12676 13280 14188 13308
rect 12676 13268 12682 13280
rect 14182 13268 14188 13280
rect 14240 13268 14246 13320
rect 18690 13308 18696 13320
rect 15686 13280 18696 13308
rect 18690 13268 18696 13280
rect 18748 13268 18754 13320
rect 21085 13311 21143 13317
rect 21085 13277 21097 13311
rect 21131 13308 21143 13311
rect 21358 13308 21364 13320
rect 21131 13280 21364 13308
rect 21131 13277 21143 13280
rect 21085 13271 21143 13277
rect 21358 13268 21364 13280
rect 21416 13308 21422 13320
rect 21729 13311 21787 13317
rect 21729 13308 21741 13311
rect 21416 13280 21741 13308
rect 21416 13268 21422 13280
rect 21729 13277 21741 13280
rect 21775 13308 21787 13311
rect 21775 13280 21864 13308
rect 21775 13277 21787 13280
rect 21729 13271 21787 13277
rect 5474 13212 9352 13240
rect 6454 13132 6460 13184
rect 6512 13172 6518 13184
rect 9217 13175 9275 13181
rect 9217 13172 9229 13175
rect 6512 13144 9229 13172
rect 6512 13132 6518 13144
rect 9217 13141 9229 13144
rect 9263 13141 9275 13175
rect 9324 13172 9352 13212
rect 10778 13200 10784 13252
rect 10836 13240 10842 13252
rect 11333 13243 11391 13249
rect 11333 13240 11345 13243
rect 10836 13212 11345 13240
rect 10836 13200 10842 13212
rect 11333 13209 11345 13212
rect 11379 13209 11391 13243
rect 21542 13240 21548 13252
rect 12558 13212 14964 13240
rect 11333 13203 11391 13209
rect 12710 13172 12716 13184
rect 9324 13144 12716 13172
rect 9217 13135 9275 13141
rect 12710 13132 12716 13144
rect 12768 13132 12774 13184
rect 12805 13175 12863 13181
rect 12805 13141 12817 13175
rect 12851 13172 12863 13175
rect 12894 13172 12900 13184
rect 12851 13144 12900 13172
rect 12851 13141 12863 13144
rect 12805 13135 12863 13141
rect 12894 13132 12900 13144
rect 12952 13132 12958 13184
rect 14936 13172 14964 13212
rect 15856 13212 21548 13240
rect 15856 13172 15884 13212
rect 21542 13200 21548 13212
rect 21600 13200 21606 13252
rect 21836 13240 21864 13280
rect 22002 13268 22008 13320
rect 22060 13308 22066 13320
rect 22373 13311 22431 13317
rect 22373 13308 22385 13311
rect 22060 13280 22385 13308
rect 22060 13268 22066 13280
rect 22373 13277 22385 13280
rect 22419 13277 22431 13311
rect 22373 13271 22431 13277
rect 26329 13311 26387 13317
rect 26329 13277 26341 13311
rect 26375 13308 26387 13311
rect 27430 13308 27436 13320
rect 26375 13280 27436 13308
rect 26375 13277 26387 13280
rect 26329 13271 26387 13277
rect 27430 13268 27436 13280
rect 27488 13268 27494 13320
rect 28905 13311 28963 13317
rect 28905 13277 28917 13311
rect 28951 13308 28963 13311
rect 29638 13308 29644 13320
rect 28951 13280 29644 13308
rect 28951 13277 28963 13280
rect 28905 13271 28963 13277
rect 29638 13268 29644 13280
rect 29696 13268 29702 13320
rect 29914 13308 29920 13320
rect 29875 13280 29920 13308
rect 29914 13268 29920 13280
rect 29972 13268 29978 13320
rect 32122 13308 32128 13320
rect 32083 13280 32128 13308
rect 32122 13268 32128 13280
rect 32180 13268 32186 13320
rect 22738 13240 22744 13252
rect 21836 13212 22744 13240
rect 22738 13200 22744 13212
rect 22796 13200 22802 13252
rect 30650 13200 30656 13252
rect 30708 13240 30714 13252
rect 30708 13212 30753 13240
rect 30708 13200 30714 13212
rect 16022 13172 16028 13184
rect 14936 13144 15884 13172
rect 15983 13144 16028 13172
rect 16022 13132 16028 13144
rect 16080 13132 16086 13184
rect 17494 13132 17500 13184
rect 17552 13172 17558 13184
rect 19242 13172 19248 13184
rect 17552 13144 19248 13172
rect 17552 13132 17558 13144
rect 19242 13132 19248 13144
rect 19300 13132 19306 13184
rect 19334 13132 19340 13184
rect 19392 13172 19398 13184
rect 21177 13175 21235 13181
rect 21177 13172 21189 13175
rect 19392 13144 21189 13172
rect 19392 13132 19398 13144
rect 21177 13141 21189 13144
rect 21223 13141 21235 13175
rect 21177 13135 21235 13141
rect 21634 13132 21640 13184
rect 21692 13172 21698 13184
rect 21910 13172 21916 13184
rect 21692 13144 21916 13172
rect 21692 13132 21698 13144
rect 21910 13132 21916 13144
rect 21968 13132 21974 13184
rect 22002 13132 22008 13184
rect 22060 13172 22066 13184
rect 22465 13175 22523 13181
rect 22465 13172 22477 13175
rect 22060 13144 22477 13172
rect 22060 13132 22066 13144
rect 22465 13141 22477 13144
rect 22511 13141 22523 13175
rect 22465 13135 22523 13141
rect 29733 13175 29791 13181
rect 29733 13141 29745 13175
rect 29779 13172 29791 13175
rect 30926 13172 30932 13184
rect 29779 13144 30932 13172
rect 29779 13141 29791 13144
rect 29733 13135 29791 13141
rect 30926 13132 30932 13144
rect 30984 13132 30990 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 1578 12968 1584 12980
rect 1539 12940 1584 12968
rect 1578 12928 1584 12940
rect 1636 12928 1642 12980
rect 3786 12928 3792 12980
rect 3844 12968 3850 12980
rect 3844 12940 10272 12968
rect 3844 12928 3850 12940
rect 6822 12900 6828 12912
rect 6783 12872 6828 12900
rect 6822 12860 6828 12872
rect 6880 12860 6886 12912
rect 7374 12900 7380 12912
rect 7335 12872 7380 12900
rect 7374 12860 7380 12872
rect 7432 12860 7438 12912
rect 9398 12860 9404 12912
rect 9456 12860 9462 12912
rect 10244 12900 10272 12940
rect 12158 12928 12164 12980
rect 12216 12968 12222 12980
rect 12894 12968 12900 12980
rect 12216 12940 12900 12968
rect 12216 12928 12222 12940
rect 12894 12928 12900 12940
rect 12952 12968 12958 12980
rect 12952 12940 15792 12968
rect 12952 12928 12958 12940
rect 12618 12900 12624 12912
rect 10244 12872 12624 12900
rect 12618 12860 12624 12872
rect 12676 12860 12682 12912
rect 14274 12900 14280 12912
rect 14235 12872 14280 12900
rect 14274 12860 14280 12872
rect 14332 12860 14338 12912
rect 1762 12832 1768 12844
rect 1723 12804 1768 12832
rect 1762 12792 1768 12804
rect 1820 12792 1826 12844
rect 8662 12832 8668 12844
rect 8623 12804 8668 12832
rect 8662 12792 8668 12804
rect 8720 12792 8726 12844
rect 10226 12792 10232 12844
rect 10284 12832 10290 12844
rect 10594 12832 10600 12844
rect 10284 12804 10600 12832
rect 10284 12792 10290 12804
rect 10594 12792 10600 12804
rect 10652 12832 10658 12844
rect 10689 12835 10747 12841
rect 10689 12832 10701 12835
rect 10652 12804 10701 12832
rect 10652 12792 10658 12804
rect 10689 12801 10701 12804
rect 10735 12801 10747 12835
rect 10689 12795 10747 12801
rect 12066 12792 12072 12844
rect 12124 12832 12130 12844
rect 12253 12835 12311 12841
rect 12253 12832 12265 12835
rect 12124 12804 12265 12832
rect 12124 12792 12130 12804
rect 12253 12801 12265 12804
rect 12299 12801 12311 12835
rect 15654 12832 15660 12844
rect 13662 12804 15660 12832
rect 12253 12795 12311 12801
rect 15654 12792 15660 12804
rect 15712 12792 15718 12844
rect 4614 12724 4620 12776
rect 4672 12764 4678 12776
rect 6733 12767 6791 12773
rect 6733 12764 6745 12767
rect 4672 12736 6745 12764
rect 4672 12724 4678 12736
rect 6733 12733 6745 12736
rect 6779 12733 6791 12767
rect 8941 12767 8999 12773
rect 8941 12764 8953 12767
rect 6733 12727 6791 12733
rect 6840 12736 8953 12764
rect 1854 12656 1860 12708
rect 1912 12696 1918 12708
rect 6840 12696 6868 12736
rect 8941 12733 8953 12736
rect 8987 12733 8999 12767
rect 8941 12727 8999 12733
rect 9030 12724 9036 12776
rect 9088 12764 9094 12776
rect 11054 12764 11060 12776
rect 9088 12736 11060 12764
rect 9088 12724 9094 12736
rect 11054 12724 11060 12736
rect 11112 12724 11118 12776
rect 12529 12767 12587 12773
rect 12529 12764 12541 12767
rect 11900 12736 12541 12764
rect 1912 12668 6868 12696
rect 1912 12656 1918 12668
rect 3878 12588 3884 12640
rect 3936 12628 3942 12640
rect 9030 12628 9036 12640
rect 3936 12600 9036 12628
rect 3936 12588 3942 12600
rect 9030 12588 9036 12600
rect 9088 12588 9094 12640
rect 9122 12588 9128 12640
rect 9180 12628 9186 12640
rect 11606 12628 11612 12640
rect 9180 12600 11612 12628
rect 9180 12588 9186 12600
rect 11606 12588 11612 12600
rect 11664 12588 11670 12640
rect 11698 12588 11704 12640
rect 11756 12628 11762 12640
rect 11900 12637 11928 12736
rect 12529 12733 12541 12736
rect 12575 12764 12587 12767
rect 15562 12764 15568 12776
rect 12575 12736 15568 12764
rect 12575 12733 12587 12736
rect 12529 12727 12587 12733
rect 15562 12724 15568 12736
rect 15620 12724 15626 12776
rect 15764 12764 15792 12940
rect 17862 12928 17868 12980
rect 17920 12928 17926 12980
rect 19150 12968 19156 12980
rect 19111 12940 19156 12968
rect 19150 12928 19156 12940
rect 19208 12928 19214 12980
rect 19242 12928 19248 12980
rect 19300 12968 19306 12980
rect 25225 12971 25283 12977
rect 19300 12940 23520 12968
rect 19300 12928 19306 12940
rect 17880 12900 17908 12928
rect 22097 12903 22155 12909
rect 22097 12900 22109 12903
rect 17420 12872 17908 12900
rect 18906 12872 22109 12900
rect 17310 12792 17316 12844
rect 17368 12832 17374 12844
rect 17420 12841 17448 12872
rect 22097 12869 22109 12872
rect 22143 12869 22155 12903
rect 22097 12863 22155 12869
rect 17405 12835 17463 12841
rect 17405 12832 17417 12835
rect 17368 12804 17417 12832
rect 17368 12792 17374 12804
rect 17405 12801 17417 12804
rect 17451 12801 17463 12835
rect 21082 12832 21088 12844
rect 20995 12804 21088 12832
rect 17405 12795 17463 12801
rect 21082 12792 21088 12804
rect 21140 12832 21146 12844
rect 21726 12832 21732 12844
rect 21140 12804 21732 12832
rect 21140 12792 21146 12804
rect 21726 12792 21732 12804
rect 21784 12792 21790 12844
rect 21818 12792 21824 12844
rect 21876 12832 21882 12844
rect 23492 12841 23520 12940
rect 25225 12937 25237 12971
rect 25271 12968 25283 12971
rect 25498 12968 25504 12980
rect 25271 12940 25504 12968
rect 25271 12937 25283 12940
rect 25225 12931 25283 12937
rect 25498 12928 25504 12940
rect 25556 12928 25562 12980
rect 27893 12971 27951 12977
rect 27893 12937 27905 12971
rect 27939 12968 27951 12971
rect 28442 12968 28448 12980
rect 27939 12940 28448 12968
rect 27939 12937 27951 12940
rect 27893 12931 27951 12937
rect 28442 12928 28448 12940
rect 28500 12928 28506 12980
rect 24121 12903 24179 12909
rect 24121 12869 24133 12903
rect 24167 12900 24179 12903
rect 25406 12900 25412 12912
rect 24167 12872 25412 12900
rect 24167 12869 24179 12872
rect 24121 12863 24179 12869
rect 25406 12860 25412 12872
rect 25464 12860 25470 12912
rect 30926 12900 30932 12912
rect 30887 12872 30932 12900
rect 30926 12860 30932 12872
rect 30984 12860 30990 12912
rect 22005 12835 22063 12841
rect 22005 12832 22017 12835
rect 21876 12804 22017 12832
rect 21876 12792 21882 12804
rect 22005 12801 22017 12804
rect 22051 12801 22063 12835
rect 22005 12795 22063 12801
rect 23477 12835 23535 12841
rect 23477 12801 23489 12835
rect 23523 12801 23535 12835
rect 23477 12795 23535 12801
rect 24581 12835 24639 12841
rect 24581 12801 24593 12835
rect 24627 12832 24639 12835
rect 26602 12832 26608 12844
rect 24627 12804 26608 12832
rect 24627 12801 24639 12804
rect 24581 12795 24639 12801
rect 26602 12792 26608 12804
rect 26660 12792 26666 12844
rect 27798 12832 27804 12844
rect 27759 12804 27804 12832
rect 27798 12792 27804 12804
rect 27856 12792 27862 12844
rect 27890 12792 27896 12844
rect 27948 12832 27954 12844
rect 28629 12835 28687 12841
rect 28629 12832 28641 12835
rect 27948 12804 28641 12832
rect 27948 12792 27954 12804
rect 28629 12801 28641 12804
rect 28675 12801 28687 12835
rect 28629 12795 28687 12801
rect 36722 12792 36728 12844
rect 36780 12832 36786 12844
rect 38013 12835 38071 12841
rect 38013 12832 38025 12835
rect 36780 12804 38025 12832
rect 36780 12792 36786 12804
rect 38013 12801 38025 12804
rect 38059 12801 38071 12835
rect 38013 12795 38071 12801
rect 15764 12736 22508 12764
rect 14182 12656 14188 12708
rect 14240 12696 14246 12708
rect 16206 12696 16212 12708
rect 14240 12668 16212 12696
rect 14240 12656 14246 12668
rect 16206 12656 16212 12668
rect 16264 12656 16270 12708
rect 18690 12656 18696 12708
rect 18748 12696 18754 12708
rect 22186 12696 22192 12708
rect 18748 12668 21312 12696
rect 18748 12656 18754 12668
rect 11885 12631 11943 12637
rect 11885 12628 11897 12631
rect 11756 12600 11897 12628
rect 11756 12588 11762 12600
rect 11885 12597 11897 12600
rect 11931 12597 11943 12631
rect 11885 12591 11943 12597
rect 12618 12588 12624 12640
rect 12676 12628 12682 12640
rect 15378 12628 15384 12640
rect 12676 12600 15384 12628
rect 12676 12588 12682 12600
rect 15378 12588 15384 12600
rect 15436 12588 15442 12640
rect 16482 12588 16488 12640
rect 16540 12628 16546 12640
rect 17662 12631 17720 12637
rect 17662 12628 17674 12631
rect 16540 12600 17674 12628
rect 16540 12588 16546 12600
rect 17662 12597 17674 12600
rect 17708 12597 17720 12631
rect 17662 12591 17720 12597
rect 17770 12588 17776 12640
rect 17828 12628 17834 12640
rect 21177 12631 21235 12637
rect 21177 12628 21189 12631
rect 17828 12600 21189 12628
rect 17828 12588 17834 12600
rect 21177 12597 21189 12600
rect 21223 12597 21235 12631
rect 21284 12628 21312 12668
rect 22066 12668 22192 12696
rect 22066 12628 22094 12668
rect 22186 12656 22192 12668
rect 22244 12656 22250 12708
rect 22480 12696 22508 12736
rect 22554 12724 22560 12776
rect 22612 12764 22618 12776
rect 23661 12767 23719 12773
rect 23661 12764 23673 12767
rect 22612 12736 23673 12764
rect 22612 12724 22618 12736
rect 23661 12733 23673 12736
rect 23707 12733 23719 12767
rect 23661 12727 23719 12733
rect 24765 12767 24823 12773
rect 24765 12733 24777 12767
rect 24811 12764 24823 12767
rect 24946 12764 24952 12776
rect 24811 12736 24952 12764
rect 24811 12733 24823 12736
rect 24765 12727 24823 12733
rect 24946 12724 24952 12736
rect 25004 12724 25010 12776
rect 27908 12696 27936 12792
rect 30834 12764 30840 12776
rect 30795 12736 30840 12764
rect 30834 12724 30840 12736
rect 30892 12724 30898 12776
rect 31110 12764 31116 12776
rect 31071 12736 31116 12764
rect 31110 12724 31116 12736
rect 31168 12764 31174 12776
rect 31294 12764 31300 12776
rect 31168 12736 31300 12764
rect 31168 12724 31174 12736
rect 31294 12724 31300 12736
rect 31352 12724 31358 12776
rect 22480 12668 27936 12696
rect 28445 12699 28503 12705
rect 28445 12665 28457 12699
rect 28491 12696 28503 12699
rect 29914 12696 29920 12708
rect 28491 12668 29920 12696
rect 28491 12665 28503 12668
rect 28445 12659 28503 12665
rect 29914 12656 29920 12668
rect 29972 12656 29978 12708
rect 38194 12628 38200 12640
rect 21284 12600 22094 12628
rect 38155 12600 38200 12628
rect 21177 12591 21235 12597
rect 38194 12588 38200 12600
rect 38252 12588 38258 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 1946 12424 1952 12436
rect 1907 12396 1952 12424
rect 1946 12384 1952 12396
rect 2004 12384 2010 12436
rect 7374 12424 7380 12436
rect 2746 12396 7380 12424
rect 2746 12288 2774 12396
rect 7374 12384 7380 12396
rect 7432 12384 7438 12436
rect 10502 12384 10508 12436
rect 10560 12424 10566 12436
rect 17034 12424 17040 12436
rect 10560 12396 17040 12424
rect 10560 12384 10566 12396
rect 17034 12384 17040 12396
rect 17092 12384 17098 12436
rect 21358 12424 21364 12436
rect 17144 12396 21364 12424
rect 14369 12359 14427 12365
rect 14369 12356 14381 12359
rect 1872 12260 2774 12288
rect 5368 12328 14381 12356
rect 1872 12229 1900 12260
rect 1857 12223 1915 12229
rect 1857 12189 1869 12223
rect 1903 12189 1915 12223
rect 3970 12220 3976 12232
rect 3931 12192 3976 12220
rect 1857 12183 1915 12189
rect 3970 12180 3976 12192
rect 4028 12180 4034 12232
rect 5368 12206 5396 12328
rect 14369 12325 14381 12328
rect 14415 12325 14427 12359
rect 14369 12319 14427 12325
rect 5626 12248 5632 12300
rect 5684 12288 5690 12300
rect 6362 12288 6368 12300
rect 5684 12260 6368 12288
rect 5684 12248 5690 12260
rect 6362 12248 6368 12260
rect 6420 12288 6426 12300
rect 9214 12288 9220 12300
rect 6420 12260 9220 12288
rect 6420 12248 6426 12260
rect 9214 12248 9220 12260
rect 9272 12248 9278 12300
rect 11054 12248 11060 12300
rect 11112 12288 11118 12300
rect 11793 12291 11851 12297
rect 11793 12288 11805 12291
rect 11112 12260 11805 12288
rect 11112 12248 11118 12260
rect 11793 12257 11805 12260
rect 11839 12257 11851 12291
rect 12250 12288 12256 12300
rect 12211 12260 12256 12288
rect 11793 12251 11851 12257
rect 12250 12248 12256 12260
rect 12308 12248 12314 12300
rect 17144 12288 17172 12396
rect 21358 12384 21364 12396
rect 21416 12384 21422 12436
rect 24946 12424 24952 12436
rect 24907 12396 24952 12424
rect 24946 12384 24952 12396
rect 25004 12384 25010 12436
rect 30377 12427 30435 12433
rect 30377 12393 30389 12427
rect 30423 12424 30435 12427
rect 30650 12424 30656 12436
rect 30423 12396 30656 12424
rect 30423 12393 30435 12396
rect 30377 12387 30435 12393
rect 30650 12384 30656 12396
rect 30708 12384 30714 12436
rect 31665 12427 31723 12433
rect 31665 12393 31677 12427
rect 31711 12424 31723 12427
rect 32122 12424 32128 12436
rect 31711 12396 32128 12424
rect 31711 12393 31723 12396
rect 31665 12387 31723 12393
rect 32122 12384 32128 12396
rect 32180 12384 32186 12436
rect 35805 12427 35863 12433
rect 35805 12393 35817 12427
rect 35851 12424 35863 12427
rect 36722 12424 36728 12436
rect 35851 12396 36728 12424
rect 35851 12393 35863 12396
rect 35805 12387 35863 12393
rect 36722 12384 36728 12396
rect 36780 12384 36786 12436
rect 17218 12316 17224 12368
rect 17276 12356 17282 12368
rect 23290 12356 23296 12368
rect 17276 12328 23296 12356
rect 17276 12316 17282 12328
rect 23290 12316 23296 12328
rect 23348 12316 23354 12368
rect 26326 12356 26332 12368
rect 26287 12328 26332 12356
rect 26326 12316 26332 12328
rect 26384 12316 26390 12368
rect 27062 12316 27068 12368
rect 27120 12356 27126 12368
rect 28261 12359 28319 12365
rect 28261 12356 28273 12359
rect 27120 12328 28273 12356
rect 27120 12316 27126 12328
rect 28261 12325 28273 12328
rect 28307 12356 28319 12359
rect 31938 12356 31944 12368
rect 28307 12328 31944 12356
rect 28307 12325 28319 12328
rect 28261 12319 28319 12325
rect 31938 12316 31944 12328
rect 31996 12316 32002 12368
rect 14292 12260 17172 12288
rect 17328 12260 30788 12288
rect 5810 12180 5816 12232
rect 5868 12220 5874 12232
rect 5997 12223 6055 12229
rect 5997 12220 6009 12223
rect 5868 12192 6009 12220
rect 5868 12180 5874 12192
rect 5997 12189 6009 12192
rect 6043 12220 6055 12223
rect 6270 12220 6276 12232
rect 6043 12192 6276 12220
rect 6043 12189 6055 12192
rect 5997 12183 6055 12189
rect 6270 12180 6276 12192
rect 6328 12180 6334 12232
rect 7190 12180 7196 12232
rect 7248 12220 7254 12232
rect 14292 12229 14320 12260
rect 14277 12223 14335 12229
rect 7248 12192 11652 12220
rect 7248 12180 7254 12192
rect 4249 12155 4307 12161
rect 4249 12121 4261 12155
rect 4295 12121 4307 12155
rect 9122 12152 9128 12164
rect 4249 12115 4307 12121
rect 6104 12124 9128 12152
rect 4264 12084 4292 12115
rect 6104 12084 6132 12124
rect 9122 12112 9128 12124
rect 9180 12152 9186 12164
rect 11238 12152 11244 12164
rect 9180 12124 11244 12152
rect 9180 12112 9186 12124
rect 11238 12112 11244 12124
rect 11296 12112 11302 12164
rect 4264 12056 6132 12084
rect 6178 12044 6184 12096
rect 6236 12084 6242 12096
rect 11514 12084 11520 12096
rect 6236 12056 11520 12084
rect 6236 12044 6242 12056
rect 11514 12044 11520 12056
rect 11572 12044 11578 12096
rect 11624 12084 11652 12192
rect 14277 12189 14289 12223
rect 14323 12189 14335 12223
rect 14277 12183 14335 12189
rect 14366 12180 14372 12232
rect 14424 12220 14430 12232
rect 17328 12220 17356 12260
rect 14424 12192 17356 12220
rect 14424 12180 14430 12192
rect 21818 12180 21824 12232
rect 21876 12220 21882 12232
rect 21913 12223 21971 12229
rect 21913 12220 21925 12223
rect 21876 12192 21925 12220
rect 21876 12180 21882 12192
rect 21913 12189 21925 12192
rect 21959 12189 21971 12223
rect 22557 12223 22615 12229
rect 22557 12220 22569 12223
rect 21913 12183 21971 12189
rect 22066 12192 22569 12220
rect 11882 12112 11888 12164
rect 11940 12152 11946 12164
rect 11940 12124 11985 12152
rect 11940 12112 11946 12124
rect 14550 12112 14556 12164
rect 14608 12152 14614 12164
rect 21450 12152 21456 12164
rect 14608 12124 21456 12152
rect 14608 12112 14614 12124
rect 21450 12112 21456 12124
rect 21508 12112 21514 12164
rect 21542 12112 21548 12164
rect 21600 12152 21606 12164
rect 22066 12152 22094 12192
rect 22557 12189 22569 12192
rect 22603 12189 22615 12223
rect 24854 12220 24860 12232
rect 24815 12192 24860 12220
rect 22557 12183 22615 12189
rect 24854 12180 24860 12192
rect 24912 12180 24918 12232
rect 25498 12180 25504 12232
rect 25556 12220 25562 12232
rect 25961 12223 26019 12229
rect 25961 12220 25973 12223
rect 25556 12192 25973 12220
rect 25556 12180 25562 12192
rect 25961 12189 25973 12192
rect 26007 12189 26019 12223
rect 25961 12183 26019 12189
rect 26145 12223 26203 12229
rect 26145 12189 26157 12223
rect 26191 12220 26203 12223
rect 26694 12220 26700 12232
rect 26191 12192 26700 12220
rect 26191 12189 26203 12192
rect 26145 12183 26203 12189
rect 26694 12180 26700 12192
rect 26752 12180 26758 12232
rect 28828 12229 28856 12260
rect 28813 12223 28871 12229
rect 28813 12189 28825 12223
rect 28859 12189 28871 12223
rect 28813 12183 28871 12189
rect 30285 12223 30343 12229
rect 30285 12189 30297 12223
rect 30331 12189 30343 12223
rect 30760 12220 30788 12260
rect 30834 12248 30840 12300
rect 30892 12288 30898 12300
rect 30929 12291 30987 12297
rect 30929 12288 30941 12291
rect 30892 12260 30941 12288
rect 30892 12248 30898 12260
rect 30929 12257 30941 12260
rect 30975 12257 30987 12291
rect 33226 12288 33232 12300
rect 30929 12251 30987 12257
rect 31726 12260 33232 12288
rect 31726 12220 31754 12260
rect 33226 12248 33232 12260
rect 33284 12248 33290 12300
rect 31846 12220 31852 12232
rect 30760 12192 31754 12220
rect 31807 12192 31852 12220
rect 30285 12183 30343 12189
rect 21600 12124 22094 12152
rect 21600 12112 21606 12124
rect 22738 12112 22744 12164
rect 22796 12152 22802 12164
rect 22833 12155 22891 12161
rect 22833 12152 22845 12155
rect 22796 12124 22845 12152
rect 22796 12112 22802 12124
rect 22833 12121 22845 12124
rect 22879 12121 22891 12155
rect 27706 12152 27712 12164
rect 27667 12124 27712 12152
rect 22833 12115 22891 12121
rect 27706 12112 27712 12124
rect 27764 12112 27770 12164
rect 27801 12155 27859 12161
rect 27801 12121 27813 12155
rect 27847 12152 27859 12155
rect 28074 12152 28080 12164
rect 27847 12124 28080 12152
rect 27847 12121 27859 12124
rect 27801 12115 27859 12121
rect 28074 12112 28080 12124
rect 28132 12112 28138 12164
rect 28718 12112 28724 12164
rect 28776 12152 28782 12164
rect 30300 12152 30328 12183
rect 31846 12180 31852 12192
rect 31904 12180 31910 12232
rect 32674 12180 32680 12232
rect 32732 12220 32738 12232
rect 33321 12223 33379 12229
rect 33321 12220 33333 12223
rect 32732 12192 33333 12220
rect 32732 12180 32738 12192
rect 33321 12189 33333 12192
rect 33367 12189 33379 12223
rect 33321 12183 33379 12189
rect 33413 12223 33471 12229
rect 33413 12189 33425 12223
rect 33459 12220 33471 12223
rect 35989 12223 36047 12229
rect 35989 12220 36001 12223
rect 33459 12192 36001 12220
rect 33459 12189 33471 12192
rect 33413 12183 33471 12189
rect 35989 12189 36001 12192
rect 36035 12189 36047 12223
rect 35989 12183 36047 12189
rect 28776 12124 30328 12152
rect 28776 12112 28782 12124
rect 17218 12084 17224 12096
rect 11624 12056 17224 12084
rect 17218 12044 17224 12056
rect 17276 12044 17282 12096
rect 20898 12044 20904 12096
rect 20956 12084 20962 12096
rect 21082 12084 21088 12096
rect 20956 12056 21088 12084
rect 20956 12044 20962 12056
rect 21082 12044 21088 12056
rect 21140 12044 21146 12096
rect 21910 12044 21916 12096
rect 21968 12084 21974 12096
rect 22005 12087 22063 12093
rect 22005 12084 22017 12087
rect 21968 12056 22017 12084
rect 21968 12044 21974 12056
rect 22005 12053 22017 12056
rect 22051 12053 22063 12087
rect 22005 12047 22063 12053
rect 28905 12087 28963 12093
rect 28905 12053 28917 12087
rect 28951 12084 28963 12087
rect 29178 12084 29184 12096
rect 28951 12056 29184 12084
rect 28951 12053 28963 12056
rect 28905 12047 28963 12053
rect 29178 12044 29184 12056
rect 29236 12044 29242 12096
rect 32309 12087 32367 12093
rect 32309 12053 32321 12087
rect 32355 12084 32367 12087
rect 32398 12084 32404 12096
rect 32355 12056 32404 12084
rect 32355 12053 32367 12056
rect 32309 12047 32367 12053
rect 32398 12044 32404 12056
rect 32456 12044 32462 12096
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 5997 11883 6055 11889
rect 5997 11849 6009 11883
rect 6043 11880 6055 11883
rect 6178 11880 6184 11892
rect 6043 11852 6184 11880
rect 6043 11849 6055 11852
rect 5997 11843 6055 11849
rect 6178 11840 6184 11852
rect 6236 11840 6242 11892
rect 8294 11840 8300 11892
rect 8352 11880 8358 11892
rect 9306 11880 9312 11892
rect 8352 11852 9312 11880
rect 8352 11840 8358 11852
rect 9306 11840 9312 11852
rect 9364 11840 9370 11892
rect 12618 11880 12624 11892
rect 11716 11852 12624 11880
rect 7926 11812 7932 11824
rect 5750 11784 7932 11812
rect 7926 11772 7932 11784
rect 7984 11772 7990 11824
rect 10502 11812 10508 11824
rect 8878 11784 10508 11812
rect 10502 11772 10508 11784
rect 10560 11772 10566 11824
rect 11716 11753 11744 11852
rect 12618 11840 12624 11852
rect 12676 11880 12682 11892
rect 13722 11880 13728 11892
rect 12676 11852 13728 11880
rect 12676 11840 12682 11852
rect 13722 11840 13728 11852
rect 13780 11840 13786 11892
rect 16209 11883 16267 11889
rect 16209 11849 16221 11883
rect 16255 11880 16267 11883
rect 18138 11880 18144 11892
rect 16255 11852 18144 11880
rect 16255 11849 16267 11852
rect 16209 11843 16267 11849
rect 18138 11840 18144 11852
rect 18196 11840 18202 11892
rect 20438 11880 20444 11892
rect 18248 11852 20444 11880
rect 11882 11772 11888 11824
rect 11940 11812 11946 11824
rect 11940 11784 12466 11812
rect 11940 11772 11946 11784
rect 11701 11747 11759 11753
rect 11701 11713 11713 11747
rect 11747 11713 11759 11747
rect 13740 11744 13768 11840
rect 14734 11812 14740 11824
rect 14695 11784 14740 11812
rect 14734 11772 14740 11784
rect 14792 11772 14798 11824
rect 17770 11812 17776 11824
rect 15962 11784 17776 11812
rect 17770 11772 17776 11784
rect 17828 11772 17834 11824
rect 14461 11747 14519 11753
rect 14461 11744 14473 11747
rect 13740 11716 14473 11744
rect 11701 11707 11759 11713
rect 14461 11713 14473 11716
rect 14507 11713 14519 11747
rect 14461 11707 14519 11713
rect 17034 11704 17040 11756
rect 17092 11744 17098 11756
rect 18248 11744 18276 11852
rect 20438 11840 20444 11852
rect 20496 11840 20502 11892
rect 20990 11840 20996 11892
rect 21048 11880 21054 11892
rect 21361 11883 21419 11889
rect 21361 11880 21373 11883
rect 21048 11852 21373 11880
rect 21048 11840 21054 11852
rect 21361 11849 21373 11852
rect 21407 11849 21419 11883
rect 21361 11843 21419 11849
rect 21450 11840 21456 11892
rect 21508 11880 21514 11892
rect 28718 11880 28724 11892
rect 21508 11852 28724 11880
rect 21508 11840 21514 11852
rect 28718 11840 28724 11852
rect 28776 11840 28782 11892
rect 22002 11812 22008 11824
rect 19734 11784 22008 11812
rect 22002 11772 22008 11784
rect 22060 11772 22066 11824
rect 29178 11812 29184 11824
rect 29139 11784 29184 11812
rect 29178 11772 29184 11784
rect 29236 11772 29242 11824
rect 29733 11815 29791 11821
rect 29733 11781 29745 11815
rect 29779 11812 29791 11815
rect 32214 11812 32220 11824
rect 29779 11784 32220 11812
rect 29779 11781 29791 11784
rect 29733 11775 29791 11781
rect 32214 11772 32220 11784
rect 32272 11772 32278 11824
rect 32398 11812 32404 11824
rect 32359 11784 32404 11812
rect 32398 11772 32404 11784
rect 32456 11772 32462 11824
rect 32490 11772 32496 11824
rect 32548 11812 32554 11824
rect 32548 11784 32593 11812
rect 32548 11772 32554 11784
rect 17092 11716 18276 11744
rect 17092 11704 17098 11716
rect 20346 11704 20352 11756
rect 20404 11744 20410 11756
rect 20714 11744 20720 11756
rect 20404 11716 20720 11744
rect 20404 11704 20410 11716
rect 20714 11704 20720 11716
rect 20772 11704 20778 11756
rect 20806 11704 20812 11756
rect 20864 11744 20870 11756
rect 21269 11747 21327 11753
rect 21269 11744 21281 11747
rect 20864 11716 21281 11744
rect 20864 11704 20870 11716
rect 21269 11713 21281 11716
rect 21315 11713 21327 11747
rect 21269 11707 21327 11713
rect 3970 11636 3976 11688
rect 4028 11676 4034 11688
rect 4249 11679 4307 11685
rect 4249 11676 4261 11679
rect 4028 11648 4261 11676
rect 4028 11636 4034 11648
rect 4249 11645 4261 11648
rect 4295 11645 4307 11679
rect 4249 11639 4307 11645
rect 4525 11679 4583 11685
rect 4525 11645 4537 11679
rect 4571 11676 4583 11679
rect 5166 11676 5172 11688
rect 4571 11648 5172 11676
rect 4571 11645 4583 11648
rect 4525 11639 4583 11645
rect 5166 11636 5172 11648
rect 5224 11636 5230 11688
rect 7377 11679 7435 11685
rect 7377 11645 7389 11679
rect 7423 11645 7435 11679
rect 7377 11639 7435 11645
rect 7653 11679 7711 11685
rect 7653 11645 7665 11679
rect 7699 11676 7711 11679
rect 8294 11676 8300 11688
rect 7699 11648 8300 11676
rect 7699 11645 7711 11648
rect 7653 11639 7711 11645
rect 7392 11540 7420 11639
rect 8294 11636 8300 11648
rect 8352 11636 8358 11688
rect 9122 11676 9128 11688
rect 9083 11648 9128 11676
rect 9122 11636 9128 11648
rect 9180 11636 9186 11688
rect 9214 11636 9220 11688
rect 9272 11676 9278 11688
rect 11977 11679 12035 11685
rect 11977 11676 11989 11679
rect 9272 11648 11989 11676
rect 9272 11636 9278 11648
rect 11977 11645 11989 11648
rect 12023 11645 12035 11679
rect 11977 11639 12035 11645
rect 17126 11636 17132 11688
rect 17184 11676 17190 11688
rect 17310 11676 17316 11688
rect 17184 11648 17316 11676
rect 17184 11636 17190 11648
rect 17310 11636 17316 11648
rect 17368 11676 17374 11688
rect 18233 11679 18291 11685
rect 18233 11676 18245 11679
rect 17368 11648 18245 11676
rect 17368 11636 17374 11648
rect 18233 11645 18245 11648
rect 18279 11645 18291 11679
rect 18509 11679 18567 11685
rect 18509 11676 18521 11679
rect 18233 11639 18291 11645
rect 18340 11648 18521 11676
rect 8754 11568 8760 11620
rect 8812 11608 8818 11620
rect 11146 11608 11152 11620
rect 8812 11580 11152 11608
rect 8812 11568 8818 11580
rect 11146 11568 11152 11580
rect 11204 11568 11210 11620
rect 18340 11608 18368 11648
rect 18509 11645 18521 11648
rect 18555 11676 18567 11679
rect 20257 11679 20315 11685
rect 18555 11648 19564 11676
rect 18555 11645 18567 11648
rect 18509 11639 18567 11645
rect 16960 11580 18368 11608
rect 19536 11608 19564 11648
rect 20257 11645 20269 11679
rect 20303 11676 20315 11679
rect 21174 11676 21180 11688
rect 20303 11648 21180 11676
rect 20303 11645 20315 11648
rect 20257 11639 20315 11645
rect 21174 11636 21180 11648
rect 21232 11636 21238 11688
rect 21284 11676 21312 11707
rect 21542 11704 21548 11756
rect 21600 11744 21606 11756
rect 22373 11747 22431 11753
rect 22373 11744 22385 11747
rect 21600 11716 22385 11744
rect 21600 11704 21606 11716
rect 22373 11713 22385 11716
rect 22419 11713 22431 11747
rect 25314 11744 25320 11756
rect 25275 11716 25320 11744
rect 22373 11707 22431 11713
rect 25314 11704 25320 11716
rect 25372 11704 25378 11756
rect 21726 11676 21732 11688
rect 21284 11648 21732 11676
rect 21726 11636 21732 11648
rect 21784 11676 21790 11688
rect 22557 11679 22615 11685
rect 22557 11676 22569 11679
rect 21784 11648 22569 11676
rect 21784 11636 21790 11648
rect 22557 11645 22569 11648
rect 22603 11645 22615 11679
rect 22557 11639 22615 11645
rect 29089 11679 29147 11685
rect 29089 11645 29101 11679
rect 29135 11676 29147 11679
rect 29270 11676 29276 11688
rect 29135 11648 29276 11676
rect 29135 11645 29147 11648
rect 29089 11639 29147 11645
rect 29270 11636 29276 11648
rect 29328 11636 29334 11688
rect 32674 11676 32680 11688
rect 32635 11648 32680 11676
rect 32674 11636 32680 11648
rect 32732 11636 32738 11688
rect 22922 11608 22928 11620
rect 19536 11580 22928 11608
rect 8662 11540 8668 11552
rect 7392 11512 8668 11540
rect 8662 11500 8668 11512
rect 8720 11540 8726 11552
rect 9122 11540 9128 11552
rect 8720 11512 9128 11540
rect 8720 11500 8726 11512
rect 9122 11500 9128 11512
rect 9180 11500 9186 11552
rect 9582 11500 9588 11552
rect 9640 11540 9646 11552
rect 13449 11543 13507 11549
rect 13449 11540 13461 11543
rect 9640 11512 13461 11540
rect 9640 11500 9646 11512
rect 13449 11509 13461 11512
rect 13495 11509 13507 11543
rect 13449 11503 13507 11509
rect 13722 11500 13728 11552
rect 13780 11540 13786 11552
rect 16960 11540 16988 11580
rect 22922 11568 22928 11580
rect 22980 11568 22986 11620
rect 13780 11512 16988 11540
rect 13780 11500 13786 11512
rect 17034 11500 17040 11552
rect 17092 11540 17098 11552
rect 23474 11540 23480 11552
rect 17092 11512 23480 11540
rect 17092 11500 17098 11512
rect 23474 11500 23480 11512
rect 23532 11500 23538 11552
rect 25133 11543 25191 11549
rect 25133 11509 25145 11543
rect 25179 11540 25191 11543
rect 29086 11540 29092 11552
rect 25179 11512 29092 11540
rect 25179 11509 25191 11512
rect 25133 11503 25191 11509
rect 29086 11500 29092 11512
rect 29144 11500 29150 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 5902 11296 5908 11348
rect 5960 11336 5966 11348
rect 9842 11339 9900 11345
rect 9842 11336 9854 11339
rect 5960 11308 9854 11336
rect 5960 11296 5966 11308
rect 9842 11305 9854 11308
rect 9888 11305 9900 11339
rect 9842 11299 9900 11305
rect 11333 11339 11391 11345
rect 11333 11305 11345 11339
rect 11379 11336 11391 11339
rect 11422 11336 11428 11348
rect 11379 11308 11428 11336
rect 11379 11305 11391 11308
rect 11333 11299 11391 11305
rect 11422 11296 11428 11308
rect 11480 11296 11486 11348
rect 20714 11336 20720 11348
rect 12406 11308 20720 11336
rect 1581 11271 1639 11277
rect 1581 11237 1593 11271
rect 1627 11268 1639 11271
rect 1946 11268 1952 11280
rect 1627 11240 1952 11268
rect 1627 11237 1639 11240
rect 1581 11231 1639 11237
rect 1946 11228 1952 11240
rect 2004 11228 2010 11280
rect 6178 11268 6184 11280
rect 5368 11240 6184 11268
rect 4341 11203 4399 11209
rect 4341 11169 4353 11203
rect 4387 11200 4399 11203
rect 5368 11200 5396 11240
rect 6178 11228 6184 11240
rect 6236 11228 6242 11280
rect 7650 11228 7656 11280
rect 7708 11268 7714 11280
rect 9582 11268 9588 11280
rect 7708 11240 9588 11268
rect 7708 11228 7714 11240
rect 9582 11228 9588 11240
rect 9640 11228 9646 11280
rect 12406 11268 12434 11308
rect 20714 11296 20720 11308
rect 20772 11296 20778 11348
rect 25225 11339 25283 11345
rect 25225 11305 25237 11339
rect 25271 11336 25283 11339
rect 25406 11336 25412 11348
rect 25271 11308 25412 11336
rect 25271 11305 25283 11308
rect 25225 11299 25283 11305
rect 25406 11296 25412 11308
rect 25464 11296 25470 11348
rect 26694 11336 26700 11348
rect 26655 11308 26700 11336
rect 26694 11296 26700 11308
rect 26752 11296 26758 11348
rect 28074 11336 28080 11348
rect 28035 11308 28080 11336
rect 28074 11296 28080 11308
rect 28132 11296 28138 11348
rect 28905 11339 28963 11345
rect 28905 11305 28917 11339
rect 28951 11336 28963 11339
rect 32490 11336 32496 11348
rect 28951 11308 32496 11336
rect 28951 11305 28963 11308
rect 28905 11299 28963 11305
rect 32490 11296 32496 11308
rect 32548 11296 32554 11348
rect 38102 11336 38108 11348
rect 38063 11308 38108 11336
rect 38102 11296 38108 11308
rect 38160 11296 38166 11348
rect 10888 11240 12434 11268
rect 23109 11271 23167 11277
rect 10888 11200 10916 11240
rect 23109 11237 23121 11271
rect 23155 11237 23167 11271
rect 23109 11231 23167 11237
rect 4387 11172 5396 11200
rect 5460 11172 10916 11200
rect 4387 11169 4399 11172
rect 4341 11163 4399 11169
rect 1762 11132 1768 11144
rect 1723 11104 1768 11132
rect 1762 11092 1768 11104
rect 1820 11092 1826 11144
rect 3970 11092 3976 11144
rect 4028 11132 4034 11144
rect 4065 11135 4123 11141
rect 4065 11132 4077 11135
rect 4028 11104 4077 11132
rect 4028 11092 4034 11104
rect 4065 11101 4077 11104
rect 4111 11101 4123 11135
rect 5460 11118 5488 11172
rect 11054 11160 11060 11212
rect 11112 11160 11118 11212
rect 11146 11160 11152 11212
rect 11204 11200 11210 11212
rect 17034 11200 17040 11212
rect 11204 11172 17040 11200
rect 11204 11160 11210 11172
rect 17034 11160 17040 11172
rect 17092 11160 17098 11212
rect 17405 11203 17463 11209
rect 17405 11169 17417 11203
rect 17451 11200 17463 11203
rect 17770 11200 17776 11212
rect 17451 11172 17776 11200
rect 17451 11169 17463 11172
rect 17405 11163 17463 11169
rect 17770 11160 17776 11172
rect 17828 11200 17834 11212
rect 18877 11203 18935 11209
rect 17828 11172 18828 11200
rect 17828 11160 17834 11172
rect 4065 11095 4123 11101
rect 5626 11092 5632 11144
rect 5684 11132 5690 11144
rect 6089 11135 6147 11141
rect 6089 11132 6101 11135
rect 5684 11104 6101 11132
rect 5684 11092 5690 11104
rect 6089 11101 6101 11104
rect 6135 11101 6147 11135
rect 6089 11095 6147 11101
rect 6178 11092 6184 11144
rect 6236 11132 6242 11144
rect 6457 11135 6515 11141
rect 6457 11132 6469 11135
rect 6236 11104 6469 11132
rect 6236 11092 6242 11104
rect 6457 11101 6469 11104
rect 6503 11132 6515 11135
rect 8754 11132 8760 11144
rect 6503 11104 8760 11132
rect 6503 11101 6515 11104
rect 6457 11095 6515 11101
rect 8754 11092 8760 11104
rect 8812 11092 8818 11144
rect 9122 11092 9128 11144
rect 9180 11132 9186 11144
rect 9585 11135 9643 11141
rect 9585 11132 9597 11135
rect 9180 11104 9597 11132
rect 9180 11092 9186 11104
rect 9585 11101 9597 11104
rect 9631 11101 9643 11135
rect 11072 11132 11100 11160
rect 11072 11104 16528 11132
rect 9585 11095 9643 11101
rect 9306 11024 9312 11076
rect 9364 11064 9370 11076
rect 16500 11064 16528 11104
rect 16574 11092 16580 11144
rect 16632 11132 16638 11144
rect 17126 11132 17132 11144
rect 16632 11104 17132 11132
rect 16632 11092 16638 11104
rect 17126 11092 17132 11104
rect 17184 11092 17190 11144
rect 18800 11132 18828 11172
rect 18877 11169 18889 11203
rect 18923 11200 18935 11203
rect 18966 11200 18972 11212
rect 18923 11172 18972 11200
rect 18923 11169 18935 11172
rect 18877 11163 18935 11169
rect 18966 11160 18972 11172
rect 19024 11160 19030 11212
rect 19978 11160 19984 11212
rect 20036 11200 20042 11212
rect 23124 11200 23152 11231
rect 31846 11200 31852 11212
rect 20036 11172 22094 11200
rect 23124 11172 23980 11200
rect 20036 11160 20042 11172
rect 21174 11132 21180 11144
rect 18800 11104 21180 11132
rect 21174 11092 21180 11104
rect 21232 11092 21238 11144
rect 21542 11132 21548 11144
rect 21503 11104 21548 11132
rect 21542 11092 21548 11104
rect 21600 11092 21606 11144
rect 17310 11064 17316 11076
rect 9364 11036 9812 11064
rect 9364 11024 9370 11036
rect 6730 10956 6736 11008
rect 6788 10996 6794 11008
rect 6825 10999 6883 11005
rect 6825 10996 6837 10999
rect 6788 10968 6837 10996
rect 6788 10956 6794 10968
rect 6825 10965 6837 10968
rect 6871 10965 6883 10999
rect 9784 10996 9812 11036
rect 9968 11036 10350 11064
rect 16500 11036 17316 11064
rect 9968 10996 9996 11036
rect 17310 11024 17316 11036
rect 17368 11024 17374 11076
rect 20162 11064 20168 11076
rect 18630 11036 20168 11064
rect 20162 11024 20168 11036
rect 20220 11024 20226 11076
rect 21634 11024 21640 11076
rect 21692 11064 21698 11076
rect 21821 11067 21879 11073
rect 21821 11064 21833 11067
rect 21692 11036 21833 11064
rect 21692 11024 21698 11036
rect 21821 11033 21833 11036
rect 21867 11033 21879 11067
rect 22066 11064 22094 11172
rect 23290 11132 23296 11144
rect 23251 11104 23296 11132
rect 23290 11092 23296 11104
rect 23348 11092 23354 11144
rect 23952 11141 23980 11172
rect 28000 11172 31852 11200
rect 23937 11135 23995 11141
rect 23937 11101 23949 11135
rect 23983 11101 23995 11135
rect 23937 11095 23995 11101
rect 24581 11135 24639 11141
rect 24581 11101 24593 11135
rect 24627 11132 24639 11135
rect 24670 11132 24676 11144
rect 24627 11104 24676 11132
rect 24627 11101 24639 11104
rect 24581 11095 24639 11101
rect 24670 11092 24676 11104
rect 24728 11092 24734 11144
rect 24765 11135 24823 11141
rect 24765 11101 24777 11135
rect 24811 11132 24823 11135
rect 25038 11132 25044 11144
rect 24811 11104 25044 11132
rect 24811 11101 24823 11104
rect 24765 11095 24823 11101
rect 25038 11092 25044 11104
rect 25096 11092 25102 11144
rect 26510 11092 26516 11144
rect 26568 11132 26574 11144
rect 28000 11141 28028 11172
rect 31846 11160 31852 11172
rect 31904 11160 31910 11212
rect 26605 11135 26663 11141
rect 26605 11132 26617 11135
rect 26568 11104 26617 11132
rect 26568 11092 26574 11104
rect 26605 11101 26617 11104
rect 26651 11101 26663 11135
rect 26605 11095 26663 11101
rect 27985 11135 28043 11141
rect 27985 11101 27997 11135
rect 28031 11101 28043 11135
rect 29086 11132 29092 11144
rect 29047 11104 29092 11132
rect 27985 11095 28043 11101
rect 28000 11064 28028 11095
rect 29086 11092 29092 11104
rect 29144 11092 29150 11144
rect 31294 11092 31300 11144
rect 31352 11132 31358 11144
rect 31389 11135 31447 11141
rect 31389 11132 31401 11135
rect 31352 11104 31401 11132
rect 31352 11092 31358 11104
rect 31389 11101 31401 11104
rect 31435 11101 31447 11135
rect 38286 11132 38292 11144
rect 38247 11104 38292 11132
rect 31389 11095 31447 11101
rect 38286 11092 38292 11104
rect 38344 11092 38350 11144
rect 22066 11036 28028 11064
rect 31481 11067 31539 11073
rect 21821 11027 21879 11033
rect 31481 11033 31493 11067
rect 31527 11064 31539 11067
rect 33042 11064 33048 11076
rect 31527 11036 33048 11064
rect 31527 11033 31539 11036
rect 31481 11027 31539 11033
rect 33042 11024 33048 11036
rect 33100 11024 33106 11076
rect 9784 10968 9996 10996
rect 6825 10959 6883 10965
rect 12250 10956 12256 11008
rect 12308 10996 12314 11008
rect 14918 10996 14924 11008
rect 12308 10968 14924 10996
rect 12308 10956 12314 10968
rect 14918 10956 14924 10968
rect 14976 10956 14982 11008
rect 15102 10956 15108 11008
rect 15160 10996 15166 11008
rect 21450 10996 21456 11008
rect 15160 10968 21456 10996
rect 15160 10956 15166 10968
rect 21450 10956 21456 10968
rect 21508 10956 21514 11008
rect 23753 10999 23811 11005
rect 23753 10965 23765 10999
rect 23799 10996 23811 10999
rect 24762 10996 24768 11008
rect 23799 10968 24768 10996
rect 23799 10965 23811 10968
rect 23753 10959 23811 10965
rect 24762 10956 24768 10968
rect 24820 10956 24826 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 6546 10752 6552 10804
rect 6604 10792 6610 10804
rect 6604 10764 6868 10792
rect 6604 10752 6610 10764
rect 5442 10724 5448 10736
rect 5403 10696 5448 10724
rect 5442 10684 5448 10696
rect 5500 10684 5506 10736
rect 5997 10727 6055 10733
rect 5997 10693 6009 10727
rect 6043 10724 6055 10727
rect 6086 10724 6092 10736
rect 6043 10696 6092 10724
rect 6043 10693 6055 10696
rect 5997 10687 6055 10693
rect 6086 10684 6092 10696
rect 6144 10684 6150 10736
rect 6730 10724 6736 10736
rect 6691 10696 6736 10724
rect 6730 10684 6736 10696
rect 6788 10684 6794 10736
rect 6840 10733 6868 10764
rect 7926 10752 7932 10804
rect 7984 10792 7990 10804
rect 10597 10795 10655 10801
rect 10597 10792 10609 10795
rect 7984 10764 10609 10792
rect 7984 10752 7990 10764
rect 10597 10761 10609 10764
rect 10643 10761 10655 10795
rect 10597 10755 10655 10761
rect 15010 10752 15016 10804
rect 15068 10792 15074 10804
rect 18601 10795 18659 10801
rect 18601 10792 18613 10795
rect 15068 10764 18613 10792
rect 15068 10752 15074 10764
rect 18601 10761 18613 10764
rect 18647 10761 18659 10795
rect 18601 10755 18659 10761
rect 20714 10752 20720 10804
rect 20772 10792 20778 10804
rect 22462 10792 22468 10804
rect 20772 10764 22468 10792
rect 20772 10752 20778 10764
rect 22462 10752 22468 10764
rect 22520 10752 22526 10804
rect 25038 10792 25044 10804
rect 24999 10764 25044 10792
rect 25038 10752 25044 10764
rect 25096 10752 25102 10804
rect 6825 10727 6883 10733
rect 6825 10693 6837 10727
rect 6871 10693 6883 10727
rect 6825 10687 6883 10693
rect 12897 10727 12955 10733
rect 12897 10693 12909 10727
rect 12943 10724 12955 10727
rect 13170 10724 13176 10736
rect 12943 10696 13176 10724
rect 12943 10693 12955 10696
rect 12897 10687 12955 10693
rect 13170 10684 13176 10696
rect 13228 10684 13234 10736
rect 17402 10724 17408 10736
rect 14936 10696 17408 10724
rect 1578 10616 1584 10668
rect 1636 10656 1642 10668
rect 1857 10659 1915 10665
rect 1857 10656 1869 10659
rect 1636 10628 1869 10656
rect 1636 10616 1642 10628
rect 1857 10625 1869 10628
rect 1903 10625 1915 10659
rect 1857 10619 1915 10625
rect 10505 10659 10563 10665
rect 10505 10625 10517 10659
rect 10551 10656 10563 10659
rect 11330 10656 11336 10668
rect 10551 10628 11336 10656
rect 10551 10625 10563 10628
rect 10505 10619 10563 10625
rect 11330 10616 11336 10628
rect 11388 10616 11394 10668
rect 12618 10656 12624 10668
rect 12579 10628 12624 10656
rect 12618 10616 12624 10628
rect 12676 10616 12682 10668
rect 13998 10616 14004 10668
rect 14056 10616 14062 10668
rect 1949 10591 2007 10597
rect 1949 10557 1961 10591
rect 1995 10588 2007 10591
rect 5353 10591 5411 10597
rect 5353 10588 5365 10591
rect 1995 10560 5365 10588
rect 1995 10557 2007 10560
rect 1949 10551 2007 10557
rect 5353 10557 5365 10560
rect 5399 10557 5411 10591
rect 7006 10588 7012 10600
rect 6967 10560 7012 10588
rect 5353 10551 5411 10557
rect 7006 10548 7012 10560
rect 7064 10548 7070 10600
rect 8386 10548 8392 10600
rect 8444 10588 8450 10600
rect 14936 10588 14964 10696
rect 17402 10684 17408 10696
rect 17460 10684 17466 10736
rect 21910 10724 21916 10736
rect 18354 10696 21916 10724
rect 21910 10684 21916 10696
rect 21968 10684 21974 10736
rect 22281 10727 22339 10733
rect 22281 10693 22293 10727
rect 22327 10724 22339 10727
rect 22370 10724 22376 10736
rect 22327 10696 22376 10724
rect 22327 10693 22339 10696
rect 22281 10687 22339 10693
rect 22370 10684 22376 10696
rect 22428 10684 22434 10736
rect 23658 10724 23664 10736
rect 23619 10696 23664 10724
rect 23658 10684 23664 10696
rect 23716 10684 23722 10736
rect 20806 10656 20812 10668
rect 20767 10628 20812 10656
rect 20806 10616 20812 10628
rect 20864 10656 20870 10668
rect 21542 10656 21548 10668
rect 20864 10628 21548 10656
rect 20864 10616 20870 10628
rect 21542 10616 21548 10628
rect 21600 10656 21606 10668
rect 22005 10659 22063 10665
rect 22005 10656 22017 10659
rect 21600 10628 22017 10656
rect 21600 10616 21606 10628
rect 22005 10625 22017 10628
rect 22051 10625 22063 10659
rect 25222 10656 25228 10668
rect 25183 10628 25228 10656
rect 22005 10619 22063 10625
rect 25222 10616 25228 10628
rect 25280 10616 25286 10668
rect 28718 10656 28724 10668
rect 28679 10628 28724 10656
rect 28718 10616 28724 10628
rect 28776 10616 28782 10668
rect 29362 10656 29368 10668
rect 29323 10628 29368 10656
rect 29362 10616 29368 10628
rect 29420 10616 29426 10668
rect 29825 10659 29883 10665
rect 29825 10625 29837 10659
rect 29871 10656 29883 10659
rect 30098 10656 30104 10668
rect 29871 10628 30104 10656
rect 29871 10625 29883 10628
rect 29825 10619 29883 10625
rect 30098 10616 30104 10628
rect 30156 10616 30162 10668
rect 33042 10616 33048 10668
rect 33100 10656 33106 10668
rect 33965 10659 34023 10665
rect 33965 10656 33977 10659
rect 33100 10628 33977 10656
rect 33100 10616 33106 10628
rect 33965 10625 33977 10628
rect 34011 10625 34023 10659
rect 33965 10619 34023 10625
rect 8444 10560 14964 10588
rect 8444 10548 8450 10560
rect 16574 10548 16580 10600
rect 16632 10588 16638 10600
rect 16853 10591 16911 10597
rect 16853 10588 16865 10591
rect 16632 10560 16865 10588
rect 16632 10548 16638 10560
rect 16853 10557 16865 10560
rect 16899 10557 16911 10591
rect 16853 10551 16911 10557
rect 17129 10591 17187 10597
rect 17129 10557 17141 10591
rect 17175 10588 17187 10591
rect 19150 10588 19156 10600
rect 17175 10560 19156 10588
rect 17175 10557 17187 10560
rect 17129 10551 17187 10557
rect 19150 10548 19156 10560
rect 19208 10548 19214 10600
rect 20898 10548 20904 10600
rect 20956 10588 20962 10600
rect 20993 10591 21051 10597
rect 20993 10588 21005 10591
rect 20956 10560 21005 10588
rect 20956 10548 20962 10560
rect 20993 10557 21005 10560
rect 21039 10557 21051 10591
rect 20993 10551 21051 10557
rect 22830 10548 22836 10600
rect 22888 10588 22894 10600
rect 23569 10591 23627 10597
rect 23569 10588 23581 10591
rect 22888 10560 23581 10588
rect 22888 10548 22894 10560
rect 23569 10557 23581 10560
rect 23615 10557 23627 10591
rect 23569 10551 23627 10557
rect 23845 10591 23903 10597
rect 23845 10557 23857 10591
rect 23891 10557 23903 10591
rect 23845 10551 23903 10557
rect 6638 10480 6644 10532
rect 6696 10520 6702 10532
rect 9858 10520 9864 10532
rect 6696 10492 9864 10520
rect 6696 10480 6702 10492
rect 9858 10480 9864 10492
rect 9916 10480 9922 10532
rect 13924 10492 14504 10520
rect 13630 10412 13636 10464
rect 13688 10452 13694 10464
rect 13924 10452 13952 10492
rect 14366 10452 14372 10464
rect 13688 10424 13952 10452
rect 14327 10424 14372 10452
rect 13688 10412 13694 10424
rect 14366 10412 14372 10424
rect 14424 10412 14430 10464
rect 14476 10452 14504 10492
rect 21266 10480 21272 10532
rect 21324 10520 21330 10532
rect 23860 10520 23888 10551
rect 29914 10548 29920 10600
rect 29972 10588 29978 10600
rect 30009 10591 30067 10597
rect 30009 10588 30021 10591
rect 29972 10560 30021 10588
rect 29972 10548 29978 10560
rect 30009 10557 30021 10560
rect 30055 10557 30067 10591
rect 30009 10551 30067 10557
rect 21324 10492 23888 10520
rect 28537 10523 28595 10529
rect 21324 10480 21330 10492
rect 28537 10489 28549 10523
rect 28583 10520 28595 10523
rect 30374 10520 30380 10532
rect 28583 10492 30380 10520
rect 28583 10489 28595 10492
rect 28537 10483 28595 10489
rect 30374 10480 30380 10492
rect 30432 10480 30438 10532
rect 21358 10452 21364 10464
rect 14476 10424 21364 10452
rect 21358 10412 21364 10424
rect 21416 10412 21422 10464
rect 21450 10412 21456 10464
rect 21508 10452 21514 10464
rect 23934 10452 23940 10464
rect 21508 10424 23940 10452
rect 21508 10412 21514 10424
rect 23934 10412 23940 10424
rect 23992 10412 23998 10464
rect 24026 10412 24032 10464
rect 24084 10452 24090 10464
rect 27798 10452 27804 10464
rect 24084 10424 27804 10452
rect 24084 10412 24090 10424
rect 27798 10412 27804 10424
rect 27856 10412 27862 10464
rect 29181 10455 29239 10461
rect 29181 10421 29193 10455
rect 29227 10452 29239 10455
rect 30006 10452 30012 10464
rect 29227 10424 30012 10452
rect 29227 10421 29239 10424
rect 29181 10415 29239 10421
rect 30006 10412 30012 10424
rect 30064 10412 30070 10464
rect 30469 10455 30527 10461
rect 30469 10421 30481 10455
rect 30515 10452 30527 10455
rect 30558 10452 30564 10464
rect 30515 10424 30564 10452
rect 30515 10421 30527 10424
rect 30469 10415 30527 10421
rect 30558 10412 30564 10424
rect 30616 10412 30622 10464
rect 33781 10455 33839 10461
rect 33781 10421 33793 10455
rect 33827 10452 33839 10455
rect 34790 10452 34796 10464
rect 33827 10424 34796 10452
rect 33827 10421 33839 10424
rect 33781 10415 33839 10421
rect 34790 10412 34796 10424
rect 34848 10412 34854 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 4614 10208 4620 10260
rect 4672 10248 4678 10260
rect 12158 10248 12164 10260
rect 4672 10220 12164 10248
rect 4672 10208 4678 10220
rect 12158 10208 12164 10220
rect 12216 10208 12222 10260
rect 13998 10208 14004 10260
rect 14056 10248 14062 10260
rect 22741 10251 22799 10257
rect 22741 10248 22753 10251
rect 14056 10220 22753 10248
rect 14056 10208 14062 10220
rect 22741 10217 22753 10220
rect 22787 10217 22799 10251
rect 22741 10211 22799 10217
rect 23477 10251 23535 10257
rect 23477 10217 23489 10251
rect 23523 10248 23535 10251
rect 25222 10248 25228 10260
rect 23523 10220 25228 10248
rect 23523 10217 23535 10220
rect 23477 10211 23535 10217
rect 25222 10208 25228 10220
rect 25280 10208 25286 10260
rect 29825 10251 29883 10257
rect 29825 10217 29837 10251
rect 29871 10248 29883 10251
rect 29914 10248 29920 10260
rect 29871 10220 29920 10248
rect 29871 10217 29883 10220
rect 29825 10211 29883 10217
rect 29914 10208 29920 10220
rect 29972 10208 29978 10260
rect 10870 10140 10876 10192
rect 10928 10180 10934 10192
rect 15194 10180 15200 10192
rect 10928 10152 15200 10180
rect 10928 10140 10934 10152
rect 15194 10140 15200 10152
rect 15252 10140 15258 10192
rect 17310 10140 17316 10192
rect 17368 10180 17374 10192
rect 21453 10183 21511 10189
rect 21453 10180 21465 10183
rect 17368 10152 21465 10180
rect 17368 10140 17374 10152
rect 21453 10149 21465 10152
rect 21499 10149 21511 10183
rect 24026 10180 24032 10192
rect 21453 10143 21511 10149
rect 21560 10152 24032 10180
rect 4249 10115 4307 10121
rect 4249 10081 4261 10115
rect 4295 10112 4307 10115
rect 5258 10112 5264 10124
rect 4295 10084 5264 10112
rect 4295 10081 4307 10084
rect 4249 10075 4307 10081
rect 5258 10072 5264 10084
rect 5316 10072 5322 10124
rect 5368 10084 12434 10112
rect 1762 10044 1768 10056
rect 1723 10016 1768 10044
rect 1762 10004 1768 10016
rect 1820 10004 1826 10056
rect 3970 10044 3976 10056
rect 3931 10016 3976 10044
rect 3970 10004 3976 10016
rect 4028 10004 4034 10056
rect 5368 10030 5396 10084
rect 12406 10044 12434 10084
rect 14366 10072 14372 10124
rect 14424 10112 14430 10124
rect 14550 10112 14556 10124
rect 14424 10084 14556 10112
rect 14424 10072 14430 10084
rect 14550 10072 14556 10084
rect 14608 10112 14614 10124
rect 21560 10112 21588 10152
rect 24026 10140 24032 10152
rect 24084 10140 24090 10192
rect 24210 10140 24216 10192
rect 24268 10180 24274 10192
rect 24946 10180 24952 10192
rect 24268 10152 24952 10180
rect 24268 10140 24274 10152
rect 24946 10140 24952 10152
rect 25004 10140 25010 10192
rect 14608 10084 21588 10112
rect 14608 10072 14614 10084
rect 22094 10072 22100 10124
rect 22152 10112 22158 10124
rect 24673 10115 24731 10121
rect 22152 10084 22197 10112
rect 22152 10072 22158 10084
rect 24673 10081 24685 10115
rect 24719 10112 24731 10115
rect 25038 10112 25044 10124
rect 24719 10084 25044 10112
rect 24719 10081 24731 10084
rect 24673 10075 24731 10081
rect 25038 10072 25044 10084
rect 25096 10072 25102 10124
rect 20441 10047 20499 10053
rect 12406 10016 20392 10044
rect 5902 9936 5908 9988
rect 5960 9976 5966 9988
rect 5997 9979 6055 9985
rect 5997 9976 6009 9979
rect 5960 9948 6009 9976
rect 5960 9936 5966 9948
rect 5997 9945 6009 9948
rect 6043 9945 6055 9979
rect 5997 9939 6055 9945
rect 6086 9936 6092 9988
rect 6144 9976 6150 9988
rect 6549 9979 6607 9985
rect 6549 9976 6561 9979
rect 6144 9948 6561 9976
rect 6144 9936 6150 9948
rect 6549 9945 6561 9948
rect 6595 9945 6607 9979
rect 6549 9939 6607 9945
rect 6641 9979 6699 9985
rect 6641 9945 6653 9979
rect 6687 9945 6699 9979
rect 6641 9939 6699 9945
rect 7193 9979 7251 9985
rect 7193 9945 7205 9979
rect 7239 9976 7251 9979
rect 12526 9976 12532 9988
rect 7239 9948 12532 9976
rect 7239 9945 7251 9948
rect 7193 9939 7251 9945
rect 1581 9911 1639 9917
rect 1581 9877 1593 9911
rect 1627 9908 1639 9911
rect 1854 9908 1860 9920
rect 1627 9880 1860 9908
rect 1627 9877 1639 9880
rect 1581 9871 1639 9877
rect 1854 9868 1860 9880
rect 1912 9868 1918 9920
rect 4890 9868 4896 9920
rect 4948 9908 4954 9920
rect 6656 9908 6684 9939
rect 12526 9936 12532 9948
rect 12584 9976 12590 9988
rect 13630 9976 13636 9988
rect 12584 9948 13636 9976
rect 12584 9936 12590 9948
rect 13630 9936 13636 9948
rect 13688 9936 13694 9988
rect 14918 9936 14924 9988
rect 14976 9976 14982 9988
rect 20070 9976 20076 9988
rect 14976 9948 20076 9976
rect 14976 9936 14982 9948
rect 20070 9936 20076 9948
rect 20128 9936 20134 9988
rect 20364 9976 20392 10016
rect 20441 10013 20453 10047
rect 20487 10044 20499 10047
rect 20714 10044 20720 10056
rect 20487 10016 20720 10044
rect 20487 10013 20499 10016
rect 20441 10007 20499 10013
rect 20714 10004 20720 10016
rect 20772 10004 20778 10056
rect 21361 10047 21419 10053
rect 21361 10013 21373 10047
rect 21407 10044 21419 10047
rect 22005 10047 22063 10053
rect 22005 10044 22017 10047
rect 21407 10016 22017 10044
rect 21407 10013 21419 10016
rect 21361 10007 21419 10013
rect 22005 10013 22017 10016
rect 22051 10013 22063 10047
rect 22005 10007 22063 10013
rect 21542 9976 21548 9988
rect 20364 9948 21548 9976
rect 21542 9936 21548 9948
rect 21600 9936 21606 9988
rect 22020 9976 22048 10007
rect 22370 10004 22376 10056
rect 22428 10044 22434 10056
rect 22649 10047 22707 10053
rect 22649 10044 22661 10047
rect 22428 10016 22661 10044
rect 22428 10004 22434 10016
rect 22649 10013 22661 10016
rect 22695 10013 22707 10047
rect 22649 10007 22707 10013
rect 23661 10047 23719 10053
rect 23661 10013 23673 10047
rect 23707 10044 23719 10047
rect 23934 10044 23940 10056
rect 23707 10016 23940 10044
rect 23707 10013 23719 10016
rect 23661 10007 23719 10013
rect 23934 10004 23940 10016
rect 23992 10004 23998 10056
rect 30006 10044 30012 10056
rect 29967 10016 30012 10044
rect 30006 10004 30012 10016
rect 30064 10004 30070 10056
rect 22738 9976 22744 9988
rect 22020 9948 22744 9976
rect 22738 9936 22744 9948
rect 22796 9936 22802 9988
rect 24762 9936 24768 9988
rect 24820 9976 24826 9988
rect 25685 9979 25743 9985
rect 24820 9948 24865 9976
rect 24820 9936 24826 9948
rect 25685 9945 25697 9979
rect 25731 9945 25743 9979
rect 25685 9939 25743 9945
rect 4948 9880 6684 9908
rect 4948 9868 4954 9880
rect 9306 9868 9312 9920
rect 9364 9908 9370 9920
rect 20533 9911 20591 9917
rect 20533 9908 20545 9911
rect 9364 9880 20545 9908
rect 9364 9868 9370 9880
rect 20533 9877 20545 9880
rect 20579 9877 20591 9911
rect 20533 9871 20591 9877
rect 22094 9868 22100 9920
rect 22152 9908 22158 9920
rect 25130 9908 25136 9920
rect 22152 9880 25136 9908
rect 22152 9868 22158 9880
rect 25130 9868 25136 9880
rect 25188 9908 25194 9920
rect 25700 9908 25728 9939
rect 25188 9880 25728 9908
rect 25188 9868 25194 9880
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 15749 9707 15807 9713
rect 15749 9673 15761 9707
rect 15795 9673 15807 9707
rect 15749 9667 15807 9673
rect 18892 9676 19840 9704
rect 9401 9639 9459 9645
rect 9401 9636 9413 9639
rect 9140 9608 9413 9636
rect 8110 9528 8116 9580
rect 8168 9528 8174 9580
rect 9140 9568 9168 9608
rect 9401 9605 9413 9608
rect 9447 9605 9459 9639
rect 15764 9636 15792 9667
rect 18892 9636 18920 9676
rect 15764 9608 18920 9636
rect 19812 9636 19840 9676
rect 20438 9664 20444 9716
rect 20496 9704 20502 9716
rect 20496 9676 21312 9704
rect 20496 9664 20502 9676
rect 19978 9636 19984 9648
rect 19812 9608 19984 9636
rect 9401 9599 9459 9605
rect 19978 9596 19984 9608
rect 20036 9596 20042 9648
rect 20162 9596 20168 9648
rect 20220 9636 20226 9648
rect 20625 9639 20683 9645
rect 20625 9636 20637 9639
rect 20220 9608 20637 9636
rect 20220 9596 20226 9608
rect 20625 9605 20637 9608
rect 20671 9605 20683 9639
rect 21082 9636 21088 9648
rect 20625 9599 20683 9605
rect 20732 9608 21088 9636
rect 8220 9540 9168 9568
rect 6546 9460 6552 9512
rect 6604 9500 6610 9512
rect 6733 9503 6791 9509
rect 6733 9500 6745 9503
rect 6604 9472 6745 9500
rect 6604 9460 6610 9472
rect 6733 9469 6745 9472
rect 6779 9469 6791 9503
rect 6733 9463 6791 9469
rect 7650 9460 7656 9512
rect 7708 9500 7714 9512
rect 8220 9500 8248 9540
rect 10502 9528 10508 9580
rect 10560 9528 10566 9580
rect 18138 9568 18144 9580
rect 15410 9540 18144 9568
rect 18138 9528 18144 9540
rect 18196 9528 18202 9580
rect 7708 9472 8248 9500
rect 7708 9460 7714 9472
rect 8294 9460 8300 9512
rect 8352 9500 8358 9512
rect 8481 9503 8539 9509
rect 8481 9500 8493 9503
rect 8352 9472 8493 9500
rect 8352 9460 8358 9472
rect 8481 9469 8493 9472
rect 8527 9469 8539 9503
rect 9122 9500 9128 9512
rect 9083 9472 9128 9500
rect 8481 9463 8539 9469
rect 9122 9460 9128 9472
rect 9180 9460 9186 9512
rect 11149 9503 11207 9509
rect 9232 9472 11100 9500
rect 8018 9392 8024 9444
rect 8076 9432 8082 9444
rect 9232 9432 9260 9472
rect 8076 9404 9260 9432
rect 11072 9432 11100 9472
rect 11149 9469 11161 9503
rect 11195 9500 11207 9503
rect 14001 9503 14059 9509
rect 11195 9472 12434 9500
rect 11195 9469 11207 9472
rect 11149 9463 11207 9469
rect 12250 9432 12256 9444
rect 11072 9404 12256 9432
rect 8076 9392 8082 9404
rect 12250 9392 12256 9404
rect 12308 9392 12314 9444
rect 12406 9432 12434 9472
rect 14001 9469 14013 9503
rect 14047 9469 14059 9503
rect 14001 9463 14059 9469
rect 14277 9503 14335 9509
rect 14277 9469 14289 9503
rect 14323 9500 14335 9503
rect 14323 9472 17908 9500
rect 14323 9469 14335 9472
rect 14277 9463 14335 9469
rect 13906 9432 13912 9444
rect 12406 9404 13912 9432
rect 13906 9392 13912 9404
rect 13964 9392 13970 9444
rect 6996 9367 7054 9373
rect 6996 9333 7008 9367
rect 7042 9364 7054 9367
rect 11974 9364 11980 9376
rect 7042 9336 11980 9364
rect 7042 9333 7054 9336
rect 6996 9327 7054 9333
rect 11974 9324 11980 9336
rect 12032 9324 12038 9376
rect 14016 9364 14044 9463
rect 14274 9364 14280 9376
rect 14016 9336 14280 9364
rect 14274 9324 14280 9336
rect 14332 9324 14338 9376
rect 17880 9364 17908 9472
rect 17954 9460 17960 9512
rect 18012 9500 18018 9512
rect 18233 9503 18291 9509
rect 18233 9500 18245 9503
rect 18012 9472 18245 9500
rect 18012 9460 18018 9472
rect 18233 9469 18245 9472
rect 18279 9469 18291 9503
rect 18233 9463 18291 9469
rect 18509 9503 18567 9509
rect 18509 9469 18521 9503
rect 18555 9500 18567 9503
rect 19150 9500 19156 9512
rect 18555 9472 19156 9500
rect 18555 9469 18567 9472
rect 18509 9463 18567 9469
rect 19150 9460 19156 9472
rect 19208 9460 19214 9512
rect 19242 9460 19248 9512
rect 19300 9500 19306 9512
rect 19628 9500 19656 9554
rect 20070 9528 20076 9580
rect 20128 9568 20134 9580
rect 20438 9568 20444 9580
rect 20128 9540 20444 9568
rect 20128 9528 20134 9540
rect 20438 9528 20444 9540
rect 20496 9528 20502 9580
rect 20533 9571 20591 9577
rect 20533 9537 20545 9571
rect 20579 9568 20591 9571
rect 20732 9568 20760 9608
rect 21082 9596 21088 9608
rect 21140 9596 21146 9648
rect 21284 9645 21312 9676
rect 21358 9664 21364 9716
rect 21416 9704 21422 9716
rect 22830 9704 22836 9716
rect 21416 9676 22836 9704
rect 21416 9664 21422 9676
rect 22830 9664 22836 9676
rect 22888 9664 22894 9716
rect 23658 9704 23664 9716
rect 23619 9676 23664 9704
rect 23658 9664 23664 9676
rect 23716 9664 23722 9716
rect 21269 9639 21327 9645
rect 21269 9605 21281 9639
rect 21315 9605 21327 9639
rect 21269 9599 21327 9605
rect 20579 9540 20760 9568
rect 20579 9537 20591 9540
rect 20533 9531 20591 9537
rect 20806 9528 20812 9580
rect 20864 9568 20870 9580
rect 21177 9571 21235 9577
rect 21177 9568 21189 9571
rect 20864 9540 21189 9568
rect 20864 9528 20870 9540
rect 21177 9537 21189 9540
rect 21223 9568 21235 9571
rect 22002 9568 22008 9580
rect 21223 9540 22008 9568
rect 21223 9537 21235 9540
rect 21177 9531 21235 9537
rect 22002 9528 22008 9540
rect 22060 9528 22066 9580
rect 22554 9568 22560 9580
rect 22467 9540 22560 9568
rect 22554 9528 22560 9540
rect 22612 9568 22618 9580
rect 23569 9571 23627 9577
rect 22612 9540 23520 9568
rect 22612 9528 22618 9540
rect 19300 9472 19564 9500
rect 19628 9472 22094 9500
rect 19300 9460 19306 9472
rect 19536 9432 19564 9472
rect 21910 9432 21916 9444
rect 19536 9404 21916 9432
rect 21910 9392 21916 9404
rect 21968 9392 21974 9444
rect 22066 9432 22094 9472
rect 23492 9432 23520 9540
rect 23569 9537 23581 9571
rect 23615 9568 23627 9571
rect 24762 9568 24768 9580
rect 23615 9540 24768 9568
rect 23615 9537 23627 9540
rect 23569 9531 23627 9537
rect 24762 9528 24768 9540
rect 24820 9528 24826 9580
rect 29273 9571 29331 9577
rect 29273 9537 29285 9571
rect 29319 9568 29331 9571
rect 30558 9568 30564 9580
rect 29319 9540 30564 9568
rect 29319 9537 29331 9540
rect 29273 9531 29331 9537
rect 30558 9528 30564 9540
rect 30616 9528 30622 9580
rect 25222 9460 25228 9512
rect 25280 9500 25286 9512
rect 28629 9503 28687 9509
rect 28629 9500 28641 9503
rect 25280 9472 28641 9500
rect 25280 9460 25286 9472
rect 28629 9469 28641 9472
rect 28675 9469 28687 9503
rect 28629 9463 28687 9469
rect 28718 9460 28724 9512
rect 28776 9500 28782 9512
rect 28813 9503 28871 9509
rect 28813 9500 28825 9503
rect 28776 9472 28825 9500
rect 28776 9460 28782 9472
rect 28813 9469 28825 9472
rect 28859 9469 28871 9503
rect 28813 9463 28871 9469
rect 37734 9432 37740 9444
rect 22066 9404 23428 9432
rect 23492 9404 37740 9432
rect 19981 9367 20039 9373
rect 19981 9364 19993 9367
rect 17880 9336 19993 9364
rect 19981 9333 19993 9336
rect 20027 9364 20039 9367
rect 20530 9364 20536 9376
rect 20027 9336 20536 9364
rect 20027 9333 20039 9336
rect 19981 9327 20039 9333
rect 20530 9324 20536 9336
rect 20588 9324 20594 9376
rect 21082 9324 21088 9376
rect 21140 9364 21146 9376
rect 21634 9364 21640 9376
rect 21140 9336 21640 9364
rect 21140 9324 21146 9336
rect 21634 9324 21640 9336
rect 21692 9324 21698 9376
rect 22002 9324 22008 9376
rect 22060 9364 22066 9376
rect 22649 9367 22707 9373
rect 22649 9364 22661 9367
rect 22060 9336 22661 9364
rect 22060 9324 22066 9336
rect 22649 9333 22661 9336
rect 22695 9333 22707 9367
rect 23400 9364 23428 9404
rect 37734 9392 37740 9404
rect 37792 9392 37798 9444
rect 23474 9364 23480 9376
rect 23400 9336 23480 9364
rect 22649 9327 22707 9333
rect 23474 9324 23480 9336
rect 23532 9324 23538 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 7006 9120 7012 9172
rect 7064 9160 7070 9172
rect 8018 9160 8024 9172
rect 7064 9132 8024 9160
rect 7064 9120 7070 9132
rect 8018 9120 8024 9132
rect 8076 9120 8082 9172
rect 8110 9120 8116 9172
rect 8168 9160 8174 9172
rect 21082 9160 21088 9172
rect 8168 9132 21088 9160
rect 8168 9120 8174 9132
rect 21082 9120 21088 9132
rect 21140 9120 21146 9172
rect 21174 9120 21180 9172
rect 21232 9160 21238 9172
rect 28718 9160 28724 9172
rect 21232 9132 25820 9160
rect 28679 9132 28724 9160
rect 21232 9120 21238 9132
rect 8478 9052 8484 9104
rect 8536 9092 8542 9104
rect 14458 9092 14464 9104
rect 8536 9064 14464 9092
rect 8536 9052 8542 9064
rect 14458 9052 14464 9064
rect 14516 9052 14522 9104
rect 18138 9052 18144 9104
rect 18196 9092 18202 9104
rect 23569 9095 23627 9101
rect 23569 9092 23581 9095
rect 18196 9064 23581 9092
rect 18196 9052 18202 9064
rect 23569 9061 23581 9064
rect 23615 9061 23627 9095
rect 25222 9092 25228 9104
rect 25183 9064 25228 9092
rect 23569 9055 23627 9061
rect 25222 9052 25228 9064
rect 25280 9052 25286 9104
rect 6638 9024 6644 9036
rect 6599 8996 6644 9024
rect 6638 8984 6644 8996
rect 6696 8984 6702 9036
rect 11425 9027 11483 9033
rect 11425 8993 11437 9027
rect 11471 9024 11483 9027
rect 11882 9024 11888 9036
rect 11471 8996 11888 9024
rect 11471 8993 11483 8996
rect 11425 8987 11483 8993
rect 11882 8984 11888 8996
rect 11940 8984 11946 9036
rect 12250 8984 12256 9036
rect 12308 9024 12314 9036
rect 18598 9024 18604 9036
rect 12308 8996 18184 9024
rect 18559 8996 18604 9024
rect 12308 8984 12314 8996
rect 1854 8956 1860 8968
rect 1815 8928 1860 8956
rect 1854 8916 1860 8928
rect 1912 8916 1918 8968
rect 11330 8956 11336 8968
rect 11291 8928 11336 8956
rect 11330 8916 11336 8928
rect 11388 8916 11394 8968
rect 11514 8916 11520 8968
rect 11572 8956 11578 8968
rect 11977 8959 12035 8965
rect 11977 8956 11989 8959
rect 11572 8928 11989 8956
rect 11572 8916 11578 8928
rect 11977 8925 11989 8928
rect 12023 8956 12035 8959
rect 12434 8956 12440 8968
rect 12023 8928 12440 8956
rect 12023 8925 12035 8928
rect 11977 8919 12035 8925
rect 12434 8916 12440 8928
rect 12492 8916 12498 8968
rect 16574 8956 16580 8968
rect 16487 8928 16580 8956
rect 16574 8916 16580 8928
rect 16632 8916 16638 8968
rect 5994 8888 6000 8900
rect 5955 8860 6000 8888
rect 5994 8848 6000 8860
rect 6052 8848 6058 8900
rect 6089 8891 6147 8897
rect 6089 8857 6101 8891
rect 6135 8888 6147 8891
rect 6454 8888 6460 8900
rect 6135 8860 6460 8888
rect 6135 8857 6147 8860
rect 6089 8851 6147 8857
rect 6454 8848 6460 8860
rect 6512 8848 6518 8900
rect 8110 8848 8116 8900
rect 8168 8888 8174 8900
rect 11238 8888 11244 8900
rect 8168 8860 11244 8888
rect 8168 8848 8174 8860
rect 11238 8848 11244 8860
rect 11296 8848 11302 8900
rect 1949 8823 2007 8829
rect 1949 8789 1961 8823
rect 1995 8820 2007 8823
rect 8570 8820 8576 8832
rect 1995 8792 8576 8820
rect 1995 8789 2007 8792
rect 1949 8783 2007 8789
rect 8570 8780 8576 8792
rect 8628 8780 8634 8832
rect 11974 8780 11980 8832
rect 12032 8820 12038 8832
rect 12069 8823 12127 8829
rect 12069 8820 12081 8823
rect 12032 8792 12081 8820
rect 12032 8780 12038 8792
rect 12069 8789 12081 8792
rect 12115 8789 12127 8823
rect 16592 8820 16620 8916
rect 16850 8848 16856 8900
rect 16908 8888 16914 8900
rect 16908 8860 16953 8888
rect 16908 8848 16914 8860
rect 17862 8820 17868 8832
rect 16592 8792 17868 8820
rect 12069 8783 12127 8789
rect 17862 8780 17868 8792
rect 17920 8780 17926 8832
rect 17972 8820 18000 8942
rect 18156 8888 18184 8996
rect 18598 8984 18604 8996
rect 18656 8984 18662 9036
rect 25240 9024 25268 9052
rect 18708 8996 25268 9024
rect 18230 8916 18236 8968
rect 18288 8956 18294 8968
rect 18708 8956 18736 8996
rect 18288 8928 18736 8956
rect 18288 8916 18294 8928
rect 19334 8916 19340 8968
rect 19392 8956 19398 8968
rect 20162 8956 20168 8968
rect 19392 8928 20168 8956
rect 19392 8916 19398 8928
rect 20162 8916 20168 8928
rect 20220 8956 20226 8968
rect 20533 8959 20591 8965
rect 20533 8956 20545 8959
rect 20220 8928 20545 8956
rect 20220 8916 20226 8928
rect 20533 8925 20545 8928
rect 20579 8956 20591 8959
rect 20622 8956 20628 8968
rect 20579 8928 20628 8956
rect 20579 8925 20591 8928
rect 20533 8919 20591 8925
rect 20622 8916 20628 8928
rect 20680 8916 20686 8968
rect 21634 8956 21640 8968
rect 21547 8928 21640 8956
rect 21634 8916 21640 8928
rect 21692 8956 21698 8968
rect 21910 8956 21916 8968
rect 21692 8928 21916 8956
rect 21692 8916 21698 8928
rect 21910 8916 21916 8928
rect 21968 8916 21974 8968
rect 22554 8956 22560 8968
rect 22515 8928 22560 8956
rect 22554 8916 22560 8928
rect 22612 8916 22618 8968
rect 23477 8959 23535 8965
rect 23477 8925 23489 8959
rect 23523 8956 23535 8959
rect 23566 8956 23572 8968
rect 23523 8928 23572 8956
rect 23523 8925 23535 8928
rect 23477 8919 23535 8925
rect 23566 8916 23572 8928
rect 23624 8916 23630 8968
rect 25792 8965 25820 9132
rect 28718 9120 28724 9132
rect 28776 9120 28782 9172
rect 25777 8959 25835 8965
rect 25777 8925 25789 8959
rect 25823 8925 25835 8959
rect 25777 8919 25835 8925
rect 27982 8916 27988 8968
rect 28040 8956 28046 8968
rect 28169 8959 28227 8965
rect 28169 8956 28181 8959
rect 28040 8928 28181 8956
rect 28040 8916 28046 8928
rect 28169 8925 28181 8928
rect 28215 8925 28227 8959
rect 28626 8956 28632 8968
rect 28587 8928 28632 8956
rect 28169 8919 28227 8925
rect 28626 8916 28632 8928
rect 28684 8956 28690 8968
rect 29362 8956 29368 8968
rect 28684 8928 29368 8956
rect 28684 8916 28690 8928
rect 29362 8916 29368 8928
rect 29420 8916 29426 8968
rect 30558 8956 30564 8968
rect 30519 8928 30564 8956
rect 30558 8916 30564 8928
rect 30616 8916 30622 8968
rect 34790 8916 34796 8968
rect 34848 8956 34854 8968
rect 38013 8959 38071 8965
rect 38013 8956 38025 8959
rect 34848 8928 38025 8956
rect 34848 8916 34854 8928
rect 38013 8925 38025 8928
rect 38059 8925 38071 8959
rect 38013 8919 38071 8925
rect 22646 8888 22652 8900
rect 18156 8860 22652 8888
rect 22646 8848 22652 8860
rect 22704 8848 22710 8900
rect 22833 8891 22891 8897
rect 22833 8857 22845 8891
rect 22879 8888 22891 8891
rect 22879 8860 22913 8888
rect 22879 8857 22891 8860
rect 22833 8851 22891 8857
rect 20070 8820 20076 8832
rect 17972 8792 20076 8820
rect 20070 8780 20076 8792
rect 20128 8780 20134 8832
rect 20622 8820 20628 8832
rect 20583 8792 20628 8820
rect 20622 8780 20628 8792
rect 20680 8780 20686 8832
rect 20714 8780 20720 8832
rect 20772 8820 20778 8832
rect 21729 8823 21787 8829
rect 21729 8820 21741 8823
rect 20772 8792 21741 8820
rect 20772 8780 20778 8792
rect 21729 8789 21741 8792
rect 21775 8789 21787 8823
rect 21729 8783 21787 8789
rect 21818 8780 21824 8832
rect 21876 8820 21882 8832
rect 22848 8820 22876 8851
rect 23750 8848 23756 8900
rect 23808 8888 23814 8900
rect 24673 8891 24731 8897
rect 24673 8888 24685 8891
rect 23808 8860 24685 8888
rect 23808 8848 23814 8860
rect 24673 8857 24685 8860
rect 24719 8857 24731 8891
rect 24673 8851 24731 8857
rect 24765 8891 24823 8897
rect 24765 8857 24777 8891
rect 24811 8857 24823 8891
rect 24765 8851 24823 8857
rect 24210 8820 24216 8832
rect 21876 8792 24216 8820
rect 21876 8780 21882 8792
rect 24210 8780 24216 8792
rect 24268 8780 24274 8832
rect 24780 8820 24808 8851
rect 25869 8823 25927 8829
rect 25869 8820 25881 8823
rect 24780 8792 25881 8820
rect 25869 8789 25881 8792
rect 25915 8789 25927 8823
rect 25869 8783 25927 8789
rect 26513 8823 26571 8829
rect 26513 8789 26525 8823
rect 26559 8820 26571 8823
rect 27154 8820 27160 8832
rect 26559 8792 27160 8820
rect 26559 8789 26571 8792
rect 26513 8783 26571 8789
rect 27154 8780 27160 8792
rect 27212 8780 27218 8832
rect 27985 8823 28043 8829
rect 27985 8789 27997 8823
rect 28031 8820 28043 8823
rect 28442 8820 28448 8832
rect 28031 8792 28448 8820
rect 28031 8789 28043 8792
rect 27985 8783 28043 8789
rect 28442 8780 28448 8792
rect 28500 8780 28506 8832
rect 30653 8823 30711 8829
rect 30653 8789 30665 8823
rect 30699 8820 30711 8823
rect 32490 8820 32496 8832
rect 30699 8792 32496 8820
rect 30699 8789 30711 8792
rect 30653 8783 30711 8789
rect 32490 8780 32496 8792
rect 32548 8780 32554 8832
rect 38194 8820 38200 8832
rect 38155 8792 38200 8820
rect 38194 8780 38200 8792
rect 38252 8780 38258 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 2038 8616 2044 8628
rect 1999 8588 2044 8616
rect 2038 8576 2044 8588
rect 2096 8576 2102 8628
rect 8294 8616 8300 8628
rect 8207 8588 8300 8616
rect 8110 8548 8116 8560
rect 5198 8520 8116 8548
rect 8110 8508 8116 8520
rect 8168 8508 8174 8560
rect 1949 8483 2007 8489
rect 1949 8449 1961 8483
rect 1995 8480 2007 8483
rect 2314 8480 2320 8492
rect 1995 8452 2320 8480
rect 1995 8449 2007 8452
rect 1949 8443 2007 8449
rect 2314 8440 2320 8452
rect 2372 8440 2378 8492
rect 5721 8483 5779 8489
rect 5721 8449 5733 8483
rect 5767 8480 5779 8483
rect 6362 8480 6368 8492
rect 5767 8452 6368 8480
rect 5767 8449 5779 8452
rect 5721 8443 5779 8449
rect 6362 8440 6368 8452
rect 6420 8440 6426 8492
rect 8220 8489 8248 8588
rect 8294 8576 8300 8588
rect 8352 8616 8358 8628
rect 9214 8616 9220 8628
rect 8352 8588 9220 8616
rect 8352 8576 8358 8588
rect 9214 8576 9220 8588
rect 9272 8576 9278 8628
rect 9953 8619 10011 8625
rect 9953 8585 9965 8619
rect 9999 8616 10011 8619
rect 10134 8616 10140 8628
rect 9999 8588 10140 8616
rect 9999 8585 10011 8588
rect 9953 8579 10011 8585
rect 10134 8576 10140 8588
rect 10192 8576 10198 8628
rect 10502 8576 10508 8628
rect 10560 8616 10566 8628
rect 15105 8619 15163 8625
rect 15105 8616 15117 8619
rect 10560 8588 15117 8616
rect 10560 8576 10566 8588
rect 15105 8585 15117 8588
rect 15151 8585 15163 8619
rect 15105 8579 15163 8585
rect 15470 8576 15476 8628
rect 15528 8616 15534 8628
rect 15528 8588 15976 8616
rect 15528 8576 15534 8588
rect 8478 8548 8484 8560
rect 8439 8520 8484 8548
rect 8478 8508 8484 8520
rect 8536 8508 8542 8560
rect 11974 8548 11980 8560
rect 11935 8520 11980 8548
rect 11974 8508 11980 8520
rect 12032 8508 12038 8560
rect 12529 8551 12587 8557
rect 12529 8517 12541 8551
rect 12575 8548 12587 8551
rect 15838 8548 15844 8560
rect 12575 8520 15844 8548
rect 12575 8517 12587 8520
rect 12529 8511 12587 8517
rect 15838 8508 15844 8520
rect 15896 8508 15902 8560
rect 15948 8548 15976 8588
rect 16850 8576 16856 8628
rect 16908 8616 16914 8628
rect 18966 8616 18972 8628
rect 16908 8588 18972 8616
rect 16908 8576 16914 8588
rect 18966 8576 18972 8588
rect 19024 8616 19030 8628
rect 19702 8616 19708 8628
rect 19024 8588 19708 8616
rect 19024 8576 19030 8588
rect 19702 8576 19708 8588
rect 19760 8576 19766 8628
rect 20438 8576 20444 8628
rect 20496 8616 20502 8628
rect 20898 8616 20904 8628
rect 20496 8588 20904 8616
rect 20496 8576 20502 8588
rect 20898 8576 20904 8588
rect 20956 8576 20962 8628
rect 21082 8616 21088 8628
rect 21043 8588 21088 8616
rect 21082 8576 21088 8588
rect 21140 8576 21146 8628
rect 21928 8588 23244 8616
rect 18230 8548 18236 8560
rect 15948 8520 18236 8548
rect 18230 8508 18236 8520
rect 18288 8508 18294 8560
rect 19610 8548 19616 8560
rect 19550 8520 19616 8548
rect 19610 8508 19616 8520
rect 19668 8508 19674 8560
rect 8205 8483 8263 8489
rect 8205 8449 8217 8483
rect 8251 8449 8263 8483
rect 8205 8443 8263 8449
rect 9582 8440 9588 8492
rect 9640 8440 9646 8492
rect 15013 8483 15071 8489
rect 15013 8449 15025 8483
rect 15059 8449 15071 8483
rect 15013 8443 15071 8449
rect 3697 8415 3755 8421
rect 3697 8381 3709 8415
rect 3743 8381 3755 8415
rect 3697 8375 3755 8381
rect 3973 8415 4031 8421
rect 3973 8381 3985 8415
rect 4019 8412 4031 8415
rect 5810 8412 5816 8424
rect 4019 8384 5816 8412
rect 4019 8381 4031 8384
rect 3973 8375 4031 8381
rect 3712 8276 3740 8375
rect 5810 8372 5816 8384
rect 5868 8372 5874 8424
rect 8570 8372 8576 8424
rect 8628 8412 8634 8424
rect 11885 8415 11943 8421
rect 11885 8412 11897 8415
rect 8628 8384 11897 8412
rect 8628 8372 8634 8384
rect 11885 8381 11897 8384
rect 11931 8381 11943 8415
rect 15028 8412 15056 8443
rect 19794 8440 19800 8492
rect 19852 8480 19858 8492
rect 20346 8480 20352 8492
rect 19852 8452 20352 8480
rect 19852 8440 19858 8452
rect 20346 8440 20352 8452
rect 20404 8440 20410 8492
rect 20806 8440 20812 8492
rect 20864 8480 20870 8492
rect 20993 8483 21051 8489
rect 20993 8480 21005 8483
rect 20864 8452 21005 8480
rect 20864 8440 20870 8452
rect 20993 8449 21005 8452
rect 21039 8449 21051 8483
rect 20993 8443 21051 8449
rect 17862 8412 17868 8424
rect 11885 8375 11943 8381
rect 12406 8384 17868 8412
rect 11330 8304 11336 8356
rect 11388 8344 11394 8356
rect 12406 8344 12434 8384
rect 17862 8372 17868 8384
rect 17920 8372 17926 8424
rect 17954 8372 17960 8424
rect 18012 8412 18018 8424
rect 18049 8415 18107 8421
rect 18049 8412 18061 8415
rect 18012 8384 18061 8412
rect 18012 8372 18018 8384
rect 18049 8381 18061 8384
rect 18095 8381 18107 8415
rect 18325 8415 18383 8421
rect 18325 8412 18337 8415
rect 18049 8375 18107 8381
rect 18156 8384 18337 8412
rect 11388 8316 12434 8344
rect 11388 8304 11394 8316
rect 13906 8304 13912 8356
rect 13964 8344 13970 8356
rect 14458 8344 14464 8356
rect 13964 8316 14464 8344
rect 13964 8304 13970 8316
rect 14458 8304 14464 8316
rect 14516 8304 14522 8356
rect 16114 8304 16120 8356
rect 16172 8344 16178 8356
rect 18156 8344 18184 8384
rect 18325 8381 18337 8384
rect 18371 8412 18383 8415
rect 21928 8412 21956 8588
rect 22186 8508 22192 8560
rect 22244 8548 22250 8560
rect 22244 8520 22289 8548
rect 22244 8508 22250 8520
rect 22646 8508 22652 8560
rect 22704 8548 22710 8560
rect 23109 8551 23167 8557
rect 23109 8548 23121 8551
rect 22704 8520 23121 8548
rect 22704 8508 22710 8520
rect 23109 8517 23121 8520
rect 23155 8517 23167 8551
rect 23216 8548 23244 8588
rect 23382 8576 23388 8628
rect 23440 8616 23446 8628
rect 23842 8616 23848 8628
rect 23440 8588 23848 8616
rect 23440 8576 23446 8588
rect 23842 8576 23848 8588
rect 23900 8616 23906 8628
rect 23900 8588 29776 8616
rect 23900 8576 23906 8588
rect 24854 8548 24860 8560
rect 23216 8520 24860 8548
rect 23109 8511 23167 8517
rect 24854 8508 24860 8520
rect 24912 8508 24918 8560
rect 25958 8548 25964 8560
rect 25792 8520 25964 8548
rect 23566 8480 23572 8492
rect 23479 8452 23572 8480
rect 23566 8440 23572 8452
rect 23624 8480 23630 8492
rect 24026 8480 24032 8492
rect 23624 8452 24032 8480
rect 23624 8440 23630 8452
rect 24026 8440 24032 8452
rect 24084 8440 24090 8492
rect 25792 8480 25820 8520
rect 25958 8508 25964 8520
rect 26016 8508 26022 8560
rect 26053 8551 26111 8557
rect 26053 8517 26065 8551
rect 26099 8548 26111 8551
rect 26142 8548 26148 8560
rect 26099 8520 26148 8548
rect 26099 8517 26111 8520
rect 26053 8511 26111 8517
rect 26142 8508 26148 8520
rect 26200 8508 26206 8560
rect 26234 8508 26240 8560
rect 26292 8548 26298 8560
rect 29362 8548 29368 8560
rect 26292 8520 29368 8548
rect 26292 8508 26298 8520
rect 29362 8508 29368 8520
rect 29420 8508 29426 8560
rect 27154 8480 27160 8492
rect 24504 8452 25820 8480
rect 27115 8452 27160 8480
rect 18371 8384 19380 8412
rect 18371 8381 18383 8384
rect 18325 8375 18383 8381
rect 16172 8316 18184 8344
rect 19352 8344 19380 8384
rect 19628 8384 21956 8412
rect 22097 8415 22155 8421
rect 19628 8344 19656 8384
rect 22097 8381 22109 8415
rect 22143 8412 22155 8415
rect 24504 8412 24532 8452
rect 27154 8440 27160 8452
rect 27212 8440 27218 8492
rect 28442 8480 28448 8492
rect 28403 8452 28448 8480
rect 28442 8440 28448 8452
rect 28500 8440 28506 8492
rect 29748 8489 29776 8588
rect 30558 8548 30564 8560
rect 30519 8520 30564 8548
rect 30558 8508 30564 8520
rect 30616 8508 30622 8560
rect 31113 8551 31171 8557
rect 31113 8517 31125 8551
rect 31159 8548 31171 8551
rect 31202 8548 31208 8560
rect 31159 8520 31208 8548
rect 31159 8517 31171 8520
rect 31113 8511 31171 8517
rect 31202 8508 31208 8520
rect 31260 8508 31266 8560
rect 29089 8483 29147 8489
rect 29089 8449 29101 8483
rect 29135 8480 29147 8483
rect 29733 8483 29791 8489
rect 29135 8452 29592 8480
rect 29135 8449 29147 8452
rect 29089 8443 29147 8449
rect 24670 8412 24676 8424
rect 22143 8384 24532 8412
rect 24631 8384 24676 8412
rect 22143 8381 22155 8384
rect 22097 8375 22155 8381
rect 24670 8372 24676 8384
rect 24728 8372 24734 8424
rect 24854 8412 24860 8424
rect 24815 8384 24860 8412
rect 24854 8372 24860 8384
rect 24912 8372 24918 8424
rect 25961 8415 26019 8421
rect 25961 8381 25973 8415
rect 26007 8412 26019 8415
rect 26326 8412 26332 8424
rect 26007 8384 26332 8412
rect 26007 8381 26019 8384
rect 25961 8375 26019 8381
rect 26326 8372 26332 8384
rect 26384 8372 26390 8424
rect 27341 8415 27399 8421
rect 26436 8384 26740 8412
rect 19352 8316 19656 8344
rect 19720 8316 20024 8344
rect 16172 8304 16178 8316
rect 3970 8276 3976 8288
rect 3712 8248 3976 8276
rect 3970 8236 3976 8248
rect 4028 8236 4034 8288
rect 11054 8236 11060 8288
rect 11112 8276 11118 8288
rect 11790 8276 11796 8288
rect 11112 8248 11796 8276
rect 11112 8236 11118 8248
rect 11790 8236 11796 8248
rect 11848 8276 11854 8288
rect 13814 8276 13820 8288
rect 11848 8248 13820 8276
rect 11848 8236 11854 8248
rect 13814 8236 13820 8248
rect 13872 8236 13878 8288
rect 13998 8236 14004 8288
rect 14056 8276 14062 8288
rect 19720 8276 19748 8316
rect 14056 8248 19748 8276
rect 14056 8236 14062 8248
rect 19794 8236 19800 8288
rect 19852 8276 19858 8288
rect 19996 8276 20024 8316
rect 20162 8304 20168 8356
rect 20220 8344 20226 8356
rect 23566 8344 23572 8356
rect 20220 8316 22048 8344
rect 20220 8304 20226 8316
rect 21266 8276 21272 8288
rect 19852 8248 19897 8276
rect 19996 8248 21272 8276
rect 19852 8236 19858 8248
rect 21266 8236 21272 8248
rect 21324 8236 21330 8288
rect 22020 8276 22048 8316
rect 22112 8316 23572 8344
rect 22112 8276 22140 8316
rect 23566 8304 23572 8316
rect 23624 8304 23630 8356
rect 25038 8344 25044 8356
rect 24999 8316 25044 8344
rect 25038 8304 25044 8316
rect 25096 8344 25102 8356
rect 26436 8344 26464 8384
rect 25096 8316 26464 8344
rect 25096 8304 25102 8316
rect 26510 8304 26516 8356
rect 26568 8344 26574 8356
rect 26712 8344 26740 8384
rect 27341 8381 27353 8415
rect 27387 8412 27399 8415
rect 27387 8384 28948 8412
rect 27387 8381 27399 8384
rect 27341 8375 27399 8381
rect 28920 8353 28948 8384
rect 29564 8353 29592 8452
rect 29733 8449 29745 8483
rect 29779 8449 29791 8483
rect 32490 8480 32496 8492
rect 32451 8452 32496 8480
rect 29733 8443 29791 8449
rect 32490 8440 32496 8452
rect 32548 8440 32554 8492
rect 30469 8415 30527 8421
rect 30469 8381 30481 8415
rect 30515 8412 30527 8415
rect 31754 8412 31760 8424
rect 30515 8384 31760 8412
rect 30515 8381 30527 8384
rect 30469 8375 30527 8381
rect 31754 8372 31760 8384
rect 31812 8372 31818 8424
rect 27617 8347 27675 8353
rect 27617 8344 27629 8347
rect 26568 8316 26613 8344
rect 26712 8316 27629 8344
rect 26568 8304 26574 8316
rect 27617 8313 27629 8316
rect 27663 8313 27675 8347
rect 27617 8307 27675 8313
rect 28905 8347 28963 8353
rect 28905 8313 28917 8347
rect 28951 8313 28963 8347
rect 28905 8307 28963 8313
rect 29549 8347 29607 8353
rect 29549 8313 29561 8347
rect 29595 8313 29607 8347
rect 29549 8307 29607 8313
rect 32309 8347 32367 8353
rect 32309 8313 32321 8347
rect 32355 8344 32367 8347
rect 34422 8344 34428 8356
rect 32355 8316 34428 8344
rect 32355 8313 32367 8316
rect 32309 8307 32367 8313
rect 34422 8304 34428 8316
rect 34480 8304 34486 8356
rect 23658 8276 23664 8288
rect 22020 8248 22140 8276
rect 23619 8248 23664 8276
rect 23658 8236 23664 8248
rect 23716 8236 23722 8288
rect 28261 8279 28319 8285
rect 28261 8245 28273 8279
rect 28307 8276 28319 8279
rect 28442 8276 28448 8288
rect 28307 8248 28448 8276
rect 28307 8245 28319 8248
rect 28261 8239 28319 8245
rect 28442 8236 28448 8248
rect 28500 8236 28506 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 2406 8032 2412 8084
rect 2464 8072 2470 8084
rect 2593 8075 2651 8081
rect 2593 8072 2605 8075
rect 2464 8044 2605 8072
rect 2464 8032 2470 8044
rect 2593 8041 2605 8044
rect 2639 8041 2651 8075
rect 5718 8072 5724 8084
rect 5679 8044 5724 8072
rect 2593 8035 2651 8041
rect 5718 8032 5724 8044
rect 5776 8032 5782 8084
rect 10042 8032 10048 8084
rect 10100 8072 10106 8084
rect 10318 8072 10324 8084
rect 10100 8044 10324 8072
rect 10100 8032 10106 8044
rect 10318 8032 10324 8044
rect 10376 8072 10382 8084
rect 16025 8075 16083 8081
rect 16025 8072 16037 8075
rect 10376 8044 16037 8072
rect 10376 8032 10382 8044
rect 16025 8041 16037 8044
rect 16071 8041 16083 8075
rect 16025 8035 16083 8041
rect 18690 8032 18696 8084
rect 18748 8072 18754 8084
rect 19334 8072 19340 8084
rect 18748 8044 19340 8072
rect 18748 8032 18754 8044
rect 19334 8032 19340 8044
rect 19392 8032 19398 8084
rect 20070 8032 20076 8084
rect 20128 8072 20134 8084
rect 21821 8075 21879 8081
rect 21821 8072 21833 8075
rect 20128 8044 21833 8072
rect 20128 8032 20134 8044
rect 21821 8041 21833 8044
rect 21867 8041 21879 8075
rect 21821 8035 21879 8041
rect 22094 8032 22100 8084
rect 22152 8072 22158 8084
rect 22462 8072 22468 8084
rect 22152 8044 22324 8072
rect 22423 8044 22468 8072
rect 22152 8032 22158 8044
rect 5736 8004 5764 8032
rect 12897 8007 12955 8013
rect 5736 7976 6132 8004
rect 2041 7939 2099 7945
rect 2041 7905 2053 7939
rect 2087 7936 2099 7939
rect 5994 7936 6000 7948
rect 2087 7908 6000 7936
rect 2087 7905 2099 7908
rect 2041 7899 2099 7905
rect 5994 7896 6000 7908
rect 6052 7896 6058 7948
rect 6104 7936 6132 7976
rect 12897 7973 12909 8007
rect 12943 8004 12955 8007
rect 13722 8004 13728 8016
rect 12943 7976 13728 8004
rect 12943 7973 12955 7976
rect 12897 7967 12955 7973
rect 13722 7964 13728 7976
rect 13780 7964 13786 8016
rect 15580 7976 19564 8004
rect 6825 7939 6883 7945
rect 6825 7936 6837 7939
rect 6104 7908 6837 7936
rect 6825 7905 6837 7908
rect 6871 7905 6883 7939
rect 6825 7899 6883 7905
rect 8573 7939 8631 7945
rect 8573 7905 8585 7939
rect 8619 7936 8631 7939
rect 11054 7936 11060 7948
rect 8619 7908 11060 7936
rect 8619 7905 8631 7908
rect 8573 7899 8631 7905
rect 11054 7896 11060 7908
rect 11112 7896 11118 7948
rect 15580 7936 15608 7976
rect 12544 7908 15608 7936
rect 1854 7828 1860 7880
rect 1912 7868 1918 7880
rect 1949 7871 2007 7877
rect 1949 7868 1961 7871
rect 1912 7840 1961 7868
rect 1912 7828 1918 7840
rect 1949 7837 1961 7840
rect 1995 7837 2007 7871
rect 1949 7831 2007 7837
rect 2774 7828 2780 7880
rect 2832 7868 2838 7880
rect 3970 7868 3976 7880
rect 2832 7840 2877 7868
rect 3931 7840 3976 7868
rect 2832 7828 2838 7840
rect 3970 7828 3976 7840
rect 4028 7828 4034 7880
rect 6546 7868 6552 7880
rect 6507 7840 6552 7868
rect 6546 7828 6552 7840
rect 6604 7828 6610 7880
rect 11146 7868 11152 7880
rect 11107 7840 11152 7868
rect 11146 7828 11152 7840
rect 11204 7828 11210 7880
rect 12544 7854 12572 7908
rect 17954 7896 17960 7948
rect 18012 7936 18018 7948
rect 19429 7939 19487 7945
rect 19429 7936 19441 7939
rect 18012 7908 19441 7936
rect 18012 7896 18018 7908
rect 19429 7905 19441 7908
rect 19475 7905 19487 7939
rect 19536 7936 19564 7976
rect 20806 7964 20812 8016
rect 20864 8004 20870 8016
rect 20990 8004 20996 8016
rect 20864 7976 20996 8004
rect 20864 7964 20870 7976
rect 20990 7964 20996 7976
rect 21048 8004 21054 8016
rect 21177 8007 21235 8013
rect 21177 8004 21189 8007
rect 21048 7976 21189 8004
rect 21048 7964 21054 7976
rect 21177 7973 21189 7976
rect 21223 7973 21235 8007
rect 22296 8004 22324 8044
rect 22462 8032 22468 8044
rect 22520 8032 22526 8084
rect 23937 8075 23995 8081
rect 23937 8041 23949 8075
rect 23983 8072 23995 8075
rect 24854 8072 24860 8084
rect 23983 8044 24860 8072
rect 23983 8041 23995 8044
rect 23937 8035 23995 8041
rect 24854 8032 24860 8044
rect 24912 8032 24918 8084
rect 25961 8075 26019 8081
rect 25961 8041 25973 8075
rect 26007 8072 26019 8075
rect 26142 8072 26148 8084
rect 26007 8044 26148 8072
rect 26007 8041 26019 8044
rect 25961 8035 26019 8041
rect 26142 8032 26148 8044
rect 26200 8032 26206 8084
rect 29638 8032 29644 8084
rect 29696 8072 29702 8084
rect 29733 8075 29791 8081
rect 29733 8072 29745 8075
rect 29696 8044 29745 8072
rect 29696 8032 29702 8044
rect 29733 8041 29745 8044
rect 29779 8041 29791 8075
rect 29733 8035 29791 8041
rect 30377 8075 30435 8081
rect 30377 8041 30389 8075
rect 30423 8072 30435 8075
rect 30558 8072 30564 8084
rect 30423 8044 30564 8072
rect 30423 8041 30435 8044
rect 30377 8035 30435 8041
rect 30558 8032 30564 8044
rect 30616 8032 30622 8084
rect 31754 8072 31760 8084
rect 31715 8044 31760 8072
rect 31754 8032 31760 8044
rect 31812 8032 31818 8084
rect 22554 8004 22560 8016
rect 22296 7976 22560 8004
rect 21177 7967 21235 7973
rect 22554 7964 22560 7976
rect 22612 7964 22618 8016
rect 24581 8007 24639 8013
rect 24581 7973 24593 8007
rect 24627 7973 24639 8007
rect 24581 7967 24639 7973
rect 20714 7936 20720 7948
rect 19536 7908 20720 7936
rect 19429 7899 19487 7905
rect 20714 7896 20720 7908
rect 20772 7896 20778 7948
rect 24596 7936 24624 7967
rect 28258 7964 28264 8016
rect 28316 7964 28322 8016
rect 28276 7936 28304 7964
rect 28353 7939 28411 7945
rect 28353 7936 28365 7939
rect 24596 7908 25452 7936
rect 28276 7908 28365 7936
rect 14274 7868 14280 7880
rect 14235 7840 14280 7868
rect 14274 7828 14280 7840
rect 14332 7828 14338 7880
rect 18046 7828 18052 7880
rect 18104 7868 18110 7880
rect 18690 7868 18696 7880
rect 18104 7840 18696 7868
rect 18104 7828 18110 7840
rect 18690 7828 18696 7840
rect 18748 7828 18754 7880
rect 21729 7871 21787 7877
rect 21729 7837 21741 7871
rect 21775 7868 21787 7871
rect 21910 7868 21916 7880
rect 21775 7840 21916 7868
rect 21775 7837 21787 7840
rect 21729 7831 21787 7837
rect 21910 7828 21916 7840
rect 21968 7828 21974 7880
rect 22002 7828 22008 7880
rect 22060 7868 22066 7880
rect 22278 7868 22284 7880
rect 22060 7840 22284 7868
rect 22060 7828 22066 7840
rect 22278 7828 22284 7840
rect 22336 7868 22342 7880
rect 22373 7871 22431 7877
rect 22373 7868 22385 7871
rect 22336 7840 22385 7868
rect 22336 7828 22342 7840
rect 22373 7837 22385 7840
rect 22419 7837 22431 7871
rect 22373 7831 22431 7837
rect 22462 7828 22468 7880
rect 22520 7868 22526 7880
rect 22520 7840 23796 7868
rect 22520 7828 22526 7840
rect 4249 7803 4307 7809
rect 4249 7769 4261 7803
rect 4295 7800 4307 7803
rect 4522 7800 4528 7812
rect 4295 7772 4528 7800
rect 4295 7769 4307 7772
rect 4249 7763 4307 7769
rect 4522 7760 4528 7772
rect 4580 7760 4586 7812
rect 8478 7800 8484 7812
rect 5474 7772 7236 7800
rect 8050 7772 8484 7800
rect 7208 7732 7236 7772
rect 8478 7760 8484 7772
rect 8536 7760 8542 7812
rect 11330 7760 11336 7812
rect 11388 7800 11394 7812
rect 11425 7803 11483 7809
rect 11425 7800 11437 7803
rect 11388 7772 11437 7800
rect 11388 7760 11394 7772
rect 11425 7769 11437 7772
rect 11471 7769 11483 7803
rect 14553 7803 14611 7809
rect 14553 7800 14565 7803
rect 11425 7763 11483 7769
rect 12820 7772 14565 7800
rect 8662 7732 8668 7744
rect 7208 7704 8668 7732
rect 8662 7692 8668 7704
rect 8720 7692 8726 7744
rect 10594 7692 10600 7744
rect 10652 7732 10658 7744
rect 12820 7732 12848 7772
rect 14553 7769 14565 7772
rect 14599 7769 14611 7803
rect 14553 7763 14611 7769
rect 15194 7760 15200 7812
rect 15252 7760 15258 7812
rect 18230 7760 18236 7812
rect 18288 7800 18294 7812
rect 18288 7772 18920 7800
rect 18288 7760 18294 7772
rect 10652 7704 12848 7732
rect 10652 7692 10658 7704
rect 13814 7692 13820 7744
rect 13872 7732 13878 7744
rect 18322 7732 18328 7744
rect 13872 7704 18328 7732
rect 13872 7692 13878 7704
rect 18322 7692 18328 7704
rect 18380 7692 18386 7744
rect 18506 7692 18512 7744
rect 18564 7732 18570 7744
rect 18785 7735 18843 7741
rect 18785 7732 18797 7735
rect 18564 7704 18797 7732
rect 18564 7692 18570 7704
rect 18785 7701 18797 7704
rect 18831 7701 18843 7735
rect 18892 7732 18920 7772
rect 19334 7760 19340 7812
rect 19392 7800 19398 7812
rect 19610 7800 19616 7812
rect 19392 7772 19616 7800
rect 19392 7760 19398 7772
rect 19610 7760 19616 7772
rect 19668 7760 19674 7812
rect 19705 7803 19763 7809
rect 19705 7769 19717 7803
rect 19751 7800 19763 7803
rect 19794 7800 19800 7812
rect 19751 7772 19800 7800
rect 19751 7769 19763 7772
rect 19705 7763 19763 7769
rect 19794 7760 19800 7772
rect 19852 7760 19858 7812
rect 23658 7800 23664 7812
rect 20930 7772 23664 7800
rect 23658 7760 23664 7772
rect 23716 7760 23722 7812
rect 23768 7800 23796 7840
rect 23842 7828 23848 7880
rect 23900 7868 23906 7880
rect 24762 7868 24768 7880
rect 23900 7840 23945 7868
rect 24723 7840 24768 7868
rect 23900 7828 23906 7840
rect 24762 7828 24768 7840
rect 24820 7828 24826 7880
rect 25424 7877 25452 7908
rect 28353 7905 28365 7908
rect 28399 7905 28411 7939
rect 28626 7936 28632 7948
rect 28587 7908 28632 7936
rect 28353 7899 28411 7905
rect 28626 7896 28632 7908
rect 28684 7896 28690 7948
rect 25409 7871 25467 7877
rect 25409 7837 25421 7871
rect 25455 7837 25467 7871
rect 25409 7831 25467 7837
rect 25869 7871 25927 7877
rect 25869 7837 25881 7871
rect 25915 7868 25927 7871
rect 26881 7871 26939 7877
rect 26881 7868 26893 7871
rect 25915 7840 26893 7868
rect 25915 7837 25927 7840
rect 25869 7831 25927 7837
rect 26881 7837 26893 7840
rect 26927 7837 26939 7871
rect 26881 7831 26939 7837
rect 29917 7871 29975 7877
rect 29917 7837 29929 7871
rect 29963 7837 29975 7871
rect 29917 7831 29975 7837
rect 25884 7800 25912 7831
rect 23768 7772 25912 7800
rect 28442 7760 28448 7812
rect 28500 7800 28506 7812
rect 28500 7772 28545 7800
rect 28500 7760 28506 7772
rect 28718 7760 28724 7812
rect 28776 7800 28782 7812
rect 29932 7800 29960 7831
rect 30374 7828 30380 7880
rect 30432 7868 30438 7880
rect 30561 7871 30619 7877
rect 30561 7868 30573 7871
rect 30432 7840 30573 7868
rect 30432 7828 30438 7840
rect 30561 7837 30573 7840
rect 30607 7837 30619 7871
rect 30561 7831 30619 7837
rect 31665 7871 31723 7877
rect 31665 7837 31677 7871
rect 31711 7868 31723 7871
rect 33042 7868 33048 7880
rect 31711 7840 33048 7868
rect 31711 7837 31723 7840
rect 31665 7831 31723 7837
rect 33042 7828 33048 7840
rect 33100 7828 33106 7880
rect 38286 7868 38292 7880
rect 38247 7840 38292 7868
rect 38286 7828 38292 7840
rect 38344 7828 38350 7880
rect 28776 7772 29960 7800
rect 28776 7760 28782 7772
rect 22370 7732 22376 7744
rect 18892 7704 22376 7732
rect 18785 7695 18843 7701
rect 22370 7692 22376 7704
rect 22428 7692 22434 7744
rect 23566 7692 23572 7744
rect 23624 7732 23630 7744
rect 25225 7735 25283 7741
rect 25225 7732 25237 7735
rect 23624 7704 25237 7732
rect 23624 7692 23630 7704
rect 25225 7701 25237 7704
rect 25271 7701 25283 7735
rect 25225 7695 25283 7701
rect 26697 7735 26755 7741
rect 26697 7701 26709 7735
rect 26743 7732 26755 7735
rect 27338 7732 27344 7744
rect 26743 7704 27344 7732
rect 26743 7701 26755 7704
rect 26697 7695 26755 7701
rect 27338 7692 27344 7704
rect 27396 7692 27402 7744
rect 37274 7692 37280 7744
rect 37332 7732 37338 7744
rect 38105 7735 38163 7741
rect 38105 7732 38117 7735
rect 37332 7704 38117 7732
rect 37332 7692 37338 7704
rect 38105 7701 38117 7704
rect 38151 7701 38163 7735
rect 38105 7695 38163 7701
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 2041 7531 2099 7537
rect 2041 7497 2053 7531
rect 2087 7528 2099 7531
rect 6086 7528 6092 7540
rect 2087 7500 6092 7528
rect 2087 7497 2099 7500
rect 2041 7491 2099 7497
rect 6086 7488 6092 7500
rect 6144 7488 6150 7540
rect 8202 7488 8208 7540
rect 8260 7488 8266 7540
rect 8478 7488 8484 7540
rect 8536 7528 8542 7540
rect 13998 7528 14004 7540
rect 8536 7500 14004 7528
rect 8536 7488 8542 7500
rect 13998 7488 14004 7500
rect 14056 7488 14062 7540
rect 18322 7528 18328 7540
rect 14108 7500 18328 7528
rect 6546 7420 6552 7472
rect 6604 7460 6610 7472
rect 8220 7460 8248 7488
rect 9306 7460 9312 7472
rect 6604 7432 8248 7460
rect 9062 7432 9312 7460
rect 6604 7420 6610 7432
rect 1670 7352 1676 7404
rect 1728 7392 1734 7404
rect 7576 7401 7604 7432
rect 9306 7420 9312 7432
rect 9364 7420 9370 7472
rect 9398 7420 9404 7472
rect 9456 7460 9462 7472
rect 13906 7460 13912 7472
rect 9456 7432 13912 7460
rect 9456 7420 9462 7432
rect 13906 7420 13912 7432
rect 13964 7420 13970 7472
rect 1949 7395 2007 7401
rect 1949 7392 1961 7395
rect 1728 7364 1961 7392
rect 1728 7352 1734 7364
rect 1949 7361 1961 7364
rect 1995 7361 2007 7395
rect 1949 7355 2007 7361
rect 7561 7395 7619 7401
rect 7561 7361 7573 7395
rect 7607 7361 7619 7395
rect 7561 7355 7619 7361
rect 7834 7324 7840 7336
rect 7795 7296 7840 7324
rect 7834 7284 7840 7296
rect 7892 7284 7898 7336
rect 9582 7284 9588 7336
rect 9640 7324 9646 7336
rect 14108 7324 14136 7500
rect 18322 7488 18328 7500
rect 18380 7488 18386 7540
rect 22741 7531 22799 7537
rect 22741 7528 22753 7531
rect 18616 7500 22753 7528
rect 14550 7460 14556 7472
rect 14511 7432 14556 7460
rect 14550 7420 14556 7432
rect 14608 7420 14614 7472
rect 18616 7460 18644 7500
rect 22741 7497 22753 7500
rect 22787 7497 22799 7531
rect 27157 7531 27215 7537
rect 27157 7528 27169 7531
rect 22741 7491 22799 7497
rect 24872 7500 27169 7528
rect 21361 7463 21419 7469
rect 21361 7460 21373 7463
rect 15778 7432 18644 7460
rect 19458 7432 21373 7460
rect 21361 7429 21373 7432
rect 21407 7429 21419 7463
rect 21361 7423 21419 7429
rect 21450 7420 21456 7472
rect 21508 7460 21514 7472
rect 23566 7460 23572 7472
rect 21508 7432 23572 7460
rect 21508 7420 21514 7432
rect 23566 7420 23572 7432
rect 23624 7420 23630 7472
rect 24394 7420 24400 7472
rect 24452 7460 24458 7472
rect 24872 7469 24900 7500
rect 27157 7497 27169 7500
rect 27203 7497 27215 7531
rect 27157 7491 27215 7497
rect 24765 7463 24823 7469
rect 24765 7460 24777 7463
rect 24452 7432 24777 7460
rect 24452 7420 24458 7432
rect 24765 7429 24777 7432
rect 24811 7429 24823 7463
rect 24765 7423 24823 7429
rect 24857 7463 24915 7469
rect 24857 7429 24869 7463
rect 24903 7429 24915 7463
rect 29178 7460 29184 7472
rect 29139 7432 29184 7460
rect 24857 7423 24915 7429
rect 29178 7420 29184 7432
rect 29236 7420 29242 7472
rect 19444 7364 20116 7392
rect 14274 7324 14280 7336
rect 9640 7296 14136 7324
rect 14235 7296 14280 7324
rect 9640 7284 9646 7296
rect 14274 7284 14280 7296
rect 14332 7284 14338 7336
rect 15102 7324 15108 7336
rect 14384 7296 15108 7324
rect 13814 7216 13820 7268
rect 13872 7256 13878 7268
rect 14384 7256 14412 7296
rect 15102 7284 15108 7296
rect 15160 7284 15166 7336
rect 15562 7284 15568 7336
rect 15620 7324 15626 7336
rect 16298 7324 16304 7336
rect 15620 7296 16304 7324
rect 15620 7284 15626 7296
rect 16298 7284 16304 7296
rect 16356 7284 16362 7336
rect 17954 7324 17960 7336
rect 17915 7296 17960 7324
rect 17954 7284 17960 7296
rect 18012 7284 18018 7336
rect 18230 7324 18236 7336
rect 18191 7296 18236 7324
rect 18230 7284 18236 7296
rect 18288 7284 18294 7336
rect 18322 7284 18328 7336
rect 18380 7324 18386 7336
rect 19444 7324 19472 7364
rect 18380 7296 19472 7324
rect 18380 7284 18386 7296
rect 19886 7284 19892 7336
rect 19944 7324 19950 7336
rect 19981 7327 20039 7333
rect 19981 7324 19993 7327
rect 19944 7296 19993 7324
rect 19944 7284 19950 7296
rect 19981 7293 19993 7296
rect 20027 7293 20039 7327
rect 20088 7324 20116 7364
rect 21082 7352 21088 7404
rect 21140 7392 21146 7404
rect 21269 7395 21327 7401
rect 21269 7392 21281 7395
rect 21140 7364 21281 7392
rect 21140 7352 21146 7364
rect 21269 7361 21281 7364
rect 21315 7392 21327 7395
rect 21726 7392 21732 7404
rect 21315 7364 21732 7392
rect 21315 7361 21327 7364
rect 21269 7355 21327 7361
rect 21726 7352 21732 7364
rect 21784 7352 21790 7404
rect 22002 7392 22008 7404
rect 21963 7364 22008 7392
rect 22002 7352 22008 7364
rect 22060 7392 22066 7404
rect 22649 7395 22707 7401
rect 22649 7392 22661 7395
rect 22060 7364 22661 7392
rect 22060 7352 22066 7364
rect 22649 7361 22661 7364
rect 22695 7361 22707 7395
rect 22649 7355 22707 7361
rect 23477 7395 23535 7401
rect 23477 7361 23489 7395
rect 23523 7392 23535 7395
rect 23658 7392 23664 7404
rect 23523 7364 23664 7392
rect 23523 7361 23535 7364
rect 23477 7355 23535 7361
rect 23658 7352 23664 7364
rect 23716 7392 23722 7404
rect 24026 7392 24032 7404
rect 23716 7364 24032 7392
rect 23716 7352 23722 7364
rect 24026 7352 24032 7364
rect 24084 7352 24090 7404
rect 27338 7392 27344 7404
rect 27299 7364 27344 7392
rect 27338 7352 27344 7364
rect 27396 7352 27402 7404
rect 30190 7392 30196 7404
rect 30151 7364 30196 7392
rect 30190 7352 30196 7364
rect 30248 7352 30254 7404
rect 20088 7296 21588 7324
rect 19981 7287 20039 7293
rect 21560 7256 21588 7296
rect 21634 7284 21640 7336
rect 21692 7324 21698 7336
rect 25409 7327 25467 7333
rect 21692 7296 24716 7324
rect 21692 7284 21698 7296
rect 22097 7259 22155 7265
rect 22097 7256 22109 7259
rect 13872 7228 14412 7256
rect 19260 7228 21496 7256
rect 21560 7228 22109 7256
rect 13872 7216 13878 7228
rect 9309 7191 9367 7197
rect 9309 7157 9321 7191
rect 9355 7188 9367 7191
rect 11054 7188 11060 7200
rect 9355 7160 11060 7188
rect 9355 7157 9367 7160
rect 9309 7151 9367 7157
rect 11054 7148 11060 7160
rect 11112 7148 11118 7200
rect 12066 7148 12072 7200
rect 12124 7188 12130 7200
rect 19260 7188 19288 7228
rect 12124 7160 19288 7188
rect 21468 7188 21496 7228
rect 22097 7225 22109 7228
rect 22143 7225 22155 7259
rect 22097 7219 22155 7225
rect 23474 7216 23480 7268
rect 23532 7256 23538 7268
rect 23569 7259 23627 7265
rect 23569 7256 23581 7259
rect 23532 7228 23581 7256
rect 23532 7216 23538 7228
rect 23569 7225 23581 7228
rect 23615 7225 23627 7259
rect 24688 7256 24716 7296
rect 25409 7293 25421 7327
rect 25455 7324 25467 7327
rect 26510 7324 26516 7336
rect 25455 7296 26516 7324
rect 25455 7293 25467 7296
rect 25409 7287 25467 7293
rect 26510 7284 26516 7296
rect 26568 7284 26574 7336
rect 29086 7324 29092 7336
rect 29047 7296 29092 7324
rect 29086 7284 29092 7296
rect 29144 7284 29150 7336
rect 29362 7324 29368 7336
rect 29323 7296 29368 7324
rect 29362 7284 29368 7296
rect 29420 7284 29426 7336
rect 27246 7256 27252 7268
rect 24688 7228 27252 7256
rect 23569 7219 23627 7225
rect 27246 7216 27252 7228
rect 27304 7216 27310 7268
rect 24762 7188 24768 7200
rect 21468 7160 24768 7188
rect 12124 7148 12130 7160
rect 24762 7148 24768 7160
rect 24820 7148 24826 7200
rect 30285 7191 30343 7197
rect 30285 7157 30297 7191
rect 30331 7188 30343 7191
rect 31202 7188 31208 7200
rect 30331 7160 31208 7188
rect 30331 7157 30343 7160
rect 30285 7151 30343 7157
rect 31202 7148 31208 7160
rect 31260 7148 31266 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 6352 6987 6410 6993
rect 6352 6953 6364 6987
rect 6398 6984 6410 6987
rect 9398 6984 9404 6996
rect 6398 6956 9404 6984
rect 6398 6953 6410 6956
rect 6352 6947 6410 6953
rect 9398 6944 9404 6956
rect 9456 6944 9462 6996
rect 10124 6987 10182 6993
rect 10124 6953 10136 6987
rect 10170 6984 10182 6987
rect 19886 6984 19892 6996
rect 10170 6956 19892 6984
rect 10170 6953 10182 6956
rect 10124 6947 10182 6953
rect 19886 6944 19892 6956
rect 19944 6984 19950 6996
rect 21634 6984 21640 6996
rect 19944 6956 21640 6984
rect 19944 6944 19950 6956
rect 21634 6944 21640 6956
rect 21692 6944 21698 6996
rect 21726 6944 21732 6996
rect 21784 6984 21790 6996
rect 25590 6984 25596 6996
rect 21784 6956 25596 6984
rect 21784 6944 21790 6956
rect 25590 6944 25596 6956
rect 25648 6944 25654 6996
rect 11330 6876 11336 6928
rect 11388 6916 11394 6928
rect 13814 6916 13820 6928
rect 11388 6888 13820 6916
rect 11388 6876 11394 6888
rect 13814 6876 13820 6888
rect 13872 6876 13878 6928
rect 13906 6876 13912 6928
rect 13964 6916 13970 6928
rect 14642 6916 14648 6928
rect 13964 6888 14648 6916
rect 13964 6876 13970 6888
rect 14642 6876 14648 6888
rect 14700 6876 14706 6928
rect 16574 6876 16580 6928
rect 16632 6916 16638 6928
rect 20622 6916 20628 6928
rect 16632 6888 20628 6916
rect 16632 6876 16638 6888
rect 20622 6876 20628 6888
rect 20680 6876 20686 6928
rect 21542 6916 21548 6928
rect 21503 6888 21548 6916
rect 21542 6876 21548 6888
rect 21600 6876 21606 6928
rect 23290 6916 23296 6928
rect 22572 6888 23296 6916
rect 6089 6851 6147 6857
rect 2240 6820 6040 6848
rect 2240 6789 2268 6820
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6749 2283 6783
rect 2225 6743 2283 6749
rect 2317 6783 2375 6789
rect 2317 6749 2329 6783
rect 2363 6780 2375 6783
rect 2961 6783 3019 6789
rect 2961 6780 2973 6783
rect 2363 6752 2973 6780
rect 2363 6749 2375 6752
rect 2317 6743 2375 6749
rect 2961 6749 2973 6752
rect 3007 6749 3019 6783
rect 2961 6743 3019 6749
rect 2777 6647 2835 6653
rect 2777 6613 2789 6647
rect 2823 6644 2835 6647
rect 2866 6644 2872 6656
rect 2823 6616 2872 6644
rect 2823 6613 2835 6616
rect 2777 6607 2835 6613
rect 2866 6604 2872 6616
rect 2924 6604 2930 6656
rect 6012 6644 6040 6820
rect 6089 6817 6101 6851
rect 6135 6848 6147 6851
rect 6454 6848 6460 6860
rect 6135 6820 6460 6848
rect 6135 6817 6147 6820
rect 6089 6811 6147 6817
rect 6454 6808 6460 6820
rect 6512 6808 6518 6860
rect 10502 6848 10508 6860
rect 7484 6820 10508 6848
rect 7484 6766 7512 6820
rect 10502 6808 10508 6820
rect 10560 6808 10566 6860
rect 11609 6851 11667 6857
rect 11609 6817 11621 6851
rect 11655 6848 11667 6851
rect 11698 6848 11704 6860
rect 11655 6820 11704 6848
rect 11655 6817 11667 6820
rect 11609 6811 11667 6817
rect 11698 6808 11704 6820
rect 11756 6808 11762 6860
rect 17218 6808 17224 6860
rect 17276 6848 17282 6860
rect 22572 6857 22600 6888
rect 23290 6876 23296 6888
rect 23348 6876 23354 6928
rect 22558 6851 22616 6857
rect 17276 6820 22094 6848
rect 17276 6808 17282 6820
rect 9214 6740 9220 6792
rect 9272 6780 9278 6792
rect 9861 6783 9919 6789
rect 9861 6780 9873 6783
rect 9272 6752 9873 6780
rect 9272 6740 9278 6752
rect 9861 6749 9873 6752
rect 9907 6749 9919 6783
rect 9861 6743 9919 6749
rect 11422 6740 11428 6792
rect 11480 6780 11486 6792
rect 18230 6780 18236 6792
rect 11480 6752 18236 6780
rect 11480 6740 11486 6752
rect 18230 6740 18236 6752
rect 18288 6740 18294 6792
rect 19058 6740 19064 6792
rect 19116 6780 19122 6792
rect 20809 6783 20867 6789
rect 20809 6780 20821 6783
rect 19116 6752 20821 6780
rect 19116 6740 19122 6752
rect 20809 6749 20821 6752
rect 20855 6749 20867 6783
rect 20809 6743 20867 6749
rect 21453 6783 21511 6789
rect 21453 6749 21465 6783
rect 21499 6780 21511 6783
rect 21910 6780 21916 6792
rect 21499 6752 21916 6780
rect 21499 6749 21511 6752
rect 21453 6743 21511 6749
rect 21910 6740 21916 6752
rect 21968 6740 21974 6792
rect 22066 6780 22094 6820
rect 22558 6817 22570 6851
rect 22604 6817 22616 6851
rect 22558 6811 22616 6817
rect 28813 6851 28871 6857
rect 28813 6817 28825 6851
rect 28859 6848 28871 6851
rect 29178 6848 29184 6860
rect 28859 6820 29184 6848
rect 28859 6817 28871 6820
rect 28813 6811 28871 6817
rect 29178 6808 29184 6820
rect 29236 6808 29242 6860
rect 22373 6783 22431 6789
rect 22373 6780 22385 6783
rect 22066 6752 22385 6780
rect 22373 6749 22385 6752
rect 22419 6780 22431 6783
rect 23198 6780 23204 6792
rect 22419 6774 22508 6780
rect 22664 6774 23204 6780
rect 22419 6752 23204 6774
rect 22419 6749 22431 6752
rect 22373 6743 22431 6749
rect 22480 6746 22692 6752
rect 23198 6740 23204 6752
rect 23256 6740 23262 6792
rect 23382 6740 23388 6792
rect 23440 6780 23446 6792
rect 23477 6783 23535 6789
rect 23477 6780 23489 6783
rect 23440 6752 23489 6780
rect 23440 6740 23446 6752
rect 23477 6749 23489 6752
rect 23523 6749 23535 6783
rect 28718 6780 28724 6792
rect 28679 6752 28724 6780
rect 23477 6743 23535 6749
rect 28718 6740 28724 6752
rect 28776 6740 28782 6792
rect 9582 6712 9588 6724
rect 7668 6684 9588 6712
rect 7668 6644 7696 6684
rect 9582 6672 9588 6684
rect 9640 6672 9646 6724
rect 23569 6715 23627 6721
rect 23569 6712 23581 6715
rect 11362 6684 22508 6712
rect 7834 6644 7840 6656
rect 6012 6616 7696 6644
rect 7795 6616 7840 6644
rect 7834 6604 7840 6616
rect 7892 6604 7898 6656
rect 7926 6604 7932 6656
rect 7984 6644 7990 6656
rect 17218 6644 17224 6656
rect 7984 6616 17224 6644
rect 7984 6604 7990 6616
rect 17218 6604 17224 6616
rect 17276 6604 17282 6656
rect 17770 6604 17776 6656
rect 17828 6644 17834 6656
rect 20806 6644 20812 6656
rect 17828 6616 20812 6644
rect 17828 6604 17834 6616
rect 20806 6604 20812 6616
rect 20864 6604 20870 6656
rect 20901 6647 20959 6653
rect 20901 6613 20913 6647
rect 20947 6644 20959 6647
rect 22186 6644 22192 6656
rect 20947 6616 22192 6644
rect 20947 6613 20959 6616
rect 20901 6607 20959 6613
rect 22186 6604 22192 6616
rect 22244 6604 22250 6656
rect 22480 6644 22508 6684
rect 22664 6684 23581 6712
rect 22664 6644 22692 6684
rect 23569 6681 23581 6684
rect 23615 6681 23627 6715
rect 23569 6675 23627 6681
rect 22480 6616 22692 6644
rect 23017 6647 23075 6653
rect 23017 6613 23029 6647
rect 23063 6644 23075 6647
rect 25682 6644 25688 6656
rect 23063 6616 25688 6644
rect 23063 6613 23075 6616
rect 23017 6607 23075 6613
rect 25682 6604 25688 6616
rect 25740 6604 25746 6656
rect 25958 6604 25964 6656
rect 26016 6644 26022 6656
rect 28902 6644 28908 6656
rect 26016 6616 28908 6644
rect 26016 6604 26022 6616
rect 28902 6604 28908 6616
rect 28960 6604 28966 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 2041 6443 2099 6449
rect 2041 6409 2053 6443
rect 2087 6440 2099 6443
rect 7926 6440 7932 6452
rect 2087 6412 7932 6440
rect 2087 6409 2099 6412
rect 2041 6403 2099 6409
rect 7926 6400 7932 6412
rect 7984 6400 7990 6452
rect 10410 6440 10416 6452
rect 10371 6412 10416 6440
rect 10410 6400 10416 6412
rect 10468 6400 10474 6452
rect 10502 6400 10508 6452
rect 10560 6440 10566 6452
rect 16574 6440 16580 6452
rect 10560 6412 16580 6440
rect 10560 6400 10566 6412
rect 16574 6400 16580 6412
rect 16632 6400 16638 6452
rect 16666 6400 16672 6452
rect 16724 6440 16730 6452
rect 19334 6440 19340 6452
rect 16724 6412 19340 6440
rect 16724 6400 16730 6412
rect 19334 6400 19340 6412
rect 19392 6400 19398 6452
rect 19978 6440 19984 6452
rect 19939 6412 19984 6440
rect 19978 6400 19984 6412
rect 20036 6400 20042 6452
rect 20254 6400 20260 6452
rect 20312 6440 20318 6452
rect 23014 6440 23020 6452
rect 20312 6412 23020 6440
rect 20312 6400 20318 6412
rect 23014 6400 23020 6412
rect 23072 6400 23078 6452
rect 24305 6443 24363 6449
rect 24305 6440 24317 6443
rect 23124 6412 24317 6440
rect 23124 6372 23152 6412
rect 24305 6409 24317 6412
rect 24351 6409 24363 6443
rect 30834 6440 30840 6452
rect 24305 6403 24363 6409
rect 27264 6412 30840 6440
rect 10166 6344 23152 6372
rect 23198 6332 23204 6384
rect 23256 6372 23262 6384
rect 23256 6344 23301 6372
rect 23256 6332 23262 6344
rect 23566 6332 23572 6384
rect 23624 6372 23630 6384
rect 23753 6375 23811 6381
rect 23753 6372 23765 6375
rect 23624 6344 23765 6372
rect 23624 6332 23630 6344
rect 23753 6341 23765 6344
rect 23799 6372 23811 6375
rect 24118 6372 24124 6384
rect 23799 6344 24124 6372
rect 23799 6341 23811 6344
rect 23753 6335 23811 6341
rect 24118 6332 24124 6344
rect 24176 6332 24182 6384
rect 25314 6372 25320 6384
rect 25275 6344 25320 6372
rect 25314 6332 25320 6344
rect 25372 6332 25378 6384
rect 25869 6375 25927 6381
rect 25869 6341 25881 6375
rect 25915 6372 25927 6375
rect 25958 6372 25964 6384
rect 25915 6344 25964 6372
rect 25915 6341 25927 6344
rect 25869 6335 25927 6341
rect 25958 6332 25964 6344
rect 26016 6332 26022 6384
rect 27264 6381 27292 6412
rect 30834 6400 30840 6412
rect 30892 6440 30898 6452
rect 31297 6443 31355 6449
rect 31297 6440 31309 6443
rect 30892 6412 31309 6440
rect 30892 6400 30898 6412
rect 31297 6409 31309 6412
rect 31343 6409 31355 6443
rect 31297 6403 31355 6409
rect 27249 6375 27307 6381
rect 27249 6341 27261 6375
rect 27295 6341 27307 6375
rect 27249 6335 27307 6341
rect 27341 6375 27399 6381
rect 27341 6341 27353 6375
rect 27387 6372 27399 6375
rect 27614 6372 27620 6384
rect 27387 6344 27620 6372
rect 27387 6341 27399 6344
rect 27341 6335 27399 6341
rect 27614 6332 27620 6344
rect 27672 6332 27678 6384
rect 28537 6375 28595 6381
rect 28537 6341 28549 6375
rect 28583 6372 28595 6375
rect 28810 6372 28816 6384
rect 28583 6344 28816 6372
rect 28583 6341 28595 6344
rect 28537 6335 28595 6341
rect 28810 6332 28816 6344
rect 28868 6332 28874 6384
rect 28902 6332 28908 6384
rect 28960 6372 28966 6384
rect 29089 6375 29147 6381
rect 29089 6372 29101 6375
rect 28960 6344 29101 6372
rect 28960 6332 28966 6344
rect 29089 6341 29101 6344
rect 29135 6372 29147 6375
rect 30374 6372 30380 6384
rect 29135 6344 30380 6372
rect 29135 6341 29147 6344
rect 29089 6335 29147 6341
rect 30374 6332 30380 6344
rect 30432 6332 30438 6384
rect 1946 6304 1952 6316
rect 1907 6276 1952 6304
rect 1946 6264 1952 6276
rect 2004 6264 2010 6316
rect 5350 6264 5356 6316
rect 5408 6264 5414 6316
rect 19061 6307 19119 6313
rect 18064 6276 18276 6304
rect 3970 6236 3976 6248
rect 3931 6208 3976 6236
rect 3970 6196 3976 6208
rect 4028 6196 4034 6248
rect 4249 6239 4307 6245
rect 4249 6205 4261 6239
rect 4295 6236 4307 6239
rect 5902 6236 5908 6248
rect 4295 6208 5908 6236
rect 4295 6205 4307 6208
rect 4249 6199 4307 6205
rect 5902 6196 5908 6208
rect 5960 6196 5966 6248
rect 8665 6239 8723 6245
rect 8665 6205 8677 6239
rect 8711 6205 8723 6239
rect 8665 6199 8723 6205
rect 8941 6239 8999 6245
rect 8941 6205 8953 6239
rect 8987 6236 8999 6239
rect 9490 6236 9496 6248
rect 8987 6208 9496 6236
rect 8987 6205 8999 6208
rect 8941 6199 8999 6205
rect 5718 6168 5724 6180
rect 5631 6140 5724 6168
rect 5718 6128 5724 6140
rect 5776 6168 5782 6180
rect 7190 6168 7196 6180
rect 5776 6140 7196 6168
rect 5776 6128 5782 6140
rect 7190 6128 7196 6140
rect 7248 6128 7254 6180
rect 8680 6100 8708 6199
rect 9490 6196 9496 6208
rect 9548 6196 9554 6248
rect 9582 6196 9588 6248
rect 9640 6236 9646 6248
rect 12802 6236 12808 6248
rect 9640 6208 12808 6236
rect 9640 6196 9646 6208
rect 12802 6196 12808 6208
rect 12860 6196 12866 6248
rect 15286 6196 15292 6248
rect 15344 6236 15350 6248
rect 17957 6239 18015 6245
rect 17957 6236 17969 6239
rect 15344 6208 17969 6236
rect 15344 6196 15350 6208
rect 17957 6205 17969 6208
rect 18003 6205 18015 6239
rect 17957 6199 18015 6205
rect 10686 6128 10692 6180
rect 10744 6168 10750 6180
rect 16666 6168 16672 6180
rect 10744 6140 16672 6168
rect 10744 6128 10750 6140
rect 16666 6128 16672 6140
rect 16724 6128 16730 6180
rect 9122 6100 9128 6112
rect 8680 6072 9128 6100
rect 9122 6060 9128 6072
rect 9180 6060 9186 6112
rect 9306 6060 9312 6112
rect 9364 6100 9370 6112
rect 18064 6100 18092 6276
rect 18141 6239 18199 6245
rect 18141 6205 18153 6239
rect 18187 6205 18199 6239
rect 18248 6236 18276 6276
rect 19061 6273 19073 6307
rect 19107 6304 19119 6307
rect 19242 6304 19248 6316
rect 19107 6276 19248 6304
rect 19107 6273 19119 6276
rect 19061 6267 19119 6273
rect 19242 6264 19248 6276
rect 19300 6264 19306 6316
rect 19886 6304 19892 6316
rect 19847 6276 19892 6304
rect 19886 6264 19892 6276
rect 19944 6264 19950 6316
rect 21450 6304 21456 6316
rect 20732 6276 21456 6304
rect 20732 6236 20760 6276
rect 21450 6264 21456 6276
rect 21508 6264 21514 6316
rect 22002 6304 22008 6316
rect 21963 6276 22008 6304
rect 22002 6264 22008 6276
rect 22060 6264 22066 6316
rect 24210 6304 24216 6316
rect 24171 6276 24216 6304
rect 24210 6264 24216 6276
rect 24268 6264 24274 6316
rect 30006 6264 30012 6316
rect 30064 6304 30070 6316
rect 30193 6307 30251 6313
rect 30193 6304 30205 6307
rect 30064 6276 30205 6304
rect 30064 6264 30070 6276
rect 30193 6273 30205 6276
rect 30239 6273 30251 6307
rect 38286 6304 38292 6316
rect 38247 6276 38292 6304
rect 30193 6267 30251 6273
rect 38286 6264 38292 6276
rect 38344 6264 38350 6316
rect 18248 6208 20760 6236
rect 18141 6199 18199 6205
rect 18156 6168 18184 6199
rect 20898 6196 20904 6248
rect 20956 6236 20962 6248
rect 20993 6239 21051 6245
rect 20993 6236 21005 6239
rect 20956 6208 21005 6236
rect 20956 6196 20962 6208
rect 20993 6205 21005 6208
rect 21039 6205 21051 6239
rect 22922 6236 22928 6248
rect 20993 6199 21051 6205
rect 21376 6208 22928 6236
rect 21376 6168 21404 6208
rect 22922 6196 22928 6208
rect 22980 6196 22986 6248
rect 23109 6239 23167 6245
rect 23109 6205 23121 6239
rect 23155 6205 23167 6239
rect 23109 6199 23167 6205
rect 18156 6140 21404 6168
rect 21450 6128 21456 6180
rect 21508 6168 21514 6180
rect 22097 6171 22155 6177
rect 22097 6168 22109 6171
rect 21508 6140 22109 6168
rect 21508 6128 21514 6140
rect 22097 6137 22109 6140
rect 22143 6137 22155 6171
rect 23124 6168 23152 6199
rect 24946 6196 24952 6248
rect 25004 6236 25010 6248
rect 25225 6239 25283 6245
rect 25225 6236 25237 6239
rect 25004 6208 25237 6236
rect 25004 6196 25010 6208
rect 25225 6205 25237 6208
rect 25271 6205 25283 6239
rect 25225 6199 25283 6205
rect 28166 6196 28172 6248
rect 28224 6236 28230 6248
rect 28445 6239 28503 6245
rect 28445 6236 28457 6239
rect 28224 6208 28457 6236
rect 28224 6196 28230 6208
rect 28445 6205 28457 6208
rect 28491 6205 28503 6239
rect 30650 6236 30656 6248
rect 28445 6199 28503 6205
rect 28736 6208 30656 6236
rect 24670 6168 24676 6180
rect 23124 6140 24676 6168
rect 22097 6131 22155 6137
rect 24670 6128 24676 6140
rect 24728 6128 24734 6180
rect 27798 6168 27804 6180
rect 27759 6140 27804 6168
rect 27798 6128 27804 6140
rect 27856 6168 27862 6180
rect 28626 6168 28632 6180
rect 27856 6140 28632 6168
rect 27856 6128 27862 6140
rect 28626 6128 28632 6140
rect 28684 6128 28690 6180
rect 18598 6100 18604 6112
rect 9364 6072 18092 6100
rect 18559 6072 18604 6100
rect 9364 6060 9370 6072
rect 18598 6060 18604 6072
rect 18656 6060 18662 6112
rect 18690 6060 18696 6112
rect 18748 6100 18754 6112
rect 19153 6103 19211 6109
rect 19153 6100 19165 6103
rect 18748 6072 19165 6100
rect 18748 6060 18754 6072
rect 19153 6069 19165 6072
rect 19199 6069 19211 6103
rect 19153 6063 19211 6069
rect 21174 6060 21180 6112
rect 21232 6100 21238 6112
rect 21542 6100 21548 6112
rect 21232 6072 21548 6100
rect 21232 6060 21238 6072
rect 21542 6060 21548 6072
rect 21600 6060 21606 6112
rect 23014 6060 23020 6112
rect 23072 6100 23078 6112
rect 28736 6100 28764 6208
rect 30650 6196 30656 6208
rect 30708 6196 30714 6248
rect 30837 6239 30895 6245
rect 30837 6205 30849 6239
rect 30883 6205 30895 6239
rect 30837 6199 30895 6205
rect 30009 6171 30067 6177
rect 30009 6137 30021 6171
rect 30055 6168 30067 6171
rect 30852 6168 30880 6199
rect 30055 6140 30880 6168
rect 30055 6137 30067 6140
rect 30009 6131 30067 6137
rect 38102 6100 38108 6112
rect 23072 6072 28764 6100
rect 38063 6072 38108 6100
rect 23072 6060 23078 6072
rect 38102 6060 38108 6072
rect 38160 6060 38166 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 1578 5896 1584 5908
rect 1539 5868 1584 5896
rect 1578 5856 1584 5868
rect 1636 5856 1642 5908
rect 5721 5899 5779 5905
rect 5721 5865 5733 5899
rect 5767 5896 5779 5899
rect 6178 5896 6184 5908
rect 5767 5868 6184 5896
rect 5767 5865 5779 5868
rect 5721 5859 5779 5865
rect 6178 5856 6184 5868
rect 6236 5856 6242 5908
rect 12158 5856 12164 5908
rect 12216 5896 12222 5908
rect 13173 5899 13231 5905
rect 13173 5896 13185 5899
rect 12216 5868 13185 5896
rect 12216 5856 12222 5868
rect 13173 5865 13185 5868
rect 13219 5865 13231 5899
rect 13173 5859 13231 5865
rect 16022 5856 16028 5908
rect 16080 5896 16086 5908
rect 16380 5899 16438 5905
rect 16380 5896 16392 5899
rect 16080 5868 16392 5896
rect 16080 5856 16086 5868
rect 16380 5865 16392 5868
rect 16426 5896 16438 5899
rect 16426 5868 21772 5896
rect 16426 5865 16438 5868
rect 16380 5859 16438 5865
rect 9306 5828 9312 5840
rect 5368 5800 9312 5828
rect 1762 5692 1768 5704
rect 1723 5664 1768 5692
rect 1762 5652 1768 5664
rect 1820 5652 1826 5704
rect 3970 5692 3976 5704
rect 3931 5664 3976 5692
rect 3970 5652 3976 5664
rect 4028 5652 4034 5704
rect 5368 5678 5396 5800
rect 9306 5788 9312 5800
rect 9364 5788 9370 5840
rect 14200 5800 16252 5828
rect 8662 5720 8668 5772
rect 8720 5760 8726 5772
rect 14200 5760 14228 5800
rect 8720 5732 14228 5760
rect 16224 5760 16252 5800
rect 18598 5788 18604 5840
rect 18656 5828 18662 5840
rect 21450 5828 21456 5840
rect 18656 5800 21456 5828
rect 18656 5788 18662 5800
rect 21450 5788 21456 5800
rect 21508 5788 21514 5840
rect 21744 5828 21772 5868
rect 22094 5856 22100 5908
rect 22152 5896 22158 5908
rect 22152 5868 22197 5896
rect 22480 5868 23152 5896
rect 22152 5856 22158 5868
rect 22480 5828 22508 5868
rect 21744 5800 22508 5828
rect 20990 5760 20996 5772
rect 16224 5732 20996 5760
rect 8720 5720 8726 5732
rect 20990 5720 20996 5732
rect 21048 5720 21054 5772
rect 21634 5720 21640 5772
rect 21692 5760 21698 5772
rect 22741 5763 22799 5769
rect 22741 5760 22753 5763
rect 21692 5732 22753 5760
rect 21692 5720 21698 5732
rect 22741 5729 22753 5732
rect 22787 5729 22799 5763
rect 23124 5760 23152 5868
rect 23198 5856 23204 5908
rect 23256 5896 23262 5908
rect 25225 5899 25283 5905
rect 25225 5896 25237 5899
rect 23256 5868 25237 5896
rect 23256 5856 23262 5868
rect 25225 5865 25237 5868
rect 25271 5865 25283 5899
rect 25225 5859 25283 5865
rect 25866 5856 25872 5908
rect 25924 5896 25930 5908
rect 26053 5899 26111 5905
rect 26053 5896 26065 5899
rect 25924 5868 26065 5896
rect 25924 5856 25930 5868
rect 26053 5865 26065 5868
rect 26099 5865 26111 5899
rect 27614 5896 27620 5908
rect 27575 5868 27620 5896
rect 26053 5859 26111 5865
rect 27614 5856 27620 5868
rect 27672 5856 27678 5908
rect 28810 5896 28816 5908
rect 28771 5868 28816 5896
rect 28810 5856 28816 5868
rect 28868 5856 28874 5908
rect 30006 5896 30012 5908
rect 29967 5868 30012 5896
rect 30006 5856 30012 5868
rect 30064 5856 30070 5908
rect 30650 5856 30656 5908
rect 30708 5896 30714 5908
rect 30929 5899 30987 5905
rect 30929 5896 30941 5899
rect 30708 5868 30941 5896
rect 30708 5856 30714 5868
rect 30929 5865 30941 5868
rect 30975 5865 30987 5899
rect 30929 5859 30987 5865
rect 23290 5788 23296 5840
rect 23348 5828 23354 5840
rect 24673 5831 24731 5837
rect 24673 5828 24685 5831
rect 23348 5800 24685 5828
rect 23348 5788 23354 5800
rect 24673 5797 24685 5800
rect 24719 5797 24731 5831
rect 24673 5791 24731 5797
rect 27982 5760 27988 5772
rect 23124 5732 27988 5760
rect 22741 5723 22799 5729
rect 9214 5652 9220 5704
rect 9272 5692 9278 5704
rect 11146 5692 11152 5704
rect 9272 5664 11152 5692
rect 9272 5652 9278 5664
rect 11146 5652 11152 5664
rect 11204 5692 11210 5704
rect 11425 5695 11483 5701
rect 11425 5692 11437 5695
rect 11204 5664 11437 5692
rect 11204 5652 11210 5664
rect 11425 5661 11437 5664
rect 11471 5661 11483 5695
rect 11425 5655 11483 5661
rect 16117 5695 16175 5701
rect 16117 5661 16129 5695
rect 16163 5661 16175 5695
rect 16117 5655 16175 5661
rect 4249 5627 4307 5633
rect 4249 5593 4261 5627
rect 4295 5593 4307 5627
rect 11440 5624 11468 5655
rect 11606 5624 11612 5636
rect 11440 5596 11612 5624
rect 4249 5587 4307 5593
rect 4264 5556 4292 5587
rect 11606 5584 11612 5596
rect 11664 5584 11670 5636
rect 11701 5627 11759 5633
rect 11701 5593 11713 5627
rect 11747 5624 11759 5627
rect 11974 5624 11980 5636
rect 11747 5596 11980 5624
rect 11747 5593 11759 5596
rect 11701 5587 11759 5593
rect 11974 5584 11980 5596
rect 12032 5584 12038 5636
rect 13630 5624 13636 5636
rect 12926 5596 13636 5624
rect 13630 5584 13636 5596
rect 13688 5584 13694 5636
rect 14274 5584 14280 5636
rect 14332 5624 14338 5636
rect 16132 5624 16160 5655
rect 14332 5596 16423 5624
rect 14332 5584 14338 5596
rect 16298 5556 16304 5568
rect 4264 5528 16304 5556
rect 16298 5516 16304 5528
rect 16356 5516 16362 5568
rect 16395 5556 16423 5596
rect 17218 5556 17224 5568
rect 16395 5528 17224 5556
rect 17218 5516 17224 5528
rect 17276 5516 17282 5568
rect 17512 5556 17540 5678
rect 21726 5652 21732 5704
rect 21784 5692 21790 5704
rect 22005 5695 22063 5701
rect 22005 5692 22017 5695
rect 21784 5664 22017 5692
rect 21784 5652 21790 5664
rect 22005 5661 22017 5664
rect 22051 5661 22063 5695
rect 22005 5655 22063 5661
rect 22370 5652 22376 5704
rect 22428 5692 22434 5704
rect 22646 5692 22652 5704
rect 22428 5664 22652 5692
rect 22428 5652 22434 5664
rect 22646 5652 22652 5664
rect 22704 5652 22710 5704
rect 23293 5695 23351 5701
rect 23293 5661 23305 5695
rect 23339 5692 23351 5695
rect 23474 5692 23480 5704
rect 23339 5664 23480 5692
rect 23339 5661 23351 5664
rect 23293 5655 23351 5661
rect 23474 5652 23480 5664
rect 23532 5652 23538 5704
rect 23842 5652 23848 5704
rect 23900 5692 23906 5704
rect 24581 5695 24639 5701
rect 24581 5692 24593 5695
rect 23900 5664 24593 5692
rect 23900 5652 23906 5664
rect 24581 5661 24593 5664
rect 24627 5661 24639 5695
rect 25406 5692 25412 5704
rect 25367 5664 25412 5692
rect 24581 5655 24639 5661
rect 25406 5652 25412 5664
rect 25464 5652 25470 5704
rect 25961 5695 26019 5701
rect 25961 5661 25973 5695
rect 26007 5692 26019 5695
rect 27430 5692 27436 5704
rect 26007 5664 27436 5692
rect 26007 5661 26019 5664
rect 25961 5655 26019 5661
rect 27430 5652 27436 5664
rect 27488 5652 27494 5704
rect 27540 5701 27568 5732
rect 27982 5720 27988 5732
rect 28040 5720 28046 5772
rect 28166 5760 28172 5772
rect 28127 5732 28172 5760
rect 28166 5720 28172 5732
rect 28224 5720 28230 5772
rect 27525 5695 27583 5701
rect 27525 5661 27537 5695
rect 27571 5661 27583 5695
rect 28994 5692 29000 5704
rect 28955 5664 29000 5692
rect 27525 5655 27583 5661
rect 28994 5652 29000 5664
rect 29052 5652 29058 5704
rect 30190 5692 30196 5704
rect 30151 5664 30196 5692
rect 30190 5652 30196 5664
rect 30248 5652 30254 5704
rect 30837 5695 30895 5701
rect 30837 5661 30849 5695
rect 30883 5692 30895 5695
rect 38102 5692 38108 5704
rect 30883 5664 38108 5692
rect 30883 5661 30895 5664
rect 30837 5655 30895 5661
rect 38102 5652 38108 5664
rect 38160 5652 38166 5704
rect 18138 5584 18144 5636
rect 18196 5624 18202 5636
rect 20898 5624 20904 5636
rect 18196 5596 18241 5624
rect 20859 5596 20904 5624
rect 18196 5584 18202 5596
rect 20898 5584 20904 5596
rect 20956 5584 20962 5636
rect 20993 5627 21051 5633
rect 20993 5593 21005 5627
rect 21039 5624 21051 5627
rect 21358 5624 21364 5636
rect 21039 5596 21364 5624
rect 21039 5593 21051 5596
rect 20993 5587 21051 5593
rect 21358 5584 21364 5596
rect 21416 5584 21422 5636
rect 21542 5624 21548 5636
rect 21503 5596 21548 5624
rect 21542 5584 21548 5596
rect 21600 5584 21606 5636
rect 23385 5627 23443 5633
rect 23385 5624 23397 5627
rect 22664 5596 23397 5624
rect 20162 5556 20168 5568
rect 17512 5528 20168 5556
rect 20162 5516 20168 5528
rect 20220 5516 20226 5568
rect 20622 5516 20628 5568
rect 20680 5556 20686 5568
rect 22664 5556 22692 5596
rect 23385 5593 23397 5596
rect 23431 5593 23443 5627
rect 23385 5587 23443 5593
rect 20680 5528 22692 5556
rect 20680 5516 20686 5528
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 7006 5352 7012 5364
rect 2332 5324 7012 5352
rect 1486 5176 1492 5228
rect 1544 5216 1550 5228
rect 2332 5225 2360 5324
rect 7006 5312 7012 5324
rect 7064 5312 7070 5364
rect 8772 5324 13952 5352
rect 3970 5284 3976 5296
rect 3712 5256 3976 5284
rect 3712 5225 3740 5256
rect 3970 5244 3976 5256
rect 4028 5244 4034 5296
rect 8772 5284 8800 5324
rect 11146 5284 11152 5296
rect 5198 5256 8800 5284
rect 10718 5256 11152 5284
rect 11146 5244 11152 5256
rect 11204 5244 11210 5296
rect 1581 5219 1639 5225
rect 1581 5216 1593 5219
rect 1544 5188 1593 5216
rect 1544 5176 1550 5188
rect 1581 5185 1593 5188
rect 1627 5185 1639 5219
rect 1581 5179 1639 5185
rect 2317 5219 2375 5225
rect 2317 5185 2329 5219
rect 2363 5185 2375 5219
rect 2317 5179 2375 5185
rect 3697 5219 3755 5225
rect 3697 5185 3709 5219
rect 3743 5185 3755 5219
rect 9214 5216 9220 5228
rect 9175 5188 9220 5216
rect 3697 5179 3755 5185
rect 9214 5176 9220 5188
rect 9272 5176 9278 5228
rect 3973 5151 4031 5157
rect 3973 5117 3985 5151
rect 4019 5148 4031 5151
rect 9493 5151 9551 5157
rect 9493 5148 9505 5151
rect 4019 5120 6224 5148
rect 4019 5117 4031 5120
rect 3973 5111 4031 5117
rect 5442 5080 5448 5092
rect 5403 5052 5448 5080
rect 5442 5040 5448 5052
rect 5500 5040 5506 5092
rect 1762 5012 1768 5024
rect 1723 4984 1768 5012
rect 1762 4972 1768 4984
rect 1820 4972 1826 5024
rect 2409 5015 2467 5021
rect 2409 4981 2421 5015
rect 2455 5012 2467 5015
rect 2498 5012 2504 5024
rect 2455 4984 2504 5012
rect 2455 4981 2467 4984
rect 2409 4975 2467 4981
rect 2498 4972 2504 4984
rect 2556 4972 2562 5024
rect 6196 5012 6224 5120
rect 8956 5120 9505 5148
rect 6270 5040 6276 5092
rect 6328 5080 6334 5092
rect 8956 5080 8984 5120
rect 9493 5117 9505 5120
rect 9539 5117 9551 5151
rect 9493 5111 9551 5117
rect 10778 5108 10784 5160
rect 10836 5148 10842 5160
rect 10965 5151 11023 5157
rect 10965 5148 10977 5151
rect 10836 5120 10977 5148
rect 10836 5108 10842 5120
rect 10965 5117 10977 5120
rect 11011 5117 11023 5151
rect 13924 5148 13952 5324
rect 13998 5312 14004 5364
rect 14056 5352 14062 5364
rect 14056 5324 20760 5352
rect 14056 5312 14062 5324
rect 14182 5284 14188 5296
rect 14016 5256 14188 5284
rect 14016 5225 14044 5256
rect 14182 5244 14188 5256
rect 14240 5244 14246 5296
rect 14292 5293 14320 5324
rect 14277 5287 14335 5293
rect 14277 5253 14289 5287
rect 14323 5253 14335 5287
rect 18506 5284 18512 5296
rect 15502 5256 18512 5284
rect 14277 5247 14335 5253
rect 18506 5244 18512 5256
rect 18564 5244 18570 5296
rect 20622 5284 20628 5296
rect 19458 5256 20628 5284
rect 20622 5244 20628 5256
rect 20680 5244 20686 5296
rect 13990 5219 14048 5225
rect 13990 5185 14002 5219
rect 14036 5185 14048 5219
rect 17126 5216 17132 5228
rect 17087 5188 17132 5216
rect 13990 5179 14048 5185
rect 17126 5176 17132 5188
rect 17184 5176 17190 5228
rect 17034 5148 17040 5160
rect 13924 5120 17040 5148
rect 10965 5111 11023 5117
rect 17034 5108 17040 5120
rect 17092 5108 17098 5160
rect 17218 5108 17224 5160
rect 17276 5148 17282 5160
rect 17954 5148 17960 5160
rect 17276 5120 17960 5148
rect 17276 5108 17282 5120
rect 17954 5108 17960 5120
rect 18012 5108 18018 5160
rect 18233 5151 18291 5157
rect 18233 5117 18245 5151
rect 18279 5148 18291 5151
rect 18322 5148 18328 5160
rect 18279 5120 18328 5148
rect 18279 5117 18291 5120
rect 18233 5111 18291 5117
rect 18322 5108 18328 5120
rect 18380 5108 18386 5160
rect 18598 5108 18604 5160
rect 18656 5148 18662 5160
rect 20622 5148 20628 5160
rect 18656 5120 20628 5148
rect 18656 5108 18662 5120
rect 20622 5108 20628 5120
rect 20680 5108 20686 5160
rect 20732 5148 20760 5324
rect 21266 5312 21272 5364
rect 21324 5352 21330 5364
rect 21361 5355 21419 5361
rect 21361 5352 21373 5355
rect 21324 5324 21373 5352
rect 21324 5312 21330 5324
rect 21361 5321 21373 5324
rect 21407 5321 21419 5355
rect 21361 5315 21419 5321
rect 22922 5312 22928 5364
rect 22980 5352 22986 5364
rect 23385 5355 23443 5361
rect 23385 5352 23397 5355
rect 22980 5324 23397 5352
rect 22980 5312 22986 5324
rect 23385 5321 23397 5324
rect 23431 5321 23443 5355
rect 23385 5315 23443 5321
rect 23474 5312 23480 5364
rect 23532 5352 23538 5364
rect 24578 5352 24584 5364
rect 23532 5324 24584 5352
rect 23532 5312 23538 5324
rect 24578 5312 24584 5324
rect 24636 5312 24642 5364
rect 25406 5312 25412 5364
rect 25464 5352 25470 5364
rect 25869 5355 25927 5361
rect 25869 5352 25881 5355
rect 25464 5324 25881 5352
rect 25464 5312 25470 5324
rect 25869 5321 25881 5324
rect 25915 5321 25927 5355
rect 25869 5315 25927 5321
rect 27157 5355 27215 5361
rect 27157 5321 27169 5355
rect 27203 5352 27215 5355
rect 28994 5352 29000 5364
rect 27203 5324 29000 5352
rect 27203 5321 27215 5324
rect 27157 5315 27215 5321
rect 28994 5312 29000 5324
rect 29052 5312 29058 5364
rect 29086 5312 29092 5364
rect 29144 5352 29150 5364
rect 29825 5355 29883 5361
rect 29825 5352 29837 5355
rect 29144 5324 29837 5352
rect 29144 5312 29150 5324
rect 29825 5321 29837 5324
rect 29871 5321 29883 5355
rect 29825 5315 29883 5321
rect 22370 5284 22376 5296
rect 21284 5256 22376 5284
rect 21284 5225 21312 5256
rect 22370 5244 22376 5256
rect 22428 5244 22434 5296
rect 22646 5244 22652 5296
rect 22704 5284 22710 5296
rect 22704 5256 26096 5284
rect 22704 5244 22710 5256
rect 21269 5219 21327 5225
rect 21269 5185 21281 5219
rect 21315 5185 21327 5219
rect 21269 5179 21327 5185
rect 22097 5219 22155 5225
rect 22097 5185 22109 5219
rect 22143 5216 22155 5219
rect 22462 5216 22468 5228
rect 22143 5188 22468 5216
rect 22143 5185 22155 5188
rect 22097 5179 22155 5185
rect 22462 5176 22468 5188
rect 22520 5176 22526 5228
rect 23293 5219 23351 5225
rect 23293 5185 23305 5219
rect 23339 5185 23351 5219
rect 23293 5179 23351 5185
rect 23937 5219 23995 5225
rect 23937 5185 23949 5219
rect 23983 5216 23995 5219
rect 24026 5216 24032 5228
rect 23983 5188 24032 5216
rect 23983 5185 23995 5188
rect 23937 5179 23995 5185
rect 23308 5148 23336 5179
rect 24026 5176 24032 5188
rect 24084 5176 24090 5228
rect 24578 5216 24584 5228
rect 24539 5188 24584 5216
rect 24578 5176 24584 5188
rect 24636 5176 24642 5228
rect 24670 5176 24676 5228
rect 24728 5216 24734 5228
rect 25866 5216 25872 5228
rect 24728 5188 25872 5216
rect 24728 5176 24734 5188
rect 25866 5176 25872 5188
rect 25924 5176 25930 5228
rect 26068 5225 26096 5256
rect 26510 5244 26516 5296
rect 26568 5284 26574 5296
rect 36722 5284 36728 5296
rect 26568 5256 28488 5284
rect 26568 5244 26574 5256
rect 26053 5219 26111 5225
rect 26053 5185 26065 5219
rect 26099 5185 26111 5219
rect 26053 5179 26111 5185
rect 27341 5219 27399 5225
rect 27341 5185 27353 5219
rect 27387 5185 27399 5219
rect 27982 5216 27988 5228
rect 27943 5188 27988 5216
rect 27341 5179 27399 5185
rect 20732 5120 23336 5148
rect 6328 5052 8984 5080
rect 6328 5040 6334 5052
rect 19334 5040 19340 5092
rect 19392 5080 19398 5092
rect 22189 5083 22247 5089
rect 22189 5080 22201 5083
rect 19392 5052 22201 5080
rect 19392 5040 19398 5052
rect 22189 5049 22201 5052
rect 22235 5049 22247 5083
rect 23308 5080 23336 5120
rect 23382 5108 23388 5160
rect 23440 5148 23446 5160
rect 25225 5151 25283 5157
rect 25225 5148 25237 5151
rect 23440 5120 25237 5148
rect 23440 5108 23446 5120
rect 25225 5117 25237 5120
rect 25271 5117 25283 5151
rect 25225 5111 25283 5117
rect 26510 5080 26516 5092
rect 23308 5052 26516 5080
rect 22189 5043 22247 5049
rect 26510 5040 26516 5052
rect 26568 5040 26574 5092
rect 10686 5012 10692 5024
rect 6196 4984 10692 5012
rect 10686 4972 10692 4984
rect 10744 4972 10750 5024
rect 11054 4972 11060 5024
rect 11112 5012 11118 5024
rect 13906 5012 13912 5024
rect 11112 4984 13912 5012
rect 11112 4972 11118 4984
rect 13906 4972 13912 4984
rect 13964 4972 13970 5024
rect 15746 5012 15752 5024
rect 15707 4984 15752 5012
rect 15746 4972 15752 4984
rect 15804 4972 15810 5024
rect 16945 5015 17003 5021
rect 16945 4981 16957 5015
rect 16991 5012 17003 5015
rect 19426 5012 19432 5024
rect 16991 4984 19432 5012
rect 16991 4981 17003 4984
rect 16945 4975 17003 4981
rect 19426 4972 19432 4984
rect 19484 4972 19490 5024
rect 19518 4972 19524 5024
rect 19576 5012 19582 5024
rect 19705 5015 19763 5021
rect 19705 5012 19717 5015
rect 19576 4984 19717 5012
rect 19576 4972 19582 4984
rect 19705 4981 19717 4984
rect 19751 4981 19763 5015
rect 19705 4975 19763 4981
rect 20070 4972 20076 5024
rect 20128 5012 20134 5024
rect 21726 5012 21732 5024
rect 20128 4984 21732 5012
rect 20128 4972 20134 4984
rect 21726 4972 21732 4984
rect 21784 4972 21790 5024
rect 23934 4972 23940 5024
rect 23992 5012 23998 5024
rect 24029 5015 24087 5021
rect 24029 5012 24041 5015
rect 23992 4984 24041 5012
rect 23992 4972 23998 4984
rect 24029 4981 24041 4984
rect 24075 4981 24087 5015
rect 24670 5012 24676 5024
rect 24631 4984 24676 5012
rect 24029 4975 24087 4981
rect 24670 4972 24676 4984
rect 24728 4972 24734 5024
rect 24762 4972 24768 5024
rect 24820 5012 24826 5024
rect 27356 5012 27384 5179
rect 27982 5176 27988 5188
rect 28040 5176 28046 5228
rect 28460 5225 28488 5256
rect 29748 5256 36728 5284
rect 29748 5225 29776 5256
rect 36722 5244 36728 5256
rect 36780 5244 36786 5296
rect 28445 5219 28503 5225
rect 28445 5185 28457 5219
rect 28491 5185 28503 5219
rect 28445 5179 28503 5185
rect 29733 5219 29791 5225
rect 29733 5185 29745 5219
rect 29779 5185 29791 5219
rect 29733 5179 29791 5185
rect 30561 5219 30619 5225
rect 30561 5185 30573 5219
rect 30607 5185 30619 5219
rect 31202 5216 31208 5228
rect 31163 5188 31208 5216
rect 30561 5179 30619 5185
rect 28537 5151 28595 5157
rect 28537 5117 28549 5151
rect 28583 5148 28595 5151
rect 30576 5148 30604 5179
rect 31202 5176 31208 5188
rect 31260 5176 31266 5228
rect 28583 5120 30604 5148
rect 28583 5117 28595 5120
rect 28537 5111 28595 5117
rect 30377 5083 30435 5089
rect 30377 5049 30389 5083
rect 30423 5080 30435 5083
rect 33318 5080 33324 5092
rect 30423 5052 33324 5080
rect 30423 5049 30435 5052
rect 30377 5043 30435 5049
rect 33318 5040 33324 5052
rect 33376 5040 33382 5092
rect 24820 4984 27384 5012
rect 27801 5015 27859 5021
rect 24820 4972 24826 4984
rect 27801 4981 27813 5015
rect 27847 5012 27859 5015
rect 28074 5012 28080 5024
rect 27847 4984 28080 5012
rect 27847 4981 27859 4984
rect 27801 4975 27859 4981
rect 28074 4972 28080 4984
rect 28132 4972 28138 5024
rect 31021 5015 31079 5021
rect 31021 4981 31033 5015
rect 31067 5012 31079 5015
rect 32950 5012 32956 5024
rect 31067 4984 32956 5012
rect 31067 4981 31079 4984
rect 31021 4975 31079 4981
rect 32950 4972 32956 4984
rect 33008 4972 33014 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 11330 4808 11336 4820
rect 6012 4780 11336 4808
rect 4249 4675 4307 4681
rect 4249 4641 4261 4675
rect 4295 4672 4307 4675
rect 5718 4672 5724 4684
rect 4295 4644 5724 4672
rect 4295 4641 4307 4644
rect 4249 4635 4307 4641
rect 5718 4632 5724 4644
rect 5776 4632 5782 4684
rect 6012 4681 6040 4780
rect 11330 4768 11336 4780
rect 11388 4768 11394 4820
rect 11974 4768 11980 4820
rect 12032 4808 12038 4820
rect 12250 4808 12256 4820
rect 12032 4780 12256 4808
rect 12032 4768 12038 4780
rect 12250 4768 12256 4780
rect 12308 4768 12314 4820
rect 12342 4768 12348 4820
rect 12400 4808 12406 4820
rect 13998 4808 14004 4820
rect 12400 4780 14004 4808
rect 12400 4768 12406 4780
rect 13998 4768 14004 4780
rect 14056 4768 14062 4820
rect 16945 4811 17003 4817
rect 16945 4808 16957 4811
rect 14384 4780 16957 4808
rect 14384 4740 14412 4780
rect 16945 4777 16957 4780
rect 16991 4777 17003 4811
rect 16945 4771 17003 4777
rect 17034 4768 17040 4820
rect 17092 4808 17098 4820
rect 24670 4808 24676 4820
rect 17092 4780 24676 4808
rect 17092 4768 17098 4780
rect 24670 4768 24676 4780
rect 24728 4768 24734 4820
rect 26329 4811 26387 4817
rect 26329 4777 26341 4811
rect 26375 4808 26387 4811
rect 27982 4808 27988 4820
rect 26375 4780 27988 4808
rect 26375 4777 26387 4780
rect 26329 4771 26387 4777
rect 27982 4768 27988 4780
rect 28040 4768 28046 4820
rect 16022 4740 16028 4752
rect 11808 4712 14412 4740
rect 15983 4712 16028 4740
rect 5997 4675 6055 4681
rect 5997 4641 6009 4675
rect 6043 4641 6055 4675
rect 5997 4635 6055 4641
rect 9674 4632 9680 4684
rect 9732 4672 9738 4684
rect 11808 4672 11836 4712
rect 16022 4700 16028 4712
rect 16080 4700 16086 4752
rect 16850 4700 16856 4752
rect 16908 4740 16914 4752
rect 18138 4740 18144 4752
rect 16908 4712 18144 4740
rect 16908 4700 16914 4712
rect 18138 4700 18144 4712
rect 18196 4700 18202 4752
rect 18230 4700 18236 4752
rect 18288 4740 18294 4752
rect 18288 4712 18333 4740
rect 18288 4700 18294 4712
rect 18414 4700 18420 4752
rect 18472 4740 18478 4752
rect 19978 4740 19984 4752
rect 18472 4712 19984 4740
rect 18472 4700 18478 4712
rect 19978 4700 19984 4712
rect 20036 4700 20042 4752
rect 20622 4700 20628 4752
rect 20680 4740 20686 4752
rect 21453 4743 21511 4749
rect 21453 4740 21465 4743
rect 20680 4712 21465 4740
rect 20680 4700 20686 4712
rect 21453 4709 21465 4712
rect 21499 4709 21511 4743
rect 24026 4740 24032 4752
rect 23939 4712 24032 4740
rect 21453 4703 21511 4709
rect 24026 4700 24032 4712
rect 24084 4740 24090 4752
rect 25593 4743 25651 4749
rect 25593 4740 25605 4743
rect 24084 4712 25605 4740
rect 24084 4700 24090 4712
rect 25593 4709 25605 4712
rect 25639 4709 25651 4743
rect 25593 4703 25651 4709
rect 27341 4743 27399 4749
rect 27341 4709 27353 4743
rect 27387 4740 27399 4743
rect 27706 4740 27712 4752
rect 27387 4712 27712 4740
rect 27387 4709 27399 4712
rect 27341 4703 27399 4709
rect 27706 4700 27712 4712
rect 27764 4700 27770 4752
rect 28261 4743 28319 4749
rect 28261 4740 28273 4743
rect 27816 4712 28273 4740
rect 19334 4672 19340 4684
rect 9732 4644 11836 4672
rect 11900 4644 19340 4672
rect 9732 4632 9738 4644
rect 3970 4604 3976 4616
rect 3931 4576 3976 4604
rect 3970 4564 3976 4576
rect 4028 4564 4034 4616
rect 10502 4604 10508 4616
rect 10463 4576 10508 4604
rect 10502 4564 10508 4576
rect 10560 4564 10566 4616
rect 11900 4590 11928 4644
rect 19334 4632 19340 4644
rect 19392 4632 19398 4684
rect 22462 4672 22468 4684
rect 21376 4644 22468 4672
rect 14274 4604 14280 4616
rect 14235 4576 14280 4604
rect 14274 4564 14280 4576
rect 14332 4564 14338 4616
rect 16853 4607 16911 4613
rect 16853 4573 16865 4607
rect 16899 4604 16911 4607
rect 17034 4604 17040 4616
rect 16899 4576 17040 4604
rect 16899 4573 16911 4576
rect 16853 4567 16911 4573
rect 17034 4564 17040 4576
rect 17092 4564 17098 4616
rect 17497 4607 17555 4613
rect 17497 4573 17509 4607
rect 17543 4604 17555 4607
rect 18046 4604 18052 4616
rect 17543 4576 18052 4604
rect 17543 4573 17555 4576
rect 17497 4567 17555 4573
rect 18046 4564 18052 4576
rect 18104 4564 18110 4616
rect 18141 4607 18199 4613
rect 18141 4573 18153 4607
rect 18187 4604 18199 4607
rect 19242 4604 19248 4616
rect 18187 4576 19248 4604
rect 18187 4573 18199 4576
rect 18141 4567 18199 4573
rect 19242 4564 19248 4576
rect 19300 4564 19306 4616
rect 20070 4564 20076 4616
rect 20128 4604 20134 4616
rect 21376 4613 21404 4644
rect 22462 4632 22468 4644
rect 22520 4632 22526 4684
rect 23382 4672 23388 4684
rect 23343 4644 23388 4672
rect 23382 4632 23388 4644
rect 23440 4632 23446 4684
rect 24670 4632 24676 4684
rect 24728 4672 24734 4684
rect 25409 4675 25467 4681
rect 25409 4672 25421 4675
rect 24728 4644 25421 4672
rect 24728 4632 24734 4644
rect 25409 4641 25421 4644
rect 25455 4641 25467 4675
rect 27816 4672 27844 4712
rect 28261 4709 28273 4712
rect 28307 4709 28319 4743
rect 28261 4703 28319 4709
rect 28074 4672 28080 4684
rect 25409 4635 25467 4641
rect 25516 4644 27844 4672
rect 28035 4644 28080 4672
rect 20441 4607 20499 4613
rect 20441 4604 20453 4607
rect 20128 4576 20453 4604
rect 20128 4564 20134 4576
rect 20441 4573 20453 4576
rect 20487 4573 20499 4607
rect 20441 4567 20499 4573
rect 21361 4607 21419 4613
rect 21361 4573 21373 4607
rect 21407 4573 21419 4607
rect 21361 4567 21419 4573
rect 22005 4607 22063 4613
rect 22005 4573 22017 4607
rect 22051 4604 22063 4607
rect 22370 4604 22376 4616
rect 22051 4576 22376 4604
rect 22051 4573 22063 4576
rect 22005 4567 22063 4573
rect 22370 4564 22376 4576
rect 22428 4564 22434 4616
rect 23569 4607 23627 4613
rect 23569 4573 23581 4607
rect 23615 4573 23627 4607
rect 23569 4567 23627 4573
rect 24581 4607 24639 4613
rect 24581 4573 24593 4607
rect 24627 4604 24639 4607
rect 24762 4604 24768 4616
rect 24627 4576 24768 4604
rect 24627 4573 24639 4576
rect 24581 4567 24639 4573
rect 5902 4536 5908 4548
rect 5474 4508 5908 4536
rect 5902 4496 5908 4508
rect 5960 4496 5966 4548
rect 10781 4539 10839 4545
rect 10781 4505 10793 4539
rect 10827 4536 10839 4539
rect 11054 4536 11060 4548
rect 10827 4508 11060 4536
rect 10827 4505 10839 4508
rect 10781 4499 10839 4505
rect 11054 4496 11060 4508
rect 11112 4496 11118 4548
rect 12342 4536 12348 4548
rect 12176 4508 12348 4536
rect 7282 4428 7288 4480
rect 7340 4468 7346 4480
rect 12176 4468 12204 4508
rect 12342 4496 12348 4508
rect 12400 4496 12406 4548
rect 14458 4496 14464 4548
rect 14516 4536 14522 4548
rect 14553 4539 14611 4545
rect 14553 4536 14565 4539
rect 14516 4508 14565 4536
rect 14516 4496 14522 4508
rect 14553 4505 14565 4508
rect 14599 4505 14611 4539
rect 20533 4539 20591 4545
rect 20533 4536 20545 4539
rect 15778 4508 20545 4536
rect 14553 4499 14611 4505
rect 20533 4505 20545 4508
rect 20579 4505 20591 4539
rect 23584 4536 23612 4567
rect 24762 4564 24768 4576
rect 24820 4564 24826 4616
rect 25222 4604 25228 4616
rect 25183 4576 25228 4604
rect 25222 4564 25228 4576
rect 25280 4604 25286 4616
rect 25516 4604 25544 4644
rect 28074 4632 28080 4644
rect 28132 4632 28138 4684
rect 26510 4604 26516 4616
rect 25280 4576 25544 4604
rect 26471 4576 26516 4604
rect 25280 4564 25286 4576
rect 26510 4564 26516 4576
rect 26568 4564 26574 4616
rect 27249 4607 27307 4613
rect 27249 4573 27261 4607
rect 27295 4573 27307 4607
rect 27890 4604 27896 4616
rect 27851 4576 27896 4604
rect 27249 4567 27307 4573
rect 24673 4539 24731 4545
rect 23584 4508 24624 4536
rect 20533 4499 20591 4505
rect 7340 4440 12204 4468
rect 7340 4428 7346 4440
rect 12250 4428 12256 4480
rect 12308 4468 12314 4480
rect 17218 4468 17224 4480
rect 12308 4440 17224 4468
rect 12308 4428 12314 4440
rect 17218 4428 17224 4440
rect 17276 4428 17282 4480
rect 17586 4468 17592 4480
rect 17547 4440 17592 4468
rect 17586 4428 17592 4440
rect 17644 4428 17650 4480
rect 17678 4428 17684 4480
rect 17736 4468 17742 4480
rect 22097 4471 22155 4477
rect 22097 4468 22109 4471
rect 17736 4440 22109 4468
rect 17736 4428 17742 4440
rect 22097 4437 22109 4440
rect 22143 4437 22155 4471
rect 24596 4468 24624 4508
rect 24673 4505 24685 4539
rect 24719 4536 24731 4539
rect 25314 4536 25320 4548
rect 24719 4508 25320 4536
rect 24719 4505 24731 4508
rect 24673 4499 24731 4505
rect 25314 4496 25320 4508
rect 25372 4496 25378 4548
rect 27264 4536 27292 4567
rect 27890 4564 27896 4576
rect 27948 4564 27954 4616
rect 28997 4607 29055 4613
rect 28997 4573 29009 4607
rect 29043 4604 29055 4607
rect 32858 4604 32864 4616
rect 29043 4576 32864 4604
rect 29043 4573 29055 4576
rect 28997 4567 29055 4573
rect 32858 4564 32864 4576
rect 32916 4564 32922 4616
rect 34422 4564 34428 4616
rect 34480 4604 34486 4616
rect 38013 4607 38071 4613
rect 38013 4604 38025 4607
rect 34480 4576 38025 4604
rect 34480 4564 34486 4576
rect 38013 4573 38025 4576
rect 38059 4573 38071 4607
rect 38013 4567 38071 4573
rect 29730 4536 29736 4548
rect 27264 4508 29736 4536
rect 29730 4496 29736 4508
rect 29788 4496 29794 4548
rect 25774 4468 25780 4480
rect 24596 4440 25780 4468
rect 22097 4431 22155 4437
rect 25774 4428 25780 4440
rect 25832 4428 25838 4480
rect 25866 4428 25872 4480
rect 25924 4468 25930 4480
rect 29089 4471 29147 4477
rect 29089 4468 29101 4471
rect 25924 4440 29101 4468
rect 25924 4428 25930 4440
rect 29089 4437 29101 4440
rect 29135 4437 29147 4471
rect 38194 4468 38200 4480
rect 38155 4440 38200 4468
rect 29089 4431 29147 4437
rect 38194 4428 38200 4440
rect 38252 4428 38258 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 5902 4224 5908 4276
rect 5960 4264 5966 4276
rect 13906 4264 13912 4276
rect 5960 4236 13912 4264
rect 5960 4224 5966 4236
rect 13906 4224 13912 4236
rect 13964 4224 13970 4276
rect 13998 4224 14004 4276
rect 14056 4264 14062 4276
rect 16850 4264 16856 4276
rect 14056 4236 16856 4264
rect 14056 4224 14062 4236
rect 16850 4224 16856 4236
rect 16908 4224 16914 4276
rect 16945 4267 17003 4273
rect 16945 4233 16957 4267
rect 16991 4264 17003 4267
rect 17126 4264 17132 4276
rect 16991 4236 17132 4264
rect 16991 4233 17003 4236
rect 16945 4227 17003 4233
rect 17126 4224 17132 4236
rect 17184 4224 17190 4276
rect 17218 4224 17224 4276
rect 17276 4264 17282 4276
rect 17276 4236 19380 4264
rect 17276 4224 17282 4236
rect 17586 4196 17592 4208
rect 14214 4168 17592 4196
rect 17586 4156 17592 4168
rect 17644 4156 17650 4208
rect 17954 4196 17960 4208
rect 17788 4168 17960 4196
rect 1765 4131 1823 4137
rect 1765 4097 1777 4131
rect 1811 4128 1823 4131
rect 2774 4128 2780 4140
rect 1811 4100 2780 4128
rect 1811 4097 1823 4100
rect 1765 4091 1823 4097
rect 2774 4088 2780 4100
rect 2832 4088 2838 4140
rect 5810 4088 5816 4140
rect 5868 4128 5874 4140
rect 7282 4128 7288 4140
rect 5868 4100 7288 4128
rect 5868 4088 5874 4100
rect 7282 4088 7288 4100
rect 7340 4088 7346 4140
rect 7374 4088 7380 4140
rect 7432 4128 7438 4140
rect 8297 4131 8355 4137
rect 8297 4128 8309 4131
rect 7432 4100 8309 4128
rect 7432 4088 7438 4100
rect 8297 4097 8309 4100
rect 8343 4097 8355 4131
rect 8297 4091 8355 4097
rect 8386 4088 8392 4140
rect 8444 4128 8450 4140
rect 16853 4131 16911 4137
rect 8444 4100 8489 4128
rect 8444 4088 8450 4100
rect 16853 4097 16865 4131
rect 16899 4128 16911 4131
rect 17678 4128 17684 4140
rect 16899 4100 17684 4128
rect 16899 4097 16911 4100
rect 16853 4091 16911 4097
rect 17678 4088 17684 4100
rect 17736 4088 17742 4140
rect 17788 4137 17816 4168
rect 17954 4156 17960 4168
rect 18012 4196 18018 4208
rect 18322 4196 18328 4208
rect 18012 4168 18328 4196
rect 18012 4156 18018 4168
rect 18322 4156 18328 4168
rect 18380 4156 18386 4208
rect 18506 4156 18512 4208
rect 18564 4156 18570 4208
rect 19352 4196 19380 4236
rect 19978 4224 19984 4276
rect 20036 4264 20042 4276
rect 24762 4264 24768 4276
rect 20036 4236 24768 4264
rect 20036 4224 20042 4236
rect 24762 4224 24768 4236
rect 24820 4224 24826 4276
rect 25774 4264 25780 4276
rect 25735 4236 25780 4264
rect 25774 4224 25780 4236
rect 25832 4224 25838 4276
rect 27890 4224 27896 4276
rect 27948 4264 27954 4276
rect 28169 4267 28227 4273
rect 28169 4264 28181 4267
rect 27948 4236 28181 4264
rect 27948 4224 27954 4236
rect 28169 4233 28181 4236
rect 28215 4233 28227 4267
rect 28169 4227 28227 4233
rect 19352 4168 22692 4196
rect 22664 4140 22692 4168
rect 28552 4168 29408 4196
rect 17773 4131 17831 4137
rect 17773 4097 17785 4131
rect 17819 4097 17831 4131
rect 20070 4128 20076 4140
rect 20031 4100 20076 4128
rect 17773 4091 17831 4097
rect 20070 4088 20076 4100
rect 20128 4088 20134 4140
rect 20162 4088 20168 4140
rect 20220 4128 20226 4140
rect 21266 4128 21272 4140
rect 20220 4100 20265 4128
rect 21227 4100 21272 4128
rect 20220 4088 20226 4100
rect 21266 4088 21272 4100
rect 21324 4088 21330 4140
rect 21910 4088 21916 4140
rect 21968 4128 21974 4140
rect 22005 4131 22063 4137
rect 22005 4128 22017 4131
rect 21968 4100 22017 4128
rect 21968 4088 21974 4100
rect 22005 4097 22017 4100
rect 22051 4097 22063 4131
rect 22646 4128 22652 4140
rect 22607 4100 22652 4128
rect 22005 4091 22063 4097
rect 22646 4088 22652 4100
rect 22704 4088 22710 4140
rect 23198 4088 23204 4140
rect 23256 4128 23262 4140
rect 23293 4131 23351 4137
rect 23293 4128 23305 4131
rect 23256 4100 23305 4128
rect 23256 4088 23262 4100
rect 23293 4097 23305 4100
rect 23339 4128 23351 4131
rect 23474 4128 23480 4140
rect 23339 4100 23480 4128
rect 23339 4097 23351 4100
rect 23293 4091 23351 4097
rect 23474 4088 23480 4100
rect 23532 4088 23538 4140
rect 24486 4128 24492 4140
rect 24447 4100 24492 4128
rect 24486 4088 24492 4100
rect 24544 4088 24550 4140
rect 24581 4131 24639 4137
rect 24581 4097 24593 4131
rect 24627 4128 24639 4131
rect 24670 4128 24676 4140
rect 24627 4100 24676 4128
rect 24627 4097 24639 4100
rect 24581 4091 24639 4097
rect 24670 4088 24676 4100
rect 24728 4088 24734 4140
rect 25317 4131 25375 4137
rect 25317 4128 25329 4131
rect 24780 4100 25329 4128
rect 10502 4020 10508 4072
rect 10560 4060 10566 4072
rect 11606 4060 11612 4072
rect 10560 4032 11612 4060
rect 10560 4020 10566 4032
rect 11606 4020 11612 4032
rect 11664 4060 11670 4072
rect 12713 4063 12771 4069
rect 12713 4060 12725 4063
rect 11664 4032 12725 4060
rect 11664 4020 11670 4032
rect 12713 4029 12725 4032
rect 12759 4029 12771 4063
rect 12986 4060 12992 4072
rect 12947 4032 12992 4060
rect 12713 4023 12771 4029
rect 1581 3995 1639 4001
rect 1581 3961 1593 3995
rect 1627 3992 1639 3995
rect 1670 3992 1676 4004
rect 1627 3964 1676 3992
rect 1627 3961 1639 3964
rect 1581 3955 1639 3961
rect 1670 3952 1676 3964
rect 1728 3952 1734 4004
rect 12728 3924 12756 4023
rect 12986 4020 12992 4032
rect 13044 4020 13050 4072
rect 13446 4020 13452 4072
rect 13504 4060 13510 4072
rect 18049 4063 18107 4069
rect 18049 4060 18061 4063
rect 13504 4032 14228 4060
rect 13504 4020 13510 4032
rect 14200 3992 14228 4032
rect 17880 4032 18061 4060
rect 17880 3992 17908 4032
rect 18049 4029 18061 4032
rect 18095 4029 18107 4063
rect 18049 4023 18107 4029
rect 19058 4020 19064 4072
rect 19116 4060 19122 4072
rect 19521 4063 19579 4069
rect 19521 4060 19533 4063
rect 19116 4032 19533 4060
rect 19116 4020 19122 4032
rect 19521 4029 19533 4032
rect 19567 4029 19579 4063
rect 24394 4060 24400 4072
rect 19521 4023 19579 4029
rect 19628 4032 24400 4060
rect 14200 3964 17908 3992
rect 14274 3924 14280 3936
rect 12728 3896 14280 3924
rect 14274 3884 14280 3896
rect 14332 3884 14338 3936
rect 14461 3927 14519 3933
rect 14461 3893 14473 3927
rect 14507 3924 14519 3927
rect 14642 3924 14648 3936
rect 14507 3896 14648 3924
rect 14507 3893 14519 3896
rect 14461 3887 14519 3893
rect 14642 3884 14648 3896
rect 14700 3884 14706 3936
rect 14734 3884 14740 3936
rect 14792 3924 14798 3936
rect 17770 3924 17776 3936
rect 14792 3896 17776 3924
rect 14792 3884 14798 3896
rect 17770 3884 17776 3896
rect 17828 3884 17834 3936
rect 17880 3924 17908 3964
rect 19628 3924 19656 4032
rect 24394 4020 24400 4032
rect 24452 4020 24458 4072
rect 24504 4060 24532 4088
rect 24780 4060 24808 4100
rect 25317 4097 25329 4100
rect 25363 4097 25375 4131
rect 25317 4091 25375 4097
rect 25961 4131 26019 4137
rect 25961 4097 25973 4131
rect 26007 4097 26019 4131
rect 25961 4091 26019 4097
rect 25976 4060 26004 4091
rect 26142 4088 26148 4140
rect 26200 4128 26206 4140
rect 26605 4131 26663 4137
rect 26605 4128 26617 4131
rect 26200 4100 26617 4128
rect 26200 4088 26206 4100
rect 26605 4097 26617 4100
rect 26651 4097 26663 4131
rect 27341 4131 27399 4137
rect 27341 4128 27353 4131
rect 26605 4091 26663 4097
rect 26712 4100 27353 4128
rect 24504 4032 24808 4060
rect 25148 4032 26004 4060
rect 21361 3995 21419 4001
rect 21361 3961 21373 3995
rect 21407 3992 21419 3995
rect 23474 3992 23480 4004
rect 21407 3964 23480 3992
rect 21407 3961 21419 3964
rect 21361 3955 21419 3961
rect 23474 3952 23480 3964
rect 23532 3952 23538 4004
rect 25148 4001 25176 4032
rect 25133 3995 25191 4001
rect 25133 3961 25145 3995
rect 25179 3961 25191 3995
rect 25133 3955 25191 3961
rect 25406 3952 25412 4004
rect 25464 3992 25470 4004
rect 26421 3995 26479 4001
rect 26421 3992 26433 3995
rect 25464 3964 26433 3992
rect 25464 3952 25470 3964
rect 26421 3961 26433 3964
rect 26467 3961 26479 3995
rect 26421 3955 26479 3961
rect 17880 3896 19656 3924
rect 20714 3884 20720 3936
rect 20772 3924 20778 3936
rect 22097 3927 22155 3933
rect 22097 3924 22109 3927
rect 20772 3896 22109 3924
rect 20772 3884 20778 3896
rect 22097 3893 22109 3896
rect 22143 3893 22155 3927
rect 22097 3887 22155 3893
rect 22186 3884 22192 3936
rect 22244 3924 22250 3936
rect 22741 3927 22799 3933
rect 22741 3924 22753 3927
rect 22244 3896 22753 3924
rect 22244 3884 22250 3896
rect 22741 3893 22753 3896
rect 22787 3893 22799 3927
rect 22741 3887 22799 3893
rect 22830 3884 22836 3936
rect 22888 3924 22894 3936
rect 23385 3927 23443 3933
rect 23385 3924 23397 3927
rect 22888 3896 23397 3924
rect 22888 3884 22894 3896
rect 23385 3893 23397 3896
rect 23431 3893 23443 3927
rect 23385 3887 23443 3893
rect 23842 3884 23848 3936
rect 23900 3924 23906 3936
rect 26712 3924 26740 4100
rect 27341 4097 27353 4100
rect 27387 4097 27399 4131
rect 28166 4128 28172 4140
rect 28127 4100 28172 4128
rect 27341 4091 27399 4097
rect 28166 4088 28172 4100
rect 28224 4088 28230 4140
rect 28552 4128 28580 4168
rect 28368 4100 28580 4128
rect 28721 4131 28779 4137
rect 28368 4060 28396 4100
rect 28721 4097 28733 4131
rect 28767 4097 28779 4131
rect 28721 4091 28779 4097
rect 28813 4131 28871 4137
rect 28813 4097 28825 4131
rect 28859 4128 28871 4131
rect 29270 4128 29276 4140
rect 28859 4100 29276 4128
rect 28859 4097 28871 4100
rect 28813 4091 28871 4097
rect 27172 4032 28396 4060
rect 28736 4060 28764 4091
rect 29270 4088 29276 4100
rect 29328 4088 29334 4140
rect 29380 4128 29408 4168
rect 29549 4131 29607 4137
rect 29549 4128 29561 4131
rect 29380 4100 29561 4128
rect 29549 4097 29561 4100
rect 29595 4097 29607 4131
rect 29549 4091 29607 4097
rect 30101 4131 30159 4137
rect 30101 4097 30113 4131
rect 30147 4128 30159 4131
rect 30190 4128 30196 4140
rect 30147 4100 30196 4128
rect 30147 4097 30159 4100
rect 30101 4091 30159 4097
rect 30190 4088 30196 4100
rect 30248 4088 30254 4140
rect 30742 4060 30748 4072
rect 28736 4032 30604 4060
rect 30703 4032 30748 4060
rect 27172 4001 27200 4032
rect 27157 3995 27215 4001
rect 27157 3961 27169 3995
rect 27203 3961 27215 3995
rect 30576 3992 30604 4032
rect 30742 4020 30748 4032
rect 30800 4020 30806 4072
rect 31662 3992 31668 4004
rect 30576 3964 31668 3992
rect 27157 3955 27215 3961
rect 31662 3952 31668 3964
rect 31720 3952 31726 4004
rect 23900 3896 26740 3924
rect 23900 3884 23906 3896
rect 27062 3884 27068 3936
rect 27120 3924 27126 3936
rect 28718 3924 28724 3936
rect 27120 3896 28724 3924
rect 27120 3884 27126 3896
rect 28718 3884 28724 3896
rect 28776 3884 28782 3936
rect 29362 3924 29368 3936
rect 29323 3896 29368 3924
rect 29362 3884 29368 3896
rect 29420 3884 29426 3936
rect 30193 3927 30251 3933
rect 30193 3893 30205 3927
rect 30239 3924 30251 3927
rect 30650 3924 30656 3936
rect 30239 3896 30656 3924
rect 30239 3893 30251 3896
rect 30193 3887 30251 3893
rect 30650 3884 30656 3896
rect 30708 3884 30714 3936
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 1581 3723 1639 3729
rect 1581 3689 1593 3723
rect 1627 3720 1639 3723
rect 1854 3720 1860 3732
rect 1627 3692 1860 3720
rect 1627 3689 1639 3692
rect 1581 3683 1639 3689
rect 1854 3680 1860 3692
rect 1912 3680 1918 3732
rect 7466 3680 7472 3732
rect 7524 3720 7530 3732
rect 9030 3720 9036 3732
rect 7524 3692 9036 3720
rect 7524 3680 7530 3692
rect 9030 3680 9036 3692
rect 9088 3680 9094 3732
rect 10134 3680 10140 3732
rect 10192 3720 10198 3732
rect 11054 3720 11060 3732
rect 10192 3692 11060 3720
rect 10192 3680 10198 3692
rect 11054 3680 11060 3692
rect 11112 3720 11118 3732
rect 15378 3720 15384 3732
rect 11112 3692 15384 3720
rect 11112 3680 11118 3692
rect 15378 3680 15384 3692
rect 15436 3680 15442 3732
rect 17865 3723 17923 3729
rect 17865 3689 17877 3723
rect 17911 3720 17923 3723
rect 18506 3720 18512 3732
rect 17911 3692 18512 3720
rect 17911 3689 17923 3692
rect 17865 3683 17923 3689
rect 18506 3680 18512 3692
rect 18564 3680 18570 3732
rect 18598 3680 18604 3732
rect 18656 3720 18662 3732
rect 24486 3720 24492 3732
rect 18656 3692 24492 3720
rect 18656 3680 18662 3692
rect 24486 3680 24492 3692
rect 24544 3680 24550 3732
rect 25590 3720 25596 3732
rect 25424 3692 25596 3720
rect 6733 3655 6791 3661
rect 6733 3621 6745 3655
rect 6779 3652 6791 3655
rect 11422 3652 11428 3664
rect 6779 3624 11428 3652
rect 6779 3621 6791 3624
rect 6733 3615 6791 3621
rect 11422 3612 11428 3624
rect 11480 3612 11486 3664
rect 12986 3612 12992 3664
rect 13044 3652 13050 3664
rect 14734 3652 14740 3664
rect 13044 3624 14740 3652
rect 13044 3612 13050 3624
rect 14734 3612 14740 3624
rect 14792 3612 14798 3664
rect 17310 3612 17316 3664
rect 17368 3652 17374 3664
rect 25424 3652 25452 3692
rect 25590 3680 25596 3692
rect 25648 3680 25654 3732
rect 25682 3680 25688 3732
rect 25740 3720 25746 3732
rect 25869 3723 25927 3729
rect 25869 3720 25881 3723
rect 25740 3692 25881 3720
rect 25740 3680 25746 3692
rect 25869 3689 25881 3692
rect 25915 3689 25927 3723
rect 25869 3683 25927 3689
rect 26602 3680 26608 3732
rect 26660 3720 26666 3732
rect 26697 3723 26755 3729
rect 26697 3720 26709 3723
rect 26660 3692 26709 3720
rect 26660 3680 26666 3692
rect 26697 3689 26709 3692
rect 26743 3689 26755 3723
rect 30834 3720 30840 3732
rect 30795 3692 30840 3720
rect 26697 3683 26755 3689
rect 30834 3680 30840 3692
rect 30892 3680 30898 3732
rect 33042 3680 33048 3732
rect 33100 3720 33106 3732
rect 38105 3723 38163 3729
rect 38105 3720 38117 3723
rect 33100 3692 38117 3720
rect 33100 3680 33106 3692
rect 38105 3689 38117 3692
rect 38151 3689 38163 3723
rect 38105 3683 38163 3689
rect 17368 3624 25452 3652
rect 17368 3612 17374 3624
rect 28166 3612 28172 3664
rect 28224 3652 28230 3664
rect 37274 3652 37280 3664
rect 28224 3624 37280 3652
rect 28224 3612 28230 3624
rect 37274 3612 37280 3624
rect 37332 3612 37338 3664
rect 4062 3544 4068 3596
rect 4120 3584 4126 3596
rect 4985 3587 5043 3593
rect 4985 3584 4997 3587
rect 4120 3556 4997 3584
rect 4120 3544 4126 3556
rect 4985 3553 4997 3556
rect 5031 3584 5043 3587
rect 7190 3584 7196 3596
rect 5031 3556 7196 3584
rect 5031 3553 5043 3556
rect 4985 3547 5043 3553
rect 7190 3544 7196 3556
rect 7248 3544 7254 3596
rect 14182 3584 14188 3596
rect 8496 3556 14188 3584
rect 1762 3516 1768 3528
rect 1723 3488 1768 3516
rect 1762 3476 1768 3488
rect 1820 3476 1826 3528
rect 8496 3516 8524 3556
rect 14182 3544 14188 3556
rect 14240 3544 14246 3596
rect 15105 3587 15163 3593
rect 15105 3553 15117 3587
rect 15151 3584 15163 3587
rect 15286 3584 15292 3596
rect 15151 3556 15292 3584
rect 15151 3553 15163 3556
rect 15105 3547 15163 3553
rect 15286 3544 15292 3556
rect 15344 3544 15350 3596
rect 15378 3544 15384 3596
rect 15436 3584 15442 3596
rect 20346 3584 20352 3596
rect 15436 3556 20352 3584
rect 15436 3544 15442 3556
rect 20346 3544 20352 3556
rect 20404 3544 20410 3596
rect 25685 3587 25743 3593
rect 20640 3556 21128 3584
rect 14366 3516 14372 3528
rect 6394 3488 8524 3516
rect 8588 3488 14372 3516
rect 5261 3451 5319 3457
rect 5261 3417 5273 3451
rect 5307 3417 5319 3451
rect 5261 3411 5319 3417
rect 5276 3380 5304 3411
rect 7834 3408 7840 3460
rect 7892 3448 7898 3460
rect 8588 3448 8616 3488
rect 14366 3476 14372 3488
rect 14424 3476 14430 3528
rect 15010 3516 15016 3528
rect 14971 3488 15016 3516
rect 15010 3476 15016 3488
rect 15068 3476 15074 3528
rect 17034 3476 17040 3528
rect 17092 3516 17098 3528
rect 17129 3519 17187 3525
rect 17129 3516 17141 3519
rect 17092 3488 17141 3516
rect 17092 3476 17098 3488
rect 17129 3485 17141 3488
rect 17175 3516 17187 3519
rect 17773 3519 17831 3525
rect 17773 3516 17785 3519
rect 17175 3488 17785 3516
rect 17175 3485 17187 3488
rect 17129 3479 17187 3485
rect 17773 3485 17785 3488
rect 17819 3516 17831 3519
rect 18046 3516 18052 3528
rect 17819 3488 18052 3516
rect 17819 3485 17831 3488
rect 17773 3479 17831 3485
rect 18046 3476 18052 3488
rect 18104 3476 18110 3528
rect 18690 3476 18696 3528
rect 18748 3512 18754 3528
rect 18748 3484 18789 3512
rect 18748 3476 18754 3484
rect 18874 3476 18880 3528
rect 18932 3516 18938 3528
rect 19889 3519 19947 3525
rect 19889 3516 19901 3519
rect 18932 3488 19901 3516
rect 18932 3476 18938 3488
rect 19889 3485 19901 3488
rect 19935 3516 19947 3519
rect 20438 3516 20444 3528
rect 19935 3488 20444 3516
rect 19935 3485 19947 3488
rect 19889 3479 19947 3485
rect 20438 3476 20444 3488
rect 20496 3476 20502 3528
rect 20533 3519 20591 3525
rect 20533 3485 20545 3519
rect 20579 3516 20591 3519
rect 20640 3516 20668 3556
rect 21100 3528 21128 3556
rect 25685 3553 25697 3587
rect 25731 3584 25743 3587
rect 29362 3584 29368 3596
rect 25731 3556 29368 3584
rect 25731 3553 25743 3556
rect 25685 3547 25743 3553
rect 29362 3544 29368 3556
rect 29420 3544 29426 3596
rect 30650 3584 30656 3596
rect 30611 3556 30656 3584
rect 30650 3544 30656 3556
rect 30708 3544 30714 3596
rect 20579 3488 20668 3516
rect 20579 3485 20591 3488
rect 20533 3479 20591 3485
rect 21082 3476 21088 3528
rect 21140 3516 21146 3528
rect 21177 3519 21235 3525
rect 21177 3516 21189 3519
rect 21140 3488 21189 3516
rect 21140 3476 21146 3488
rect 21177 3485 21189 3488
rect 21223 3485 21235 3519
rect 21177 3479 21235 3485
rect 22373 3519 22431 3525
rect 22373 3485 22385 3519
rect 22419 3516 22431 3519
rect 22462 3516 22468 3528
rect 22419 3488 22468 3516
rect 22419 3485 22431 3488
rect 22373 3479 22431 3485
rect 22462 3476 22468 3488
rect 22520 3476 22526 3528
rect 22649 3519 22707 3525
rect 22649 3485 22661 3519
rect 22695 3516 22707 3519
rect 23198 3516 23204 3528
rect 22695 3488 23204 3516
rect 22695 3485 22707 3488
rect 22649 3479 22707 3485
rect 23198 3476 23204 3488
rect 23256 3476 23262 3528
rect 24578 3516 24584 3528
rect 24539 3488 24584 3516
rect 24578 3476 24584 3488
rect 24636 3476 24642 3528
rect 25509 3519 25567 3525
rect 25509 3485 25521 3519
rect 25555 3516 25567 3519
rect 25774 3516 25780 3528
rect 25555 3488 25780 3516
rect 25555 3485 25567 3488
rect 25509 3479 25567 3485
rect 25774 3476 25780 3488
rect 25832 3476 25838 3528
rect 26418 3476 26424 3528
rect 26476 3516 26482 3528
rect 26605 3519 26663 3525
rect 26605 3516 26617 3519
rect 26476 3488 26617 3516
rect 26476 3476 26482 3488
rect 26605 3485 26617 3488
rect 26651 3485 26663 3519
rect 26605 3479 26663 3485
rect 27249 3519 27307 3525
rect 27249 3485 27261 3519
rect 27295 3516 27307 3519
rect 27798 3516 27804 3528
rect 27295 3488 27804 3516
rect 27295 3485 27307 3488
rect 27249 3479 27307 3485
rect 27798 3476 27804 3488
rect 27856 3476 27862 3528
rect 28074 3516 28080 3528
rect 28035 3488 28080 3516
rect 28074 3476 28080 3488
rect 28132 3476 28138 3528
rect 29733 3519 29791 3525
rect 29733 3485 29745 3519
rect 29779 3485 29791 3519
rect 29733 3479 29791 3485
rect 30469 3519 30527 3525
rect 30469 3485 30481 3519
rect 30515 3485 30527 3519
rect 30469 3479 30527 3485
rect 18693 3475 18751 3476
rect 7892 3420 8616 3448
rect 7892 3408 7898 3420
rect 9030 3408 9036 3460
rect 9088 3448 9094 3460
rect 14458 3448 14464 3460
rect 9088 3420 14464 3448
rect 9088 3408 9094 3420
rect 14458 3408 14464 3420
rect 14516 3408 14522 3460
rect 18966 3408 18972 3460
rect 19024 3448 19030 3460
rect 20625 3451 20683 3457
rect 20625 3448 20637 3451
rect 19024 3420 20637 3448
rect 19024 3408 19030 3420
rect 20625 3417 20637 3420
rect 20671 3417 20683 3451
rect 23382 3448 23388 3460
rect 23343 3420 23388 3448
rect 20625 3411 20683 3417
rect 23382 3408 23388 3420
rect 23440 3408 23446 3460
rect 23474 3408 23480 3460
rect 23532 3448 23538 3460
rect 24026 3448 24032 3460
rect 23532 3420 23577 3448
rect 23987 3420 24032 3448
rect 23532 3408 23538 3420
rect 24026 3408 24032 3420
rect 24084 3408 24090 3460
rect 24394 3408 24400 3460
rect 24452 3448 24458 3460
rect 24452 3420 25544 3448
rect 24452 3408 24458 3420
rect 11514 3380 11520 3392
rect 5276 3352 11520 3380
rect 11514 3340 11520 3352
rect 11572 3340 11578 3392
rect 14366 3340 14372 3392
rect 14424 3380 14430 3392
rect 15746 3380 15752 3392
rect 14424 3352 15752 3380
rect 14424 3340 14430 3352
rect 15746 3340 15752 3352
rect 15804 3340 15810 3392
rect 17218 3380 17224 3392
rect 17179 3352 17224 3380
rect 17218 3340 17224 3352
rect 17276 3340 17282 3392
rect 18138 3340 18144 3392
rect 18196 3380 18202 3392
rect 18509 3383 18567 3389
rect 18509 3380 18521 3383
rect 18196 3352 18521 3380
rect 18196 3340 18202 3352
rect 18509 3349 18521 3352
rect 18555 3349 18567 3383
rect 19978 3380 19984 3392
rect 19939 3352 19984 3380
rect 18509 3343 18567 3349
rect 19978 3340 19984 3352
rect 20036 3340 20042 3392
rect 20162 3340 20168 3392
rect 20220 3380 20226 3392
rect 21269 3383 21327 3389
rect 21269 3380 21281 3383
rect 20220 3352 21281 3380
rect 20220 3340 20226 3352
rect 21269 3349 21281 3352
rect 21315 3349 21327 3383
rect 21269 3343 21327 3349
rect 21358 3340 21364 3392
rect 21416 3380 21422 3392
rect 23842 3380 23848 3392
rect 21416 3352 23848 3380
rect 21416 3340 21422 3352
rect 23842 3340 23848 3352
rect 23900 3340 23906 3392
rect 24118 3340 24124 3392
rect 24176 3380 24182 3392
rect 24673 3383 24731 3389
rect 24673 3380 24685 3383
rect 24176 3352 24685 3380
rect 24176 3340 24182 3352
rect 24673 3349 24685 3352
rect 24719 3349 24731 3383
rect 25516 3380 25544 3420
rect 25590 3408 25596 3460
rect 25648 3448 25654 3460
rect 29748 3448 29776 3479
rect 30484 3448 30512 3479
rect 31018 3476 31024 3528
rect 31076 3516 31082 3528
rect 31757 3519 31815 3525
rect 31757 3516 31769 3519
rect 31076 3488 31769 3516
rect 31076 3476 31082 3488
rect 31757 3485 31769 3488
rect 31803 3485 31815 3519
rect 31757 3479 31815 3485
rect 32217 3519 32275 3525
rect 32217 3485 32229 3519
rect 32263 3516 32275 3519
rect 33686 3516 33692 3528
rect 32263 3488 33692 3516
rect 32263 3485 32275 3488
rect 32217 3479 32275 3485
rect 33686 3476 33692 3488
rect 33744 3476 33750 3528
rect 38286 3516 38292 3528
rect 38247 3488 38292 3516
rect 38286 3476 38292 3488
rect 38344 3476 38350 3528
rect 32309 3451 32367 3457
rect 32309 3448 32321 3451
rect 25648 3420 30420 3448
rect 30484 3420 32321 3448
rect 25648 3408 25654 3420
rect 27062 3380 27068 3392
rect 25516 3352 27068 3380
rect 24673 3343 24731 3349
rect 27062 3340 27068 3352
rect 27120 3340 27126 3392
rect 27338 3380 27344 3392
rect 27299 3352 27344 3380
rect 27338 3340 27344 3352
rect 27396 3340 27402 3392
rect 27890 3380 27896 3392
rect 27851 3352 27896 3380
rect 27890 3340 27896 3352
rect 27948 3340 27954 3392
rect 28534 3380 28540 3392
rect 28495 3352 28540 3380
rect 28534 3340 28540 3352
rect 28592 3340 28598 3392
rect 28810 3340 28816 3392
rect 28868 3380 28874 3392
rect 29825 3383 29883 3389
rect 29825 3380 29837 3383
rect 28868 3352 29837 3380
rect 28868 3340 28874 3352
rect 29825 3349 29837 3352
rect 29871 3349 29883 3383
rect 30392 3380 30420 3420
rect 32309 3417 32321 3420
rect 32355 3417 32367 3451
rect 32309 3411 32367 3417
rect 31202 3380 31208 3392
rect 30392 3352 31208 3380
rect 29825 3343 29883 3349
rect 31202 3340 31208 3352
rect 31260 3340 31266 3392
rect 31570 3380 31576 3392
rect 31531 3352 31576 3380
rect 31570 3340 31576 3352
rect 31628 3340 31634 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 2317 3179 2375 3185
rect 2317 3145 2329 3179
rect 2363 3145 2375 3179
rect 2317 3139 2375 3145
rect 1581 3043 1639 3049
rect 1581 3009 1593 3043
rect 1627 3040 1639 3043
rect 2332 3040 2360 3139
rect 5810 3136 5816 3188
rect 5868 3176 5874 3188
rect 5905 3179 5963 3185
rect 5905 3176 5917 3179
rect 5868 3148 5917 3176
rect 5868 3136 5874 3148
rect 5905 3145 5917 3148
rect 5951 3145 5963 3179
rect 13446 3176 13452 3188
rect 13407 3148 13452 3176
rect 5905 3139 5963 3145
rect 13446 3136 13452 3148
rect 13504 3136 13510 3188
rect 17218 3176 17224 3188
rect 14016 3148 17224 3176
rect 6638 3108 6644 3120
rect 5658 3080 6644 3108
rect 6638 3068 6644 3080
rect 6696 3068 6702 3120
rect 7193 3111 7251 3117
rect 7193 3077 7205 3111
rect 7239 3108 7251 3111
rect 7466 3108 7472 3120
rect 7239 3080 7472 3108
rect 7239 3077 7251 3080
rect 7193 3071 7251 3077
rect 7466 3068 7472 3080
rect 7524 3068 7530 3120
rect 9674 3108 9680 3120
rect 8418 3080 9680 3108
rect 9674 3068 9680 3080
rect 9732 3068 9738 3120
rect 11149 3111 11207 3117
rect 11149 3077 11161 3111
rect 11195 3108 11207 3111
rect 11514 3108 11520 3120
rect 11195 3080 11520 3108
rect 11195 3077 11207 3080
rect 11149 3071 11207 3077
rect 11514 3068 11520 3080
rect 11572 3068 11578 3120
rect 11977 3111 12035 3117
rect 11977 3077 11989 3111
rect 12023 3108 12035 3111
rect 12066 3108 12072 3120
rect 12023 3080 12072 3108
rect 12023 3077 12035 3080
rect 11977 3071 12035 3077
rect 12066 3068 12072 3080
rect 12124 3068 12130 3120
rect 14016 3108 14044 3148
rect 17218 3136 17224 3148
rect 17276 3136 17282 3188
rect 20625 3179 20683 3185
rect 20625 3176 20637 3179
rect 17972 3148 20637 3176
rect 14274 3108 14280 3120
rect 13202 3080 14044 3108
rect 14108 3080 14280 3108
rect 2498 3040 2504 3052
rect 1627 3012 2360 3040
rect 2459 3012 2504 3040
rect 1627 3009 1639 3012
rect 1581 3003 1639 3009
rect 2498 3000 2504 3012
rect 2556 3000 2562 3052
rect 3326 3040 3332 3052
rect 3287 3012 3332 3040
rect 3326 3000 3332 3012
rect 3384 3000 3390 3052
rect 4062 3000 4068 3052
rect 4120 3040 4126 3052
rect 4157 3043 4215 3049
rect 4157 3040 4169 3043
rect 4120 3012 4169 3040
rect 4120 3000 4126 3012
rect 4157 3009 4169 3012
rect 4203 3009 4215 3043
rect 4157 3003 4215 3009
rect 6917 3043 6975 3049
rect 6917 3009 6929 3043
rect 6963 3009 6975 3043
rect 9122 3040 9128 3052
rect 9083 3012 9128 3040
rect 6917 3003 6975 3009
rect 4433 2975 4491 2981
rect 4433 2941 4445 2975
rect 4479 2972 4491 2975
rect 5442 2972 5448 2984
rect 4479 2944 5448 2972
rect 4479 2941 4491 2944
rect 4433 2935 4491 2941
rect 5442 2932 5448 2944
rect 5500 2932 5506 2984
rect 6932 2972 6960 3003
rect 9122 3000 9128 3012
rect 9180 3000 9186 3052
rect 14108 3049 14136 3080
rect 14274 3068 14280 3080
rect 14332 3068 14338 3120
rect 14366 3068 14372 3120
rect 14424 3108 14430 3120
rect 17862 3108 17868 3120
rect 14424 3080 14469 3108
rect 15594 3080 17868 3108
rect 14424 3068 14430 3080
rect 17862 3068 17868 3080
rect 17920 3068 17926 3120
rect 14093 3043 14151 3049
rect 7190 2972 7196 2984
rect 6932 2944 7196 2972
rect 7190 2932 7196 2944
rect 7248 2972 7254 2984
rect 9140 2972 9168 3000
rect 7248 2944 9168 2972
rect 9401 2975 9459 2981
rect 7248 2932 7254 2944
rect 9401 2941 9413 2975
rect 9447 2972 9459 2975
rect 10042 2972 10048 2984
rect 9447 2944 10048 2972
rect 9447 2941 9459 2944
rect 9401 2935 9459 2941
rect 10042 2932 10048 2944
rect 10100 2932 10106 2984
rect 14 2796 20 2848
rect 72 2836 78 2848
rect 1765 2839 1823 2845
rect 1765 2836 1777 2839
rect 72 2808 1777 2836
rect 72 2796 78 2808
rect 1765 2805 1777 2808
rect 1811 2805 1823 2839
rect 1765 2799 1823 2805
rect 3145 2839 3203 2845
rect 3145 2805 3157 2839
rect 3191 2836 3203 2839
rect 5810 2836 5816 2848
rect 3191 2808 5816 2836
rect 3191 2805 3203 2808
rect 3145 2799 3203 2805
rect 5810 2796 5816 2808
rect 5868 2796 5874 2848
rect 8665 2839 8723 2845
rect 8665 2805 8677 2839
rect 8711 2836 8723 2839
rect 10134 2836 10140 2848
rect 8711 2808 10140 2836
rect 8711 2805 8723 2808
rect 8665 2799 8723 2805
rect 10134 2796 10140 2808
rect 10192 2796 10198 2848
rect 10520 2836 10548 3026
rect 14093 3009 14105 3043
rect 14139 3009 14151 3043
rect 17972 3040 18000 3148
rect 20625 3145 20637 3148
rect 20671 3176 20683 3179
rect 21266 3176 21272 3188
rect 20671 3148 21272 3176
rect 20671 3145 20683 3148
rect 20625 3139 20683 3145
rect 21266 3136 21272 3148
rect 21324 3136 21330 3188
rect 23293 3179 23351 3185
rect 23293 3145 23305 3179
rect 23339 3176 23351 3179
rect 23382 3176 23388 3188
rect 23339 3148 23388 3176
rect 23339 3145 23351 3148
rect 23293 3139 23351 3145
rect 23382 3136 23388 3148
rect 23440 3136 23446 3188
rect 27801 3179 27859 3185
rect 27801 3176 27813 3179
rect 25056 3148 27813 3176
rect 18233 3111 18291 3117
rect 18233 3077 18245 3111
rect 18279 3108 18291 3111
rect 18279 3080 19642 3108
rect 18279 3077 18291 3080
rect 18233 3071 18291 3077
rect 20806 3068 20812 3120
rect 20864 3108 20870 3120
rect 21361 3111 21419 3117
rect 21361 3108 21373 3111
rect 20864 3080 21373 3108
rect 20864 3068 20870 3080
rect 21361 3077 21373 3080
rect 21407 3077 21419 3111
rect 22186 3108 22192 3120
rect 22147 3080 22192 3108
rect 21361 3071 21419 3077
rect 22186 3068 22192 3080
rect 22244 3068 22250 3120
rect 22741 3111 22799 3117
rect 22741 3077 22753 3111
rect 22787 3108 22799 3111
rect 23566 3108 23572 3120
rect 22787 3080 23572 3108
rect 22787 3077 22799 3080
rect 22741 3071 22799 3077
rect 23566 3068 23572 3080
rect 23624 3068 23630 3120
rect 14093 3003 14151 3009
rect 16040 3012 18000 3040
rect 11701 2975 11759 2981
rect 11701 2941 11713 2975
rect 11747 2972 11759 2975
rect 14108 2972 14136 3003
rect 11747 2944 14136 2972
rect 11747 2941 11759 2944
rect 11701 2935 11759 2941
rect 14458 2932 14464 2984
rect 14516 2972 14522 2984
rect 16040 2972 16068 3012
rect 18046 3000 18052 3052
rect 18104 3040 18110 3052
rect 18141 3043 18199 3049
rect 18141 3040 18153 3043
rect 18104 3012 18153 3040
rect 18104 3000 18110 3012
rect 18141 3009 18153 3012
rect 18187 3009 18199 3043
rect 18141 3003 18199 3009
rect 14516 2944 16068 2972
rect 14516 2932 14522 2944
rect 16114 2932 16120 2984
rect 16172 2972 16178 2984
rect 18156 2972 18184 3003
rect 18322 3000 18328 3052
rect 18380 3040 18386 3052
rect 18877 3043 18935 3049
rect 18877 3040 18889 3043
rect 18380 3012 18889 3040
rect 18380 3000 18386 3012
rect 18877 3009 18889 3012
rect 18923 3009 18935 3043
rect 18877 3003 18935 3009
rect 21269 3043 21327 3049
rect 21269 3009 21281 3043
rect 21315 3040 21327 3043
rect 21910 3040 21916 3052
rect 21315 3012 21916 3040
rect 21315 3009 21327 3012
rect 21269 3003 21327 3009
rect 21910 3000 21916 3012
rect 21968 3000 21974 3052
rect 23201 3043 23259 3049
rect 23201 3009 23213 3043
rect 23247 3009 23259 3043
rect 24118 3040 24124 3052
rect 24079 3012 24124 3040
rect 23201 3003 23259 3009
rect 18782 2972 18788 2984
rect 16172 2944 16217 2972
rect 18156 2944 18788 2972
rect 16172 2932 16178 2944
rect 18782 2932 18788 2944
rect 18840 2932 18846 2984
rect 19150 2972 19156 2984
rect 19111 2944 19156 2972
rect 19150 2932 19156 2944
rect 19208 2932 19214 2984
rect 22094 2932 22100 2984
rect 22152 2972 22158 2984
rect 23216 2972 23244 3003
rect 24118 3000 24124 3012
rect 24176 3000 24182 3052
rect 25056 3049 25084 3148
rect 27801 3145 27813 3148
rect 27847 3145 27859 3179
rect 31018 3176 31024 3188
rect 30979 3148 31024 3176
rect 27801 3139 27859 3145
rect 31018 3136 31024 3148
rect 31076 3136 31082 3188
rect 36722 3176 36728 3188
rect 36683 3148 36728 3176
rect 36722 3136 36728 3148
rect 36780 3136 36786 3188
rect 25133 3111 25191 3117
rect 25133 3077 25145 3111
rect 25179 3108 25191 3111
rect 26142 3108 26148 3120
rect 25179 3080 26148 3108
rect 25179 3077 25191 3080
rect 25133 3071 25191 3077
rect 26142 3068 26148 3080
rect 26200 3068 26206 3120
rect 28534 3108 28540 3120
rect 27172 3080 28540 3108
rect 27172 3049 27200 3080
rect 28534 3068 28540 3080
rect 28592 3068 28598 3120
rect 28810 3108 28816 3120
rect 28771 3080 28816 3108
rect 28810 3068 28816 3080
rect 28868 3068 28874 3120
rect 30009 3111 30067 3117
rect 30009 3077 30021 3111
rect 30055 3108 30067 3111
rect 31570 3108 31576 3120
rect 30055 3080 31576 3108
rect 30055 3077 30067 3080
rect 30009 3071 30067 3077
rect 31570 3068 31576 3080
rect 31628 3068 31634 3120
rect 32950 3068 32956 3120
rect 33008 3108 33014 3120
rect 33008 3080 38056 3108
rect 33008 3068 33014 3080
rect 24581 3043 24639 3049
rect 24581 3009 24593 3043
rect 24627 3040 24639 3043
rect 25041 3043 25099 3049
rect 25041 3040 25053 3043
rect 24627 3012 25053 3040
rect 24627 3009 24639 3012
rect 24581 3003 24639 3009
rect 25041 3009 25053 3012
rect 25087 3009 25099 3043
rect 25041 3003 25099 3009
rect 26053 3043 26111 3049
rect 26053 3009 26065 3043
rect 26099 3009 26111 3043
rect 26053 3003 26111 3009
rect 27157 3043 27215 3049
rect 27157 3009 27169 3043
rect 27203 3009 27215 3043
rect 27157 3003 27215 3009
rect 27341 3043 27399 3049
rect 27341 3009 27353 3043
rect 27387 3040 27399 3043
rect 27890 3040 27896 3052
rect 27387 3012 27896 3040
rect 27387 3009 27399 3012
rect 27341 3003 27399 3009
rect 22152 2944 22197 2972
rect 22572 2944 23244 2972
rect 23937 2975 23995 2981
rect 22152 2932 22158 2944
rect 13372 2876 13584 2904
rect 13372 2836 13400 2876
rect 10520 2808 13400 2836
rect 13556 2836 13584 2876
rect 15746 2864 15752 2916
rect 15804 2904 15810 2916
rect 18598 2904 18604 2916
rect 15804 2876 18604 2904
rect 15804 2864 15810 2876
rect 18598 2864 18604 2876
rect 18656 2864 18662 2916
rect 20714 2864 20720 2916
rect 20772 2904 20778 2916
rect 22572 2904 22600 2944
rect 23937 2941 23949 2975
rect 23983 2972 23995 2975
rect 24026 2972 24032 2984
rect 23983 2944 24032 2972
rect 23983 2941 23995 2944
rect 23937 2935 23995 2941
rect 20772 2876 22600 2904
rect 20772 2864 20778 2876
rect 20162 2836 20168 2848
rect 13556 2808 20168 2836
rect 20162 2796 20168 2808
rect 20220 2796 20226 2848
rect 20530 2796 20536 2848
rect 20588 2836 20594 2848
rect 23952 2836 23980 2935
rect 24026 2932 24032 2944
rect 24084 2932 24090 2984
rect 26068 2972 26096 3003
rect 27890 3000 27896 3012
rect 27948 3000 27954 3052
rect 27982 3000 27988 3052
rect 28040 3040 28046 3052
rect 31202 3040 31208 3052
rect 28040 3012 28580 3040
rect 31163 3012 31208 3040
rect 28040 3000 28046 3012
rect 28552 2972 28580 3012
rect 31202 3000 31208 3012
rect 31260 3000 31266 3052
rect 32490 3040 32496 3052
rect 32451 3012 32496 3040
rect 32490 3000 32496 3012
rect 32548 3000 32554 3052
rect 38028 3049 38056 3080
rect 36909 3043 36967 3049
rect 36909 3009 36921 3043
rect 36955 3009 36967 3043
rect 36909 3003 36967 3009
rect 38013 3043 38071 3049
rect 38013 3009 38025 3043
rect 38059 3009 38071 3043
rect 38013 3003 38071 3009
rect 28721 2975 28779 2981
rect 28721 2972 28733 2975
rect 26068 2944 28488 2972
rect 28552 2944 28733 2972
rect 25682 2864 25688 2916
rect 25740 2904 25746 2916
rect 25740 2876 27200 2904
rect 25740 2864 25746 2876
rect 20588 2808 23980 2836
rect 26053 2839 26111 2845
rect 20588 2796 20594 2808
rect 26053 2805 26065 2839
rect 26099 2836 26111 2839
rect 27062 2836 27068 2848
rect 26099 2808 27068 2836
rect 26099 2805 26111 2808
rect 26053 2799 26111 2805
rect 27062 2796 27068 2808
rect 27120 2796 27126 2848
rect 27172 2836 27200 2876
rect 27246 2864 27252 2916
rect 27304 2904 27310 2916
rect 28460 2904 28488 2944
rect 28721 2941 28733 2944
rect 28767 2941 28779 2975
rect 28721 2935 28779 2941
rect 28997 2975 29055 2981
rect 28997 2941 29009 2975
rect 29043 2941 29055 2975
rect 28997 2935 29055 2941
rect 29917 2975 29975 2981
rect 29917 2941 29929 2975
rect 29963 2972 29975 2975
rect 30742 2972 30748 2984
rect 29963 2944 30748 2972
rect 29963 2941 29975 2944
rect 29917 2935 29975 2941
rect 29012 2904 29040 2935
rect 30742 2932 30748 2944
rect 30800 2932 30806 2984
rect 36924 2972 36952 3003
rect 39298 2972 39304 2984
rect 36924 2944 39304 2972
rect 39298 2932 39304 2944
rect 39356 2932 39362 2984
rect 30469 2907 30527 2913
rect 30469 2904 30481 2907
rect 27304 2876 27936 2904
rect 28460 2876 30481 2904
rect 27304 2864 27310 2876
rect 27798 2836 27804 2848
rect 27172 2808 27804 2836
rect 27798 2796 27804 2808
rect 27856 2796 27862 2848
rect 27908 2836 27936 2876
rect 30469 2873 30481 2876
rect 30515 2873 30527 2907
rect 30469 2867 30527 2873
rect 30576 2876 31754 2904
rect 29914 2836 29920 2848
rect 27908 2808 29920 2836
rect 29914 2796 29920 2808
rect 29972 2796 29978 2848
rect 30282 2796 30288 2848
rect 30340 2836 30346 2848
rect 30576 2836 30604 2876
rect 30340 2808 30604 2836
rect 31726 2848 31754 2876
rect 31726 2808 31760 2848
rect 30340 2796 30346 2808
rect 31754 2796 31760 2808
rect 31812 2796 31818 2848
rect 32306 2836 32312 2848
rect 32267 2808 32312 2836
rect 32306 2796 32312 2808
rect 32364 2796 32370 2848
rect 38194 2836 38200 2848
rect 38155 2808 38200 2836
rect 38194 2796 38200 2808
rect 38252 2796 38258 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 2406 2592 2412 2644
rect 2464 2632 2470 2644
rect 2593 2635 2651 2641
rect 2593 2632 2605 2635
rect 2464 2604 2605 2632
rect 2464 2592 2470 2604
rect 2593 2601 2605 2604
rect 2639 2601 2651 2635
rect 2593 2595 2651 2601
rect 3237 2635 3295 2641
rect 3237 2601 3249 2635
rect 3283 2632 3295 2635
rect 7374 2632 7380 2644
rect 3283 2604 7380 2632
rect 3283 2601 3295 2604
rect 3237 2595 3295 2601
rect 7374 2592 7380 2604
rect 7432 2592 7438 2644
rect 7466 2592 7472 2644
rect 7524 2632 7530 2644
rect 10318 2632 10324 2644
rect 7524 2604 10324 2632
rect 7524 2592 7530 2604
rect 10318 2592 10324 2604
rect 10376 2592 10382 2644
rect 14277 2635 14335 2641
rect 14277 2601 14289 2635
rect 14323 2632 14335 2635
rect 15010 2632 15016 2644
rect 14323 2604 15016 2632
rect 14323 2601 14335 2604
rect 14277 2595 14335 2601
rect 15010 2592 15016 2604
rect 15068 2592 15074 2644
rect 17954 2632 17960 2644
rect 16546 2604 17960 2632
rect 5721 2567 5779 2573
rect 5721 2533 5733 2567
rect 5767 2564 5779 2567
rect 7006 2564 7012 2576
rect 5767 2536 7012 2564
rect 5767 2533 5779 2536
rect 5721 2527 5779 2533
rect 7006 2524 7012 2536
rect 7064 2524 7070 2576
rect 16546 2564 16574 2604
rect 17954 2592 17960 2604
rect 18012 2592 18018 2644
rect 18046 2592 18052 2644
rect 18104 2632 18110 2644
rect 20257 2635 20315 2641
rect 20257 2632 20269 2635
rect 18104 2604 20269 2632
rect 18104 2592 18110 2604
rect 20257 2601 20269 2604
rect 20303 2601 20315 2635
rect 20257 2595 20315 2601
rect 22094 2592 22100 2644
rect 22152 2632 22158 2644
rect 22189 2635 22247 2641
rect 22189 2632 22201 2635
rect 22152 2604 22201 2632
rect 22152 2592 22158 2604
rect 22189 2601 22201 2604
rect 22235 2601 22247 2635
rect 22189 2595 22247 2601
rect 23017 2635 23075 2641
rect 23017 2601 23029 2635
rect 23063 2632 23075 2635
rect 23750 2632 23756 2644
rect 23063 2604 23756 2632
rect 23063 2601 23075 2604
rect 23017 2595 23075 2601
rect 23750 2592 23756 2604
rect 23808 2592 23814 2644
rect 25498 2592 25504 2644
rect 25556 2632 25562 2644
rect 25869 2635 25927 2641
rect 25869 2632 25881 2635
rect 25556 2604 25881 2632
rect 25556 2592 25562 2604
rect 25869 2601 25881 2604
rect 25915 2601 25927 2635
rect 25869 2595 25927 2601
rect 26206 2604 28028 2632
rect 7300 2536 16574 2564
rect 2866 2496 2872 2508
rect 1596 2468 2872 2496
rect 1596 2437 1624 2468
rect 2866 2456 2872 2468
rect 2924 2456 2930 2508
rect 3970 2496 3976 2508
rect 3931 2468 3976 2496
rect 3970 2456 3976 2468
rect 4028 2456 4034 2508
rect 4249 2499 4307 2505
rect 4249 2465 4261 2499
rect 4295 2496 4307 2499
rect 7190 2496 7196 2508
rect 4295 2468 7196 2496
rect 4295 2465 4307 2468
rect 4249 2459 4307 2465
rect 7190 2456 7196 2468
rect 7248 2456 7254 2508
rect 1581 2431 1639 2437
rect 1581 2397 1593 2431
rect 1627 2397 1639 2431
rect 1581 2391 1639 2397
rect 2590 2388 2596 2440
rect 2648 2428 2654 2440
rect 2777 2431 2835 2437
rect 2777 2428 2789 2431
rect 2648 2400 2789 2428
rect 2648 2388 2654 2400
rect 2777 2397 2789 2400
rect 2823 2397 2835 2431
rect 2777 2391 2835 2397
rect 3421 2431 3479 2437
rect 3421 2397 3433 2431
rect 3467 2397 3479 2431
rect 3421 2391 3479 2397
rect 1302 2252 1308 2304
rect 1360 2292 1366 2304
rect 1765 2295 1823 2301
rect 1765 2292 1777 2295
rect 1360 2264 1777 2292
rect 1360 2252 1366 2264
rect 1765 2261 1777 2264
rect 1811 2261 1823 2295
rect 3436 2292 3464 2391
rect 5810 2388 5816 2440
rect 5868 2428 5874 2440
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 5868 2400 6561 2428
rect 5868 2388 5874 2400
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 6638 2388 6644 2440
rect 6696 2428 6702 2440
rect 7300 2428 7328 2536
rect 16666 2524 16672 2576
rect 16724 2564 16730 2576
rect 20714 2564 20720 2576
rect 16724 2536 20720 2564
rect 16724 2524 16730 2536
rect 20714 2524 20720 2536
rect 20772 2524 20778 2576
rect 23569 2567 23627 2573
rect 23569 2533 23581 2567
rect 23615 2533 23627 2567
rect 23569 2527 23627 2533
rect 19978 2496 19984 2508
rect 6696 2400 7328 2428
rect 7392 2468 19984 2496
rect 6696 2388 6702 2400
rect 7392 2360 7420 2468
rect 19978 2456 19984 2468
rect 20036 2456 20042 2508
rect 23584 2496 23612 2527
rect 22388 2468 23612 2496
rect 7742 2428 7748 2440
rect 7703 2400 7748 2428
rect 7742 2388 7748 2400
rect 7800 2388 7806 2440
rect 9125 2431 9183 2437
rect 9125 2397 9137 2431
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 10413 2431 10471 2437
rect 10413 2397 10425 2431
rect 10459 2428 10471 2431
rect 10778 2428 10784 2440
rect 10459 2400 10784 2428
rect 10459 2397 10471 2400
rect 10413 2391 10471 2397
rect 9140 2360 9168 2391
rect 10778 2388 10784 2400
rect 10836 2388 10842 2440
rect 11606 2388 11612 2440
rect 11664 2428 11670 2440
rect 11885 2431 11943 2437
rect 11885 2428 11897 2431
rect 11664 2400 11897 2428
rect 11664 2388 11670 2400
rect 11885 2397 11897 2400
rect 11931 2397 11943 2431
rect 11885 2391 11943 2397
rect 13538 2388 13544 2440
rect 13596 2428 13602 2440
rect 14461 2431 14519 2437
rect 14461 2428 14473 2431
rect 13596 2400 14473 2428
rect 13596 2388 13602 2400
rect 14461 2397 14473 2400
rect 14507 2397 14519 2431
rect 14461 2391 14519 2397
rect 14826 2388 14832 2440
rect 14884 2428 14890 2440
rect 15105 2431 15163 2437
rect 15105 2428 15117 2431
rect 14884 2400 15117 2428
rect 14884 2388 14890 2400
rect 15105 2397 15117 2400
rect 15151 2397 15163 2431
rect 15105 2391 15163 2397
rect 16758 2388 16764 2440
rect 16816 2428 16822 2440
rect 17037 2431 17095 2437
rect 17037 2428 17049 2431
rect 16816 2400 17049 2428
rect 16816 2388 16822 2400
rect 17037 2397 17049 2400
rect 17083 2397 17095 2431
rect 18138 2428 18144 2440
rect 18099 2400 18144 2428
rect 17037 2391 17095 2397
rect 18138 2388 18144 2400
rect 18196 2388 18202 2440
rect 19334 2388 19340 2440
rect 19392 2430 19398 2440
rect 19429 2431 19487 2437
rect 19429 2430 19441 2431
rect 19392 2402 19441 2430
rect 19392 2388 19398 2402
rect 19429 2397 19441 2402
rect 19475 2397 19487 2431
rect 19429 2391 19487 2397
rect 20162 2388 20168 2440
rect 20220 2428 20226 2440
rect 20220 2400 20265 2428
rect 20220 2388 20226 2400
rect 21266 2388 21272 2440
rect 21324 2428 21330 2440
rect 22388 2437 22416 2468
rect 21453 2431 21511 2437
rect 21453 2428 21465 2431
rect 21324 2400 21465 2428
rect 21324 2388 21330 2400
rect 21453 2397 21465 2400
rect 21499 2397 21511 2431
rect 21453 2391 21511 2397
rect 22373 2431 22431 2437
rect 22373 2397 22385 2431
rect 22419 2397 22431 2431
rect 22925 2431 22983 2437
rect 22925 2428 22937 2431
rect 22373 2391 22431 2397
rect 22480 2400 22937 2428
rect 22480 2360 22508 2400
rect 22925 2397 22937 2400
rect 22971 2397 22983 2431
rect 22925 2391 22983 2397
rect 23753 2431 23811 2437
rect 23753 2397 23765 2431
rect 23799 2397 23811 2431
rect 23753 2391 23811 2397
rect 24581 2431 24639 2437
rect 24581 2397 24593 2431
rect 24627 2428 24639 2431
rect 25406 2428 25412 2440
rect 24627 2400 25412 2428
rect 24627 2397 24639 2400
rect 24581 2391 24639 2397
rect 5474 2332 7420 2360
rect 7576 2332 9168 2360
rect 16868 2332 22508 2360
rect 4522 2292 4528 2304
rect 3436 2264 4528 2292
rect 1765 2255 1823 2261
rect 4522 2252 4528 2264
rect 4580 2252 4586 2304
rect 5810 2252 5816 2304
rect 5868 2292 5874 2304
rect 7576 2301 7604 2332
rect 6733 2295 6791 2301
rect 6733 2292 6745 2295
rect 5868 2264 6745 2292
rect 5868 2252 5874 2264
rect 6733 2261 6745 2264
rect 6779 2261 6791 2295
rect 6733 2255 6791 2261
rect 7561 2295 7619 2301
rect 7561 2261 7573 2295
rect 7607 2261 7619 2295
rect 7561 2255 7619 2261
rect 9030 2252 9036 2304
rect 9088 2292 9094 2304
rect 9309 2295 9367 2301
rect 9309 2292 9321 2295
rect 9088 2264 9321 2292
rect 9088 2252 9094 2264
rect 9309 2261 9321 2264
rect 9355 2261 9367 2295
rect 9309 2255 9367 2261
rect 10318 2252 10324 2304
rect 10376 2292 10382 2304
rect 10597 2295 10655 2301
rect 10597 2292 10609 2295
rect 10376 2264 10609 2292
rect 10376 2252 10382 2264
rect 10597 2261 10609 2264
rect 10643 2261 10655 2295
rect 11698 2292 11704 2304
rect 11659 2264 11704 2292
rect 10597 2255 10655 2261
rect 11698 2252 11704 2264
rect 11756 2252 11762 2304
rect 14921 2295 14979 2301
rect 14921 2261 14933 2295
rect 14967 2292 14979 2295
rect 16666 2292 16672 2304
rect 14967 2264 16672 2292
rect 14967 2261 14979 2264
rect 14921 2255 14979 2261
rect 16666 2252 16672 2264
rect 16724 2252 16730 2304
rect 16868 2301 16896 2332
rect 22554 2320 22560 2372
rect 22612 2360 22618 2372
rect 23768 2360 23796 2391
rect 25406 2388 25412 2400
rect 25464 2388 25470 2440
rect 26053 2431 26111 2437
rect 26053 2397 26065 2431
rect 26099 2397 26111 2431
rect 26053 2391 26111 2397
rect 22612 2332 23796 2360
rect 26068 2360 26096 2391
rect 26206 2360 26234 2604
rect 27893 2567 27951 2573
rect 27893 2533 27905 2567
rect 27939 2533 27951 2567
rect 28000 2564 28028 2604
rect 28074 2592 28080 2644
rect 28132 2632 28138 2644
rect 28537 2635 28595 2641
rect 28537 2632 28549 2635
rect 28132 2604 28549 2632
rect 28132 2592 28138 2604
rect 28537 2601 28549 2604
rect 28583 2601 28595 2635
rect 29730 2632 29736 2644
rect 29691 2604 29736 2632
rect 28537 2595 28595 2601
rect 29730 2592 29736 2604
rect 29788 2592 29794 2644
rect 30469 2635 30527 2641
rect 30469 2601 30481 2635
rect 30515 2632 30527 2635
rect 32490 2632 32496 2644
rect 30515 2604 32496 2632
rect 30515 2601 30527 2604
rect 30469 2595 30527 2601
rect 32490 2592 32496 2604
rect 32548 2592 32554 2644
rect 32858 2592 32864 2644
rect 32916 2632 32922 2644
rect 33686 2632 33692 2644
rect 32916 2604 33180 2632
rect 33647 2604 33692 2632
rect 32916 2592 32922 2604
rect 28000 2536 31340 2564
rect 27893 2527 27951 2533
rect 27157 2431 27215 2437
rect 27157 2397 27169 2431
rect 27203 2428 27215 2431
rect 27908 2428 27936 2527
rect 27203 2400 27936 2428
rect 28077 2431 28135 2437
rect 27203 2397 27215 2400
rect 27157 2391 27215 2397
rect 28077 2397 28089 2431
rect 28123 2397 28135 2431
rect 28718 2428 28724 2440
rect 28679 2400 28724 2428
rect 28077 2391 28135 2397
rect 26068 2332 26234 2360
rect 22612 2320 22618 2332
rect 27062 2320 27068 2372
rect 27120 2360 27126 2372
rect 28092 2360 28120 2391
rect 28718 2388 28724 2400
rect 28776 2388 28782 2440
rect 29914 2428 29920 2440
rect 29875 2400 29920 2428
rect 29914 2388 29920 2400
rect 29972 2388 29978 2440
rect 30374 2428 30380 2440
rect 30335 2400 30380 2428
rect 30374 2388 30380 2400
rect 30432 2388 30438 2440
rect 31205 2431 31263 2437
rect 31205 2397 31217 2431
rect 31251 2397 31263 2431
rect 31205 2391 31263 2397
rect 27120 2332 28120 2360
rect 27120 2320 27126 2332
rect 28994 2320 29000 2372
rect 29052 2360 29058 2372
rect 31220 2360 31248 2391
rect 29052 2332 31248 2360
rect 31312 2360 31340 2536
rect 31662 2524 31668 2576
rect 31720 2564 31726 2576
rect 33045 2567 33103 2573
rect 33045 2564 33057 2567
rect 31720 2536 33057 2564
rect 31720 2524 31726 2536
rect 33045 2533 33057 2536
rect 33091 2533 33103 2567
rect 33152 2564 33180 2604
rect 33686 2592 33692 2604
rect 33744 2592 33750 2644
rect 34885 2567 34943 2573
rect 34885 2564 34897 2567
rect 33152 2536 34897 2564
rect 33045 2527 33103 2533
rect 34885 2533 34897 2536
rect 34931 2533 34943 2567
rect 34885 2527 34943 2533
rect 31754 2456 31760 2508
rect 31812 2496 31818 2508
rect 31812 2468 33272 2496
rect 31812 2456 31818 2468
rect 32306 2428 32312 2440
rect 32267 2400 32312 2428
rect 32306 2388 32312 2400
rect 32364 2388 32370 2440
rect 33244 2437 33272 2468
rect 33318 2456 33324 2508
rect 33376 2496 33382 2508
rect 33376 2468 38056 2496
rect 33376 2456 33382 2468
rect 33229 2431 33287 2437
rect 33229 2397 33241 2431
rect 33275 2397 33287 2431
rect 33229 2391 33287 2397
rect 33502 2388 33508 2440
rect 33560 2428 33566 2440
rect 33873 2431 33931 2437
rect 33873 2428 33885 2431
rect 33560 2400 33885 2428
rect 33560 2388 33566 2400
rect 33873 2397 33885 2400
rect 33919 2397 33931 2431
rect 33873 2391 33931 2397
rect 34790 2388 34796 2440
rect 34848 2428 34854 2440
rect 35069 2431 35127 2437
rect 35069 2428 35081 2431
rect 34848 2400 35081 2428
rect 34848 2388 34854 2400
rect 35069 2397 35081 2400
rect 35115 2397 35127 2431
rect 35069 2391 35127 2397
rect 36078 2388 36084 2440
rect 36136 2428 36142 2440
rect 38028 2437 38056 2468
rect 36357 2431 36415 2437
rect 36357 2428 36369 2431
rect 36136 2400 36369 2428
rect 36136 2388 36142 2400
rect 36357 2397 36369 2400
rect 36403 2397 36415 2431
rect 36357 2391 36415 2397
rect 38013 2431 38071 2437
rect 38013 2397 38025 2431
rect 38059 2397 38071 2431
rect 38013 2391 38071 2397
rect 31312 2332 35894 2360
rect 29052 2320 29058 2332
rect 16853 2295 16911 2301
rect 16853 2261 16865 2295
rect 16899 2261 16911 2295
rect 16853 2255 16911 2261
rect 18046 2252 18052 2304
rect 18104 2292 18110 2304
rect 18325 2295 18383 2301
rect 18325 2292 18337 2295
rect 18104 2264 18337 2292
rect 18104 2252 18110 2264
rect 18325 2261 18337 2264
rect 18371 2261 18383 2295
rect 18325 2255 18383 2261
rect 19334 2252 19340 2304
rect 19392 2292 19398 2304
rect 19613 2295 19671 2301
rect 19613 2292 19625 2295
rect 19392 2264 19625 2292
rect 19392 2252 19398 2264
rect 19613 2261 19625 2264
rect 19659 2261 19671 2295
rect 19613 2255 19671 2261
rect 21174 2252 21180 2304
rect 21232 2292 21238 2304
rect 21269 2295 21327 2301
rect 21269 2292 21281 2295
rect 21232 2264 21281 2292
rect 21232 2252 21238 2264
rect 21269 2261 21281 2264
rect 21315 2261 21327 2295
rect 21269 2255 21327 2261
rect 23842 2252 23848 2304
rect 23900 2292 23906 2304
rect 24765 2295 24823 2301
rect 24765 2292 24777 2295
rect 23900 2264 24777 2292
rect 23900 2252 23906 2264
rect 24765 2261 24777 2264
rect 24811 2261 24823 2295
rect 24765 2255 24823 2261
rect 26142 2252 26148 2304
rect 26200 2292 26206 2304
rect 27341 2295 27399 2301
rect 27341 2292 27353 2295
rect 26200 2264 27353 2292
rect 26200 2252 26206 2264
rect 27341 2261 27353 2264
rect 27387 2261 27399 2295
rect 27341 2255 27399 2261
rect 27430 2252 27436 2304
rect 27488 2292 27494 2304
rect 31021 2295 31079 2301
rect 31021 2292 31033 2295
rect 27488 2264 31033 2292
rect 27488 2252 27494 2264
rect 31021 2261 31033 2264
rect 31067 2261 31079 2295
rect 31021 2255 31079 2261
rect 31570 2252 31576 2304
rect 31628 2292 31634 2304
rect 32493 2295 32551 2301
rect 32493 2292 32505 2295
rect 31628 2264 32505 2292
rect 31628 2252 31634 2264
rect 32493 2261 32505 2264
rect 32539 2261 32551 2295
rect 35866 2292 35894 2332
rect 36173 2295 36231 2301
rect 36173 2292 36185 2295
rect 35866 2264 36185 2292
rect 32493 2255 32551 2261
rect 36173 2261 36185 2264
rect 36219 2261 36231 2295
rect 36173 2255 36231 2261
rect 38010 2252 38016 2304
rect 38068 2292 38074 2304
rect 38197 2295 38255 2301
rect 38197 2292 38209 2295
rect 38068 2264 38209 2292
rect 38068 2252 38074 2264
rect 38197 2261 38209 2264
rect 38243 2261 38255 2295
rect 38197 2255 38255 2261
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 7006 2048 7012 2100
rect 7064 2088 7070 2100
rect 11974 2088 11980 2100
rect 7064 2060 11980 2088
rect 7064 2048 7070 2060
rect 11974 2048 11980 2060
rect 12032 2048 12038 2100
rect 17954 2048 17960 2100
rect 18012 2088 18018 2100
rect 22830 2088 22836 2100
rect 18012 2060 22836 2088
rect 18012 2048 18018 2060
rect 22830 2048 22836 2060
rect 22888 2048 22894 2100
rect 11698 1980 11704 2032
rect 11756 2020 11762 2032
rect 26418 2020 26424 2032
rect 11756 1992 26424 2020
rect 11756 1980 11762 1992
rect 26418 1980 26424 1992
rect 26476 1980 26482 2032
rect 7742 1912 7748 1964
rect 7800 1952 7806 1964
rect 23934 1952 23940 1964
rect 7800 1924 23940 1952
rect 7800 1912 7806 1924
rect 23934 1912 23940 1924
rect 23992 1912 23998 1964
rect 19242 1844 19248 1896
rect 19300 1884 19306 1896
rect 21174 1884 21180 1896
rect 19300 1856 21180 1884
rect 19300 1844 19306 1856
rect 21174 1844 21180 1856
rect 21232 1844 21238 1896
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 37464 37315 37516 37324
rect 2780 37204 2832 37256
rect 3148 37247 3200 37256
rect 3148 37213 3157 37247
rect 3157 37213 3191 37247
rect 3191 37213 3200 37247
rect 3148 37204 3200 37213
rect 3240 37204 3292 37256
rect 4620 37204 4672 37256
rect 7840 37247 7892 37256
rect 4068 37136 4120 37188
rect 7840 37213 7849 37247
rect 7849 37213 7883 37247
rect 7883 37213 7892 37247
rect 7840 37204 7892 37213
rect 9036 37204 9088 37256
rect 37464 37281 37473 37315
rect 37473 37281 37507 37315
rect 37507 37281 37516 37315
rect 37464 37272 37516 37281
rect 11244 37204 11296 37256
rect 11704 37204 11756 37256
rect 13544 37204 13596 37256
rect 15568 37247 15620 37256
rect 15568 37213 15577 37247
rect 15577 37213 15611 37247
rect 15611 37213 15620 37247
rect 15568 37204 15620 37213
rect 16856 37247 16908 37256
rect 16856 37213 16865 37247
rect 16865 37213 16899 37247
rect 16899 37213 16908 37247
rect 16856 37204 16908 37213
rect 18052 37204 18104 37256
rect 22008 37247 22060 37256
rect 13728 37136 13780 37188
rect 17500 37136 17552 37188
rect 22008 37213 22017 37247
rect 22017 37213 22051 37247
rect 22051 37213 22060 37247
rect 22008 37204 22060 37213
rect 22560 37204 22612 37256
rect 24492 37204 24544 37256
rect 25780 37204 25832 37256
rect 27804 37247 27856 37256
rect 27804 37213 27813 37247
rect 27813 37213 27847 37247
rect 27847 37213 27856 37247
rect 27804 37204 27856 37213
rect 28632 37204 28684 37256
rect 30380 37204 30432 37256
rect 32220 37204 32272 37256
rect 33508 37204 33560 37256
rect 33876 37204 33928 37256
rect 28908 37136 28960 37188
rect 1308 37068 1360 37120
rect 2320 37111 2372 37120
rect 2320 37077 2329 37111
rect 2329 37077 2363 37111
rect 2363 37077 2372 37111
rect 2320 37068 2372 37077
rect 2964 37111 3016 37120
rect 2964 37077 2973 37111
rect 2973 37077 3007 37111
rect 3007 37077 3016 37111
rect 2964 37068 3016 37077
rect 3976 37111 4028 37120
rect 3976 37077 3985 37111
rect 3985 37077 4019 37111
rect 4019 37077 4028 37111
rect 3976 37068 4028 37077
rect 4620 37111 4672 37120
rect 4620 37077 4629 37111
rect 4629 37077 4663 37111
rect 4663 37077 4672 37111
rect 4620 37068 4672 37077
rect 5816 37068 5868 37120
rect 7748 37068 7800 37120
rect 8944 37068 8996 37120
rect 10324 37068 10376 37120
rect 12440 37068 12492 37120
rect 14280 37111 14332 37120
rect 14280 37077 14289 37111
rect 14289 37077 14323 37111
rect 14323 37077 14332 37111
rect 14280 37068 14332 37077
rect 15476 37068 15528 37120
rect 16764 37068 16816 37120
rect 17960 37068 18012 37120
rect 19984 37068 20036 37120
rect 21272 37068 21324 37120
rect 22744 37111 22796 37120
rect 22744 37077 22753 37111
rect 22753 37077 22787 37111
rect 22787 37077 22796 37111
rect 22744 37068 22796 37077
rect 23112 37068 23164 37120
rect 25136 37068 25188 37120
rect 27712 37068 27764 37120
rect 29000 37068 29052 37120
rect 32128 37136 32180 37188
rect 37740 37247 37792 37256
rect 37740 37213 37749 37247
rect 37749 37213 37783 37247
rect 37783 37213 37792 37247
rect 37740 37204 37792 37213
rect 32404 37068 32456 37120
rect 33324 37068 33376 37120
rect 34796 37068 34848 37120
rect 36728 37068 36780 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 20 36864 72 36916
rect 4620 36864 4672 36916
rect 10692 36864 10744 36916
rect 15568 36864 15620 36916
rect 18052 36864 18104 36916
rect 39304 36864 39356 36916
rect 2320 36796 2372 36848
rect 7656 36796 7708 36848
rect 4620 36728 4672 36780
rect 36912 36771 36964 36780
rect 36912 36737 36921 36771
rect 36921 36737 36955 36771
rect 36955 36737 36964 36771
rect 36912 36728 36964 36737
rect 37004 36728 37056 36780
rect 36728 36567 36780 36576
rect 36728 36533 36737 36567
rect 36737 36533 36771 36567
rect 36771 36533 36780 36567
rect 36728 36524 36780 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 38016 36116 38068 36168
rect 37280 35980 37332 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 4068 35232 4120 35284
rect 14096 35028 14148 35080
rect 33416 35028 33468 35080
rect 38200 34935 38252 34944
rect 38200 34901 38209 34935
rect 38209 34901 38243 34935
rect 38243 34901 38252 34935
rect 38200 34892 38252 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 32128 34688 32180 34740
rect 33876 34688 33928 34740
rect 31668 34595 31720 34604
rect 31668 34561 31677 34595
rect 31677 34561 31711 34595
rect 31711 34561 31720 34595
rect 31668 34552 31720 34561
rect 28540 34484 28592 34536
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 1768 33507 1820 33516
rect 1768 33473 1777 33507
rect 1777 33473 1811 33507
rect 1811 33473 1820 33507
rect 1768 33464 1820 33473
rect 38292 33507 38344 33516
rect 38292 33473 38301 33507
rect 38301 33473 38335 33507
rect 38335 33473 38344 33507
rect 38292 33464 38344 33473
rect 7196 33260 7248 33312
rect 38108 33303 38160 33312
rect 38108 33269 38117 33303
rect 38117 33269 38151 33303
rect 38151 33269 38160 33303
rect 38108 33260 38160 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 11244 33056 11296 33108
rect 31668 33056 31720 33108
rect 37004 33056 37056 33108
rect 12532 32852 12584 32904
rect 31116 32895 31168 32904
rect 31116 32861 31125 32895
rect 31125 32861 31159 32895
rect 31159 32861 31168 32895
rect 31116 32852 31168 32861
rect 32956 32895 33008 32904
rect 32956 32861 32965 32895
rect 32965 32861 32999 32895
rect 32999 32861 33008 32895
rect 32956 32852 33008 32861
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 4620 32512 4672 32564
rect 11704 32555 11756 32564
rect 11704 32521 11713 32555
rect 11713 32521 11747 32555
rect 11747 32521 11756 32555
rect 11704 32512 11756 32521
rect 17500 32555 17552 32564
rect 17500 32521 17509 32555
rect 17509 32521 17543 32555
rect 17543 32521 17552 32555
rect 17500 32512 17552 32521
rect 28632 32555 28684 32564
rect 28632 32521 28641 32555
rect 28641 32521 28675 32555
rect 28675 32521 28684 32555
rect 28632 32512 28684 32521
rect 1768 32419 1820 32428
rect 1768 32385 1777 32419
rect 1777 32385 1811 32419
rect 1811 32385 1820 32419
rect 1768 32376 1820 32385
rect 4620 32376 4672 32428
rect 11888 32419 11940 32428
rect 11888 32385 11897 32419
rect 11897 32385 11931 32419
rect 11931 32385 11940 32419
rect 11888 32376 11940 32385
rect 16948 32376 17000 32428
rect 28816 32419 28868 32428
rect 28816 32385 28825 32419
rect 28825 32385 28859 32419
rect 28859 32385 28868 32419
rect 28816 32376 28868 32385
rect 35440 32376 35492 32428
rect 6276 32172 6328 32224
rect 38200 32215 38252 32224
rect 38200 32181 38209 32215
rect 38209 32181 38243 32215
rect 38243 32181 38252 32215
rect 38200 32172 38252 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 7840 31968 7892 32020
rect 16856 32011 16908 32020
rect 16856 31977 16865 32011
rect 16865 31977 16899 32011
rect 16899 31977 16908 32011
rect 16856 31968 16908 31977
rect 14280 31900 14332 31952
rect 10600 31764 10652 31816
rect 17040 31807 17092 31816
rect 17040 31773 17049 31807
rect 17049 31773 17083 31807
rect 17083 31773 17092 31807
rect 17040 31764 17092 31773
rect 27528 31832 27580 31884
rect 36728 31764 36780 31816
rect 26792 31671 26844 31680
rect 26792 31637 26801 31671
rect 26801 31637 26835 31671
rect 26835 31637 26844 31671
rect 26792 31628 26844 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 27804 31424 27856 31476
rect 15568 31288 15620 31340
rect 19432 31288 19484 31340
rect 26148 31331 26200 31340
rect 26148 31297 26157 31331
rect 26157 31297 26191 31331
rect 26191 31297 26200 31331
rect 26148 31288 26200 31297
rect 37280 31288 37332 31340
rect 19524 31220 19576 31272
rect 15292 31084 15344 31136
rect 19708 31084 19760 31136
rect 30472 31127 30524 31136
rect 30472 31093 30481 31127
rect 30481 31093 30515 31127
rect 30515 31093 30524 31127
rect 30472 31084 30524 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 13728 30880 13780 30932
rect 17040 30880 17092 30932
rect 18052 30923 18104 30932
rect 18052 30889 18061 30923
rect 18061 30889 18095 30923
rect 18095 30889 18104 30923
rect 18052 30880 18104 30889
rect 19524 30787 19576 30796
rect 19524 30753 19533 30787
rect 19533 30753 19567 30787
rect 19567 30753 19576 30787
rect 19524 30744 19576 30753
rect 19708 30787 19760 30796
rect 19708 30753 19717 30787
rect 19717 30753 19751 30787
rect 19751 30753 19760 30787
rect 19708 30744 19760 30753
rect 27528 30744 27580 30796
rect 1584 30719 1636 30728
rect 1584 30685 1593 30719
rect 1593 30685 1627 30719
rect 1627 30685 1636 30719
rect 1584 30676 1636 30685
rect 1860 30719 1912 30728
rect 1860 30685 1869 30719
rect 1869 30685 1903 30719
rect 1903 30685 1912 30719
rect 1860 30676 1912 30685
rect 11244 30719 11296 30728
rect 11244 30685 11253 30719
rect 11253 30685 11287 30719
rect 11287 30685 11296 30719
rect 11244 30676 11296 30685
rect 14464 30719 14516 30728
rect 14464 30685 14473 30719
rect 14473 30685 14507 30719
rect 14507 30685 14516 30719
rect 14464 30676 14516 30685
rect 19984 30676 20036 30728
rect 22560 30719 22612 30728
rect 22560 30685 22569 30719
rect 22569 30685 22603 30719
rect 22603 30685 22612 30719
rect 22560 30676 22612 30685
rect 33324 30719 33376 30728
rect 33324 30685 33333 30719
rect 33333 30685 33367 30719
rect 33367 30685 33376 30719
rect 33324 30676 33376 30685
rect 18880 30608 18932 30660
rect 11980 30540 12032 30592
rect 20168 30583 20220 30592
rect 20168 30549 20177 30583
rect 20177 30549 20211 30583
rect 20211 30549 20220 30583
rect 20168 30540 20220 30549
rect 24032 30608 24084 30660
rect 31760 30540 31812 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 14464 30336 14516 30388
rect 19432 30336 19484 30388
rect 10600 30311 10652 30320
rect 10600 30277 10609 30311
rect 10609 30277 10643 30311
rect 10643 30277 10652 30311
rect 10600 30268 10652 30277
rect 12532 30311 12584 30320
rect 12532 30277 12541 30311
rect 12541 30277 12575 30311
rect 12575 30277 12584 30311
rect 12532 30268 12584 30277
rect 14096 30268 14148 30320
rect 16948 30311 17000 30320
rect 16948 30277 16957 30311
rect 16957 30277 16991 30311
rect 16991 30277 17000 30311
rect 16948 30268 17000 30277
rect 12256 30200 12308 30252
rect 12440 30243 12492 30252
rect 12440 30209 12449 30243
rect 12449 30209 12483 30243
rect 12483 30209 12492 30243
rect 14188 30243 14240 30252
rect 12440 30200 12492 30209
rect 14188 30209 14197 30243
rect 14197 30209 14231 30243
rect 14231 30209 14240 30243
rect 14188 30200 14240 30209
rect 15016 30200 15068 30252
rect 16856 30243 16908 30252
rect 16856 30209 16865 30243
rect 16865 30209 16899 30243
rect 16899 30209 16908 30243
rect 16856 30200 16908 30209
rect 19248 30200 19300 30252
rect 22560 30336 22612 30388
rect 24952 30336 25004 30388
rect 32956 30268 33008 30320
rect 23112 30243 23164 30252
rect 23112 30209 23121 30243
rect 23121 30209 23155 30243
rect 23155 30209 23164 30243
rect 23112 30200 23164 30209
rect 24768 30200 24820 30252
rect 33600 30243 33652 30252
rect 33600 30209 33609 30243
rect 33609 30209 33643 30243
rect 33643 30209 33652 30243
rect 33600 30200 33652 30209
rect 5172 30132 5224 30184
rect 7288 30175 7340 30184
rect 7288 30141 7297 30175
rect 7297 30141 7331 30175
rect 7331 30141 7340 30175
rect 7288 30132 7340 30141
rect 33324 30132 33376 30184
rect 33416 30107 33468 30116
rect 33416 30073 33425 30107
rect 33425 30073 33459 30107
rect 33459 30073 33468 30107
rect 33416 30064 33468 30073
rect 8668 29996 8720 30048
rect 23204 30039 23256 30048
rect 23204 30005 23213 30039
rect 23213 30005 23247 30039
rect 23247 30005 23256 30039
rect 23204 29996 23256 30005
rect 38200 30039 38252 30048
rect 38200 30005 38209 30039
rect 38209 30005 38243 30039
rect 38243 30005 38252 30039
rect 38200 29996 38252 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 5172 29835 5224 29844
rect 5172 29801 5181 29835
rect 5181 29801 5215 29835
rect 5215 29801 5224 29835
rect 5172 29792 5224 29801
rect 7288 29835 7340 29844
rect 7288 29801 7297 29835
rect 7297 29801 7331 29835
rect 7331 29801 7340 29835
rect 7288 29792 7340 29801
rect 11888 29792 11940 29844
rect 14188 29792 14240 29844
rect 15108 29792 15160 29844
rect 26148 29792 26200 29844
rect 28816 29792 28868 29844
rect 16856 29724 16908 29776
rect 15292 29656 15344 29708
rect 20168 29724 20220 29776
rect 2964 29588 3016 29640
rect 8484 29588 8536 29640
rect 10784 29588 10836 29640
rect 30472 29656 30524 29708
rect 15568 29588 15620 29640
rect 19340 29588 19392 29640
rect 21088 29631 21140 29640
rect 21088 29597 21097 29631
rect 21097 29597 21131 29631
rect 21131 29597 21140 29631
rect 21088 29588 21140 29597
rect 8668 29520 8720 29572
rect 10140 29563 10192 29572
rect 10140 29529 10149 29563
rect 10149 29529 10183 29563
rect 10183 29529 10192 29563
rect 11888 29563 11940 29572
rect 10140 29520 10192 29529
rect 11888 29529 11897 29563
rect 11897 29529 11931 29563
rect 11931 29529 11940 29563
rect 11888 29520 11940 29529
rect 11980 29563 12032 29572
rect 11980 29529 11989 29563
rect 11989 29529 12023 29563
rect 12023 29529 12032 29563
rect 18144 29563 18196 29572
rect 11980 29520 12032 29529
rect 18144 29529 18153 29563
rect 18153 29529 18187 29563
rect 18187 29529 18196 29563
rect 18144 29520 18196 29529
rect 18236 29563 18288 29572
rect 18236 29529 18245 29563
rect 18245 29529 18279 29563
rect 18279 29529 18288 29563
rect 18236 29520 18288 29529
rect 18880 29520 18932 29572
rect 26240 29588 26292 29640
rect 15844 29495 15896 29504
rect 15844 29461 15853 29495
rect 15853 29461 15887 29495
rect 15887 29461 15896 29495
rect 15844 29452 15896 29461
rect 16580 29452 16632 29504
rect 20996 29452 21048 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 8668 29291 8720 29300
rect 8668 29257 8677 29291
rect 8677 29257 8711 29291
rect 8711 29257 8720 29291
rect 8668 29248 8720 29257
rect 10140 29248 10192 29300
rect 11888 29291 11940 29300
rect 11888 29257 11897 29291
rect 11897 29257 11931 29291
rect 11931 29257 11940 29291
rect 11888 29248 11940 29257
rect 15108 29291 15160 29300
rect 15108 29257 15117 29291
rect 15117 29257 15151 29291
rect 15151 29257 15160 29291
rect 15108 29248 15160 29257
rect 18144 29291 18196 29300
rect 18144 29257 18153 29291
rect 18153 29257 18187 29291
rect 18187 29257 18196 29291
rect 18144 29248 18196 29257
rect 19340 29291 19392 29300
rect 19340 29257 19349 29291
rect 19349 29257 19383 29291
rect 19383 29257 19392 29291
rect 19340 29248 19392 29257
rect 19984 29291 20036 29300
rect 19984 29257 19993 29291
rect 19993 29257 20027 29291
rect 20027 29257 20036 29291
rect 19984 29248 20036 29257
rect 22008 29248 22060 29300
rect 1768 29155 1820 29164
rect 1768 29121 1777 29155
rect 1777 29121 1811 29155
rect 1811 29121 1820 29155
rect 1768 29112 1820 29121
rect 11244 29112 11296 29164
rect 24032 29180 24084 29232
rect 15844 29112 15896 29164
rect 19248 29155 19300 29164
rect 19248 29121 19257 29155
rect 19257 29121 19291 29155
rect 19291 29121 19300 29155
rect 19248 29112 19300 29121
rect 20168 29112 20220 29164
rect 20996 29155 21048 29164
rect 20996 29121 21005 29155
rect 21005 29121 21039 29155
rect 21039 29121 21048 29155
rect 20996 29112 21048 29121
rect 38292 29155 38344 29164
rect 38292 29121 38301 29155
rect 38301 29121 38335 29155
rect 38335 29121 38344 29155
rect 38292 29112 38344 29121
rect 8024 29087 8076 29096
rect 8024 29053 8033 29087
rect 8033 29053 8067 29087
rect 8067 29053 8076 29087
rect 8024 29044 8076 29053
rect 8208 29087 8260 29096
rect 8208 29053 8217 29087
rect 8217 29053 8251 29087
rect 8251 29053 8260 29087
rect 8208 29044 8260 29053
rect 5724 28976 5776 29028
rect 34520 28976 34572 29028
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 12440 28704 12492 28756
rect 13268 28704 13320 28756
rect 13452 28704 13504 28756
rect 22100 28704 22152 28756
rect 33600 28704 33652 28756
rect 8024 28636 8076 28688
rect 14740 28636 14792 28688
rect 14004 28568 14056 28620
rect 7656 28543 7708 28552
rect 7656 28509 7665 28543
rect 7665 28509 7699 28543
rect 7699 28509 7708 28543
rect 7656 28500 7708 28509
rect 8484 28543 8536 28552
rect 8484 28509 8493 28543
rect 8493 28509 8527 28543
rect 8527 28509 8536 28543
rect 8484 28500 8536 28509
rect 10232 28543 10284 28552
rect 10232 28509 10241 28543
rect 10241 28509 10275 28543
rect 10275 28509 10284 28543
rect 10232 28500 10284 28509
rect 10692 28543 10744 28552
rect 10692 28509 10701 28543
rect 10701 28509 10735 28543
rect 10735 28509 10744 28543
rect 10692 28500 10744 28509
rect 12900 28543 12952 28552
rect 12900 28509 12909 28543
rect 12909 28509 12943 28543
rect 12943 28509 12952 28543
rect 12900 28500 12952 28509
rect 15292 28432 15344 28484
rect 8392 28364 8444 28416
rect 10048 28407 10100 28416
rect 10048 28373 10057 28407
rect 10057 28373 10091 28407
rect 10091 28373 10100 28407
rect 10048 28364 10100 28373
rect 11704 28364 11756 28416
rect 14464 28364 14516 28416
rect 15200 28407 15252 28416
rect 15200 28373 15209 28407
rect 15209 28373 15243 28407
rect 15243 28373 15252 28407
rect 15200 28364 15252 28373
rect 26424 28500 26476 28552
rect 34520 28500 34572 28552
rect 19984 28364 20036 28416
rect 29460 28364 29512 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 8208 28203 8260 28212
rect 8208 28169 8217 28203
rect 8217 28169 8251 28203
rect 8251 28169 8260 28203
rect 8208 28160 8260 28169
rect 12900 28160 12952 28212
rect 13268 28203 13320 28212
rect 13268 28169 13277 28203
rect 13277 28169 13311 28203
rect 13311 28169 13320 28203
rect 13268 28160 13320 28169
rect 14464 28135 14516 28144
rect 14464 28101 14473 28135
rect 14473 28101 14507 28135
rect 14507 28101 14516 28135
rect 14464 28092 14516 28101
rect 16120 28092 16172 28144
rect 19984 28160 20036 28212
rect 28540 28203 28592 28212
rect 20076 28092 20128 28144
rect 20904 28135 20956 28144
rect 20904 28101 20913 28135
rect 20913 28101 20947 28135
rect 20947 28101 20956 28135
rect 20904 28092 20956 28101
rect 21916 28092 21968 28144
rect 28540 28169 28549 28203
rect 28549 28169 28583 28203
rect 28583 28169 28592 28203
rect 28540 28160 28592 28169
rect 35440 28203 35492 28212
rect 35440 28169 35449 28203
rect 35449 28169 35483 28203
rect 35483 28169 35492 28203
rect 35440 28160 35492 28169
rect 3976 28024 4028 28076
rect 8392 28067 8444 28076
rect 8392 28033 8401 28067
rect 8401 28033 8435 28067
rect 8435 28033 8444 28067
rect 8392 28024 8444 28033
rect 8944 28067 8996 28076
rect 8944 28033 8953 28067
rect 8953 28033 8987 28067
rect 8987 28033 8996 28067
rect 8944 28024 8996 28033
rect 10048 28067 10100 28076
rect 10048 28033 10057 28067
rect 10057 28033 10091 28067
rect 10091 28033 10100 28067
rect 10048 28024 10100 28033
rect 14004 28024 14056 28076
rect 22744 28024 22796 28076
rect 27804 28092 27856 28144
rect 27988 28067 28040 28076
rect 9864 27999 9916 28008
rect 9864 27965 9873 27999
rect 9873 27965 9907 27999
rect 9907 27965 9916 27999
rect 9864 27956 9916 27965
rect 12624 27999 12676 28008
rect 12624 27965 12633 27999
rect 12633 27965 12667 27999
rect 12667 27965 12676 27999
rect 12624 27956 12676 27965
rect 15200 27956 15252 28008
rect 15292 27956 15344 28008
rect 15108 27888 15160 27940
rect 20168 27931 20220 27940
rect 20168 27897 20177 27931
rect 20177 27897 20211 27931
rect 20211 27897 20220 27931
rect 20168 27888 20220 27897
rect 23204 27956 23256 28008
rect 20628 27888 20680 27940
rect 22100 27931 22152 27940
rect 22100 27897 22109 27931
rect 22109 27897 22143 27931
rect 22143 27897 22152 27931
rect 22100 27888 22152 27897
rect 27988 28033 27997 28067
rect 27997 28033 28031 28067
rect 28031 28033 28040 28067
rect 27988 28024 28040 28033
rect 29460 28067 29512 28076
rect 29460 28033 29469 28067
rect 29469 28033 29503 28067
rect 29503 28033 29512 28067
rect 29460 28024 29512 28033
rect 33140 28024 33192 28076
rect 29644 27999 29696 28008
rect 29644 27965 29653 27999
rect 29653 27965 29687 27999
rect 29687 27965 29696 27999
rect 29644 27956 29696 27965
rect 6828 27820 6880 27872
rect 10508 27863 10560 27872
rect 10508 27829 10517 27863
rect 10517 27829 10551 27863
rect 10551 27829 10560 27863
rect 10508 27820 10560 27829
rect 27160 27863 27212 27872
rect 27160 27829 27169 27863
rect 27169 27829 27203 27863
rect 27203 27829 27212 27863
rect 27160 27820 27212 27829
rect 27252 27820 27304 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 5908 27616 5960 27668
rect 6828 27616 6880 27668
rect 9864 27616 9916 27668
rect 19432 27616 19484 27668
rect 29644 27616 29696 27668
rect 1768 27455 1820 27464
rect 1768 27421 1777 27455
rect 1777 27421 1811 27455
rect 1811 27421 1820 27455
rect 1768 27412 1820 27421
rect 5724 27455 5776 27464
rect 5724 27421 5733 27455
rect 5733 27421 5767 27455
rect 5767 27421 5776 27455
rect 5724 27412 5776 27421
rect 6736 27455 6788 27464
rect 6736 27421 6745 27455
rect 6745 27421 6779 27455
rect 6779 27421 6788 27455
rect 6736 27412 6788 27421
rect 7196 27455 7248 27464
rect 7196 27421 7205 27455
rect 7205 27421 7239 27455
rect 7239 27421 7248 27455
rect 7196 27412 7248 27421
rect 8944 27344 8996 27396
rect 5356 27276 5408 27328
rect 5816 27319 5868 27328
rect 5816 27285 5825 27319
rect 5825 27285 5859 27319
rect 5859 27285 5868 27319
rect 5816 27276 5868 27285
rect 7840 27319 7892 27328
rect 7840 27285 7849 27319
rect 7849 27285 7883 27319
rect 7883 27285 7892 27319
rect 7840 27276 7892 27285
rect 9128 27319 9180 27328
rect 9128 27285 9137 27319
rect 9137 27285 9171 27319
rect 9171 27285 9180 27319
rect 9128 27276 9180 27285
rect 10508 27548 10560 27600
rect 26792 27548 26844 27600
rect 11520 27480 11572 27532
rect 12624 27480 12676 27532
rect 27252 27480 27304 27532
rect 27988 27480 28040 27532
rect 33140 27548 33192 27600
rect 10324 27455 10376 27464
rect 10324 27421 10333 27455
rect 10333 27421 10367 27455
rect 10367 27421 10376 27455
rect 10784 27455 10836 27464
rect 10324 27412 10376 27421
rect 10784 27421 10793 27455
rect 10793 27421 10827 27455
rect 10827 27421 10836 27455
rect 10784 27412 10836 27421
rect 11428 27455 11480 27464
rect 11428 27421 11437 27455
rect 11437 27421 11471 27455
rect 11471 27421 11480 27455
rect 11428 27412 11480 27421
rect 16764 27455 16816 27464
rect 16764 27421 16773 27455
rect 16773 27421 16807 27455
rect 16807 27421 16816 27455
rect 16764 27412 16816 27421
rect 26608 27455 26660 27464
rect 26608 27421 26617 27455
rect 26617 27421 26651 27455
rect 26651 27421 26660 27455
rect 26608 27412 26660 27421
rect 28908 27412 28960 27464
rect 17500 27387 17552 27396
rect 17500 27353 17509 27387
rect 17509 27353 17543 27387
rect 17543 27353 17552 27387
rect 17500 27344 17552 27353
rect 18144 27387 18196 27396
rect 13268 27276 13320 27328
rect 18144 27353 18153 27387
rect 18153 27353 18187 27387
rect 18187 27353 18196 27387
rect 18144 27344 18196 27353
rect 23848 27344 23900 27396
rect 27804 27276 27856 27328
rect 28264 27276 28316 27328
rect 38200 27319 38252 27328
rect 38200 27285 38209 27319
rect 38209 27285 38243 27319
rect 38243 27285 38252 27319
rect 38200 27276 38252 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 11428 27072 11480 27124
rect 6736 27004 6788 27056
rect 5816 26936 5868 26988
rect 9128 26979 9180 26988
rect 9128 26945 9137 26979
rect 9137 26945 9171 26979
rect 9171 26945 9180 26979
rect 9128 26936 9180 26945
rect 10324 27004 10376 27056
rect 17500 27072 17552 27124
rect 18236 27072 18288 27124
rect 13268 27047 13320 27056
rect 13268 27013 13277 27047
rect 13277 27013 13311 27047
rect 13311 27013 13320 27047
rect 13268 27004 13320 27013
rect 13544 27004 13596 27056
rect 16764 27004 16816 27056
rect 26608 27072 26660 27124
rect 11520 26936 11572 26988
rect 14740 26979 14792 26988
rect 14740 26945 14749 26979
rect 14749 26945 14783 26979
rect 14783 26945 14792 26979
rect 14740 26936 14792 26945
rect 17592 26936 17644 26988
rect 17960 26979 18012 26988
rect 17960 26945 17969 26979
rect 17969 26945 18003 26979
rect 18003 26945 18012 26979
rect 17960 26936 18012 26945
rect 19340 26979 19392 26988
rect 19340 26945 19349 26979
rect 19349 26945 19383 26979
rect 19383 26945 19392 26979
rect 19340 26936 19392 26945
rect 21180 26979 21232 26988
rect 21180 26945 21189 26979
rect 21189 26945 21223 26979
rect 21223 26945 21232 26979
rect 21180 26936 21232 26945
rect 25136 26979 25188 26988
rect 8300 26868 8352 26920
rect 14924 26911 14976 26920
rect 14924 26877 14933 26911
rect 14933 26877 14967 26911
rect 14967 26877 14976 26911
rect 14924 26868 14976 26877
rect 16488 26868 16540 26920
rect 18696 26868 18748 26920
rect 25136 26945 25145 26979
rect 25145 26945 25179 26979
rect 25179 26945 25188 26979
rect 25136 26936 25188 26945
rect 25320 26936 25372 26988
rect 32404 26979 32456 26988
rect 32404 26945 32413 26979
rect 32413 26945 32447 26979
rect 32447 26945 32456 26979
rect 32404 26936 32456 26945
rect 25964 26868 26016 26920
rect 10232 26800 10284 26852
rect 20812 26800 20864 26852
rect 24308 26800 24360 26852
rect 7748 26775 7800 26784
rect 7748 26741 7757 26775
rect 7757 26741 7791 26775
rect 7791 26741 7800 26775
rect 7748 26732 7800 26741
rect 9312 26732 9364 26784
rect 15384 26775 15436 26784
rect 15384 26741 15393 26775
rect 15393 26741 15427 26775
rect 15427 26741 15436 26775
rect 15384 26732 15436 26741
rect 16672 26732 16724 26784
rect 20996 26775 21048 26784
rect 20996 26741 21005 26775
rect 21005 26741 21039 26775
rect 21039 26741 21048 26775
rect 20996 26732 21048 26741
rect 23940 26775 23992 26784
rect 23940 26741 23949 26775
rect 23949 26741 23983 26775
rect 23983 26741 23992 26775
rect 23940 26732 23992 26741
rect 25044 26732 25096 26784
rect 31852 26732 31904 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 10784 26528 10836 26580
rect 12900 26528 12952 26580
rect 13544 26571 13596 26580
rect 13544 26537 13553 26571
rect 13553 26537 13587 26571
rect 13587 26537 13596 26571
rect 13544 26528 13596 26537
rect 14924 26528 14976 26580
rect 17592 26571 17644 26580
rect 17592 26537 17601 26571
rect 17601 26537 17635 26571
rect 17635 26537 17644 26571
rect 17592 26528 17644 26537
rect 20076 26528 20128 26580
rect 27804 26571 27856 26580
rect 27804 26537 27813 26571
rect 27813 26537 27847 26571
rect 27847 26537 27856 26571
rect 27804 26528 27856 26537
rect 7748 26392 7800 26444
rect 9312 26435 9364 26444
rect 9312 26401 9321 26435
rect 9321 26401 9355 26435
rect 9355 26401 9364 26435
rect 9312 26392 9364 26401
rect 15384 26460 15436 26512
rect 16488 26435 16540 26444
rect 16488 26401 16497 26435
rect 16497 26401 16531 26435
rect 16531 26401 16540 26435
rect 16488 26392 16540 26401
rect 16672 26435 16724 26444
rect 16672 26401 16681 26435
rect 16681 26401 16715 26435
rect 16715 26401 16724 26435
rect 16672 26392 16724 26401
rect 18144 26460 18196 26512
rect 24492 26460 24544 26512
rect 26332 26460 26384 26512
rect 24216 26392 24268 26444
rect 24768 26392 24820 26444
rect 25964 26435 26016 26444
rect 25964 26401 25973 26435
rect 25973 26401 26007 26435
rect 26007 26401 26016 26435
rect 25964 26392 26016 26401
rect 27160 26392 27212 26444
rect 13084 26324 13136 26376
rect 14372 26324 14424 26376
rect 14648 26324 14700 26376
rect 20352 26367 20404 26376
rect 20352 26333 20361 26367
rect 20361 26333 20395 26367
rect 20395 26333 20404 26367
rect 20352 26324 20404 26333
rect 25320 26324 25372 26376
rect 20996 26299 21048 26308
rect 20996 26265 21005 26299
rect 21005 26265 21039 26299
rect 21039 26265 21048 26299
rect 27528 26324 27580 26376
rect 37740 26324 37792 26376
rect 20996 26256 21048 26265
rect 27804 26256 27856 26308
rect 27896 26256 27948 26308
rect 7288 26231 7340 26240
rect 7288 26197 7297 26231
rect 7297 26197 7331 26231
rect 7331 26197 7340 26231
rect 7288 26188 7340 26197
rect 23020 26188 23072 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 7748 25984 7800 26036
rect 14372 26027 14424 26036
rect 14372 25993 14381 26027
rect 14381 25993 14415 26027
rect 14415 25993 14424 26027
rect 14372 25984 14424 25993
rect 8944 25959 8996 25968
rect 8944 25925 8953 25959
rect 8953 25925 8987 25959
rect 8987 25925 8996 25959
rect 8944 25916 8996 25925
rect 9772 25916 9824 25968
rect 7288 25891 7340 25900
rect 7288 25857 7297 25891
rect 7297 25857 7331 25891
rect 7331 25857 7340 25891
rect 7288 25848 7340 25857
rect 7840 25848 7892 25900
rect 11520 25848 11572 25900
rect 11704 25891 11756 25900
rect 11704 25857 11713 25891
rect 11713 25857 11747 25891
rect 11747 25857 11756 25891
rect 11704 25848 11756 25857
rect 13636 25891 13688 25900
rect 10968 25687 11020 25696
rect 10968 25653 10977 25687
rect 10977 25653 11011 25687
rect 11011 25653 11020 25687
rect 10968 25644 11020 25653
rect 12716 25780 12768 25832
rect 13360 25712 13412 25764
rect 13636 25857 13645 25891
rect 13645 25857 13679 25891
rect 13679 25857 13688 25891
rect 13636 25848 13688 25857
rect 14280 25848 14332 25900
rect 15476 25916 15528 25968
rect 19340 25984 19392 26036
rect 20352 25984 20404 26036
rect 21180 25984 21232 26036
rect 21272 25916 21324 25968
rect 23020 25959 23072 25968
rect 23020 25925 23029 25959
rect 23029 25925 23063 25959
rect 23063 25925 23072 25959
rect 23020 25916 23072 25925
rect 23940 25916 23992 25968
rect 16580 25848 16632 25900
rect 19340 25848 19392 25900
rect 20352 25891 20404 25900
rect 20352 25857 20361 25891
rect 20361 25857 20395 25891
rect 20395 25857 20404 25891
rect 20352 25848 20404 25857
rect 22836 25848 22888 25900
rect 24308 25959 24360 25968
rect 24308 25925 24317 25959
rect 24317 25925 24351 25959
rect 24351 25925 24360 25959
rect 24308 25916 24360 25925
rect 27528 25984 27580 26036
rect 27804 26027 27856 26036
rect 27804 25993 27813 26027
rect 27813 25993 27847 26027
rect 27847 25993 27856 26027
rect 27804 25984 27856 25993
rect 26424 25916 26476 25968
rect 26332 25891 26384 25900
rect 15200 25780 15252 25832
rect 16212 25780 16264 25832
rect 23480 25780 23532 25832
rect 26332 25857 26341 25891
rect 26341 25857 26375 25891
rect 26375 25857 26384 25891
rect 26332 25848 26384 25857
rect 27804 25848 27856 25900
rect 24492 25823 24544 25832
rect 24492 25789 24501 25823
rect 24501 25789 24535 25823
rect 24535 25789 24544 25823
rect 24492 25780 24544 25789
rect 27344 25823 27396 25832
rect 27344 25789 27353 25823
rect 27353 25789 27387 25823
rect 27387 25789 27396 25823
rect 27344 25780 27396 25789
rect 27712 25712 27764 25764
rect 28448 25712 28500 25764
rect 19984 25644 20036 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 8300 25483 8352 25492
rect 8300 25449 8309 25483
rect 8309 25449 8343 25483
rect 8343 25449 8352 25483
rect 8300 25440 8352 25449
rect 9772 25483 9824 25492
rect 9772 25449 9781 25483
rect 9781 25449 9815 25483
rect 9815 25449 9824 25483
rect 9772 25440 9824 25449
rect 11520 25483 11572 25492
rect 11520 25449 11529 25483
rect 11529 25449 11563 25483
rect 11563 25449 11572 25483
rect 11520 25440 11572 25449
rect 15200 25440 15252 25492
rect 15476 25483 15528 25492
rect 15476 25449 15485 25483
rect 15485 25449 15519 25483
rect 15519 25449 15528 25483
rect 15476 25440 15528 25449
rect 16120 25483 16172 25492
rect 16120 25449 16129 25483
rect 16129 25449 16163 25483
rect 16163 25449 16172 25483
rect 16120 25440 16172 25449
rect 12716 25347 12768 25356
rect 12716 25313 12725 25347
rect 12725 25313 12759 25347
rect 12759 25313 12768 25347
rect 12716 25304 12768 25313
rect 12900 25347 12952 25356
rect 12900 25313 12909 25347
rect 12909 25313 12943 25347
rect 12943 25313 12952 25347
rect 12900 25304 12952 25313
rect 23480 25372 23532 25424
rect 25044 25347 25096 25356
rect 1768 25279 1820 25288
rect 1768 25245 1777 25279
rect 1777 25245 1811 25279
rect 1811 25245 1820 25279
rect 1768 25236 1820 25245
rect 6184 25236 6236 25288
rect 6736 25236 6788 25288
rect 9956 25279 10008 25288
rect 9956 25245 9965 25279
rect 9965 25245 9999 25279
rect 9999 25245 10008 25279
rect 9956 25236 10008 25245
rect 11704 25279 11756 25288
rect 11704 25245 11713 25279
rect 11713 25245 11747 25279
rect 11747 25245 11756 25279
rect 11704 25236 11756 25245
rect 25044 25313 25053 25347
rect 25053 25313 25087 25347
rect 25087 25313 25096 25347
rect 25044 25304 25096 25313
rect 16764 25236 16816 25288
rect 16856 25236 16908 25288
rect 18420 25236 18472 25288
rect 18696 25279 18748 25288
rect 18696 25245 18705 25279
rect 18705 25245 18739 25279
rect 18739 25245 18748 25279
rect 18696 25236 18748 25245
rect 38108 25440 38160 25492
rect 28448 25415 28500 25424
rect 28448 25381 28457 25415
rect 28457 25381 28491 25415
rect 28491 25381 28500 25415
rect 32128 25415 32180 25424
rect 28448 25372 28500 25381
rect 32128 25381 32137 25415
rect 32137 25381 32171 25415
rect 32171 25381 32180 25415
rect 32128 25372 32180 25381
rect 31760 25347 31812 25356
rect 31760 25313 31769 25347
rect 31769 25313 31803 25347
rect 31803 25313 31812 25347
rect 31760 25304 31812 25313
rect 31944 25279 31996 25288
rect 31944 25245 31953 25279
rect 31953 25245 31987 25279
rect 31987 25245 31996 25279
rect 31944 25236 31996 25245
rect 38292 25279 38344 25288
rect 38292 25245 38301 25279
rect 38301 25245 38335 25279
rect 38335 25245 38344 25279
rect 38292 25236 38344 25245
rect 13360 25168 13412 25220
rect 17868 25168 17920 25220
rect 3148 25100 3200 25152
rect 25136 25211 25188 25220
rect 25136 25177 25145 25211
rect 25145 25177 25179 25211
rect 25179 25177 25188 25211
rect 25136 25168 25188 25177
rect 27620 25168 27672 25220
rect 38108 25143 38160 25152
rect 38108 25109 38117 25143
rect 38117 25109 38151 25143
rect 38151 25109 38160 25143
rect 38108 25100 38160 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 9956 24896 10008 24948
rect 13636 24896 13688 24948
rect 21916 24896 21968 24948
rect 14924 24871 14976 24880
rect 14924 24837 14933 24871
rect 14933 24837 14967 24871
rect 14967 24837 14976 24871
rect 14924 24828 14976 24837
rect 22192 24871 22244 24880
rect 22192 24837 22201 24871
rect 22201 24837 22235 24871
rect 22235 24837 22244 24871
rect 22192 24828 22244 24837
rect 27344 24896 27396 24948
rect 5356 24803 5408 24812
rect 5356 24769 5365 24803
rect 5365 24769 5399 24803
rect 5399 24769 5408 24803
rect 5356 24760 5408 24769
rect 6276 24760 6328 24812
rect 10784 24760 10836 24812
rect 12900 24760 12952 24812
rect 12624 24692 12676 24744
rect 13452 24760 13504 24812
rect 27988 24828 28040 24880
rect 13360 24692 13412 24744
rect 14832 24735 14884 24744
rect 14832 24701 14841 24735
rect 14841 24701 14875 24735
rect 14875 24701 14884 24735
rect 14832 24692 14884 24701
rect 15476 24735 15528 24744
rect 15476 24701 15485 24735
rect 15485 24701 15519 24735
rect 15519 24701 15528 24735
rect 15476 24692 15528 24701
rect 19616 24692 19668 24744
rect 28264 24692 28316 24744
rect 14556 24624 14608 24676
rect 21916 24624 21968 24676
rect 22652 24667 22704 24676
rect 22652 24633 22661 24667
rect 22661 24633 22695 24667
rect 22695 24633 22704 24667
rect 22652 24624 22704 24633
rect 5356 24556 5408 24608
rect 8392 24556 8444 24608
rect 12808 24556 12860 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 4620 24352 4672 24404
rect 14924 24352 14976 24404
rect 20904 24352 20956 24404
rect 25136 24352 25188 24404
rect 31944 24352 31996 24404
rect 1584 24191 1636 24200
rect 1584 24157 1593 24191
rect 1593 24157 1627 24191
rect 1627 24157 1636 24191
rect 1584 24148 1636 24157
rect 6368 24148 6420 24200
rect 7748 24191 7800 24200
rect 7748 24157 7757 24191
rect 7757 24157 7791 24191
rect 7791 24157 7800 24191
rect 7748 24148 7800 24157
rect 10784 24148 10836 24200
rect 16672 24216 16724 24268
rect 22560 24284 22612 24336
rect 18880 24259 18932 24268
rect 18880 24225 18889 24259
rect 18889 24225 18923 24259
rect 18923 24225 18932 24259
rect 18880 24216 18932 24225
rect 19616 24259 19668 24268
rect 19616 24225 19625 24259
rect 19625 24225 19659 24259
rect 19659 24225 19668 24259
rect 19616 24216 19668 24225
rect 19984 24259 20036 24268
rect 19984 24225 19993 24259
rect 19993 24225 20027 24259
rect 20027 24225 20036 24259
rect 19984 24216 20036 24225
rect 20812 24216 20864 24268
rect 22652 24216 22704 24268
rect 26240 24216 26292 24268
rect 13636 24191 13688 24200
rect 13636 24157 13645 24191
rect 13645 24157 13679 24191
rect 13679 24157 13688 24191
rect 13636 24148 13688 24157
rect 16948 24148 17000 24200
rect 20720 24191 20772 24200
rect 20720 24157 20729 24191
rect 20729 24157 20763 24191
rect 20763 24157 20772 24191
rect 20720 24148 20772 24157
rect 21180 24148 21232 24200
rect 24860 24148 24912 24200
rect 38108 24216 38160 24268
rect 7288 24080 7340 24132
rect 1768 24055 1820 24064
rect 1768 24021 1777 24055
rect 1777 24021 1811 24055
rect 1811 24021 1820 24055
rect 1768 24012 1820 24021
rect 8208 24055 8260 24064
rect 8208 24021 8217 24055
rect 8217 24021 8251 24055
rect 8251 24021 8260 24055
rect 8208 24012 8260 24021
rect 10508 24055 10560 24064
rect 10508 24021 10517 24055
rect 10517 24021 10551 24055
rect 10551 24021 10560 24055
rect 10508 24012 10560 24021
rect 12348 24012 12400 24064
rect 18328 24123 18380 24132
rect 18328 24089 18337 24123
rect 18337 24089 18371 24123
rect 18371 24089 18380 24123
rect 18328 24080 18380 24089
rect 31392 24148 31444 24200
rect 38292 24191 38344 24200
rect 38292 24157 38301 24191
rect 38301 24157 38335 24191
rect 38335 24157 38344 24191
rect 38292 24148 38344 24157
rect 22652 24012 22704 24064
rect 24676 24012 24728 24064
rect 25964 24012 26016 24064
rect 28448 24055 28500 24064
rect 28448 24021 28457 24055
rect 28457 24021 28491 24055
rect 28491 24021 28500 24055
rect 28448 24012 28500 24021
rect 33508 24012 33560 24064
rect 37004 24012 37056 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 1584 23808 1636 23860
rect 8208 23808 8260 23860
rect 12808 23851 12860 23860
rect 12808 23817 12817 23851
rect 12817 23817 12851 23851
rect 12851 23817 12860 23851
rect 12808 23808 12860 23817
rect 13360 23851 13412 23860
rect 13360 23817 13369 23851
rect 13369 23817 13403 23851
rect 13403 23817 13412 23851
rect 13360 23808 13412 23817
rect 22192 23808 22244 23860
rect 14372 23740 14424 23792
rect 17040 23783 17092 23792
rect 17040 23749 17049 23783
rect 17049 23749 17083 23783
rect 17083 23749 17092 23783
rect 17040 23740 17092 23749
rect 9220 23672 9272 23724
rect 10508 23715 10560 23724
rect 10508 23681 10517 23715
rect 10517 23681 10551 23715
rect 10551 23681 10560 23715
rect 10508 23672 10560 23681
rect 10968 23672 11020 23724
rect 12348 23715 12400 23724
rect 12348 23681 12357 23715
rect 12357 23681 12391 23715
rect 12391 23681 12400 23715
rect 12348 23672 12400 23681
rect 13636 23672 13688 23724
rect 15016 23715 15068 23724
rect 15016 23681 15025 23715
rect 15025 23681 15059 23715
rect 15059 23681 15068 23715
rect 15016 23672 15068 23681
rect 21272 23715 21324 23724
rect 21272 23681 21281 23715
rect 21281 23681 21315 23715
rect 21315 23681 21324 23715
rect 21272 23672 21324 23681
rect 12164 23647 12216 23656
rect 12164 23613 12173 23647
rect 12173 23613 12207 23647
rect 12207 23613 12216 23647
rect 12164 23604 12216 23613
rect 16672 23604 16724 23656
rect 27804 23808 27856 23860
rect 28540 23808 28592 23860
rect 32128 23808 32180 23860
rect 33324 23851 33376 23860
rect 33324 23817 33333 23851
rect 33333 23817 33367 23851
rect 33367 23817 33376 23851
rect 33324 23808 33376 23817
rect 22652 23783 22704 23792
rect 22652 23749 22661 23783
rect 22661 23749 22695 23783
rect 22695 23749 22704 23783
rect 22652 23740 22704 23749
rect 29184 23715 29236 23724
rect 29184 23681 29193 23715
rect 29193 23681 29227 23715
rect 29227 23681 29236 23715
rect 29184 23672 29236 23681
rect 32496 23715 32548 23724
rect 32496 23681 32505 23715
rect 32505 23681 32539 23715
rect 32539 23681 32548 23715
rect 32496 23672 32548 23681
rect 33508 23715 33560 23724
rect 33508 23681 33517 23715
rect 33517 23681 33551 23715
rect 33551 23681 33560 23715
rect 33508 23672 33560 23681
rect 16580 23536 16632 23588
rect 14464 23468 14516 23520
rect 19984 23468 20036 23520
rect 27252 23468 27304 23520
rect 29276 23511 29328 23520
rect 29276 23477 29285 23511
rect 29285 23477 29319 23511
rect 29319 23477 29328 23511
rect 29276 23468 29328 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 7748 23264 7800 23316
rect 11704 23264 11756 23316
rect 14924 23264 14976 23316
rect 16212 23307 16264 23316
rect 16212 23273 16221 23307
rect 16221 23273 16255 23307
rect 16255 23273 16264 23307
rect 16212 23264 16264 23273
rect 16764 23264 16816 23316
rect 18328 23264 18380 23316
rect 21180 23264 21232 23316
rect 9404 23196 9456 23248
rect 16672 23196 16724 23248
rect 19432 23196 19484 23248
rect 22008 23196 22060 23248
rect 12164 23171 12216 23180
rect 12164 23137 12173 23171
rect 12173 23137 12207 23171
rect 12207 23137 12216 23171
rect 12164 23128 12216 23137
rect 14372 23171 14424 23180
rect 14372 23137 14381 23171
rect 14381 23137 14415 23171
rect 14415 23137 14424 23171
rect 14372 23128 14424 23137
rect 6460 23060 6512 23112
rect 11704 23060 11756 23112
rect 16028 23103 16080 23112
rect 14464 23035 14516 23044
rect 14464 23001 14473 23035
rect 14473 23001 14507 23035
rect 14507 23001 14516 23035
rect 14464 22992 14516 23001
rect 11336 22924 11388 22976
rect 16028 23069 16037 23103
rect 16037 23069 16071 23103
rect 16071 23069 16080 23103
rect 16028 23060 16080 23069
rect 19340 23128 19392 23180
rect 20812 23128 20864 23180
rect 27436 23264 27488 23316
rect 29184 23264 29236 23316
rect 29736 23196 29788 23248
rect 19984 23060 20036 23112
rect 18512 22992 18564 23044
rect 19340 22992 19392 23044
rect 21272 23060 21324 23112
rect 24860 23060 24912 23112
rect 28264 23171 28316 23180
rect 28264 23137 28273 23171
rect 28273 23137 28307 23171
rect 28307 23137 28316 23171
rect 28264 23128 28316 23137
rect 29276 23128 29328 23180
rect 27160 23103 27212 23112
rect 27160 23069 27169 23103
rect 27169 23069 27203 23103
rect 27203 23069 27212 23103
rect 27160 23060 27212 23069
rect 28356 23060 28408 23112
rect 32496 23264 32548 23316
rect 31392 23103 31444 23112
rect 26424 22992 26476 23044
rect 31392 23069 31401 23103
rect 31401 23069 31435 23103
rect 31435 23069 31444 23103
rect 31392 23060 31444 23069
rect 37004 23060 37056 23112
rect 31852 22992 31904 23044
rect 19432 22924 19484 22976
rect 20076 22924 20128 22976
rect 22100 22924 22152 22976
rect 25872 22924 25924 22976
rect 28264 22924 28316 22976
rect 30564 22924 30616 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 15016 22720 15068 22772
rect 17040 22720 17092 22772
rect 18512 22720 18564 22772
rect 5356 22695 5408 22704
rect 5356 22661 5365 22695
rect 5365 22661 5399 22695
rect 5399 22661 5408 22695
rect 5356 22652 5408 22661
rect 5724 22652 5776 22704
rect 8852 22695 8904 22704
rect 8852 22661 8861 22695
rect 8861 22661 8895 22695
rect 8895 22661 8904 22695
rect 8852 22652 8904 22661
rect 9404 22695 9456 22704
rect 9404 22661 9413 22695
rect 9413 22661 9447 22695
rect 9447 22661 9456 22695
rect 9404 22652 9456 22661
rect 11888 22695 11940 22704
rect 11888 22661 11897 22695
rect 11897 22661 11931 22695
rect 11931 22661 11940 22695
rect 11888 22652 11940 22661
rect 1768 22627 1820 22636
rect 1768 22593 1777 22627
rect 1777 22593 1811 22627
rect 1811 22593 1820 22627
rect 1768 22584 1820 22593
rect 3148 22627 3200 22636
rect 3148 22593 3157 22627
rect 3157 22593 3191 22627
rect 3191 22593 3200 22627
rect 3148 22584 3200 22593
rect 14188 22652 14240 22704
rect 19984 22720 20036 22772
rect 21272 22763 21324 22772
rect 21272 22729 21281 22763
rect 21281 22729 21315 22763
rect 21315 22729 21324 22763
rect 21272 22720 21324 22729
rect 22376 22695 22428 22704
rect 15660 22584 15712 22636
rect 16120 22627 16172 22636
rect 16120 22593 16129 22627
rect 16129 22593 16163 22627
rect 16163 22593 16172 22627
rect 16120 22584 16172 22593
rect 16856 22584 16908 22636
rect 17776 22584 17828 22636
rect 22376 22661 22385 22695
rect 22385 22661 22419 22695
rect 22419 22661 22428 22695
rect 22376 22652 22428 22661
rect 6000 22516 6052 22568
rect 10140 22516 10192 22568
rect 11796 22559 11848 22568
rect 11796 22525 11805 22559
rect 11805 22525 11839 22559
rect 11839 22525 11848 22559
rect 11796 22516 11848 22525
rect 11980 22516 12032 22568
rect 12256 22516 12308 22568
rect 5816 22448 5868 22500
rect 8116 22448 8168 22500
rect 16948 22491 17000 22500
rect 16948 22457 16957 22491
rect 16957 22457 16991 22491
rect 16991 22457 17000 22491
rect 16948 22448 17000 22457
rect 19156 22584 19208 22636
rect 20720 22584 20772 22636
rect 20996 22584 21048 22636
rect 22008 22516 22060 22568
rect 22560 22559 22612 22568
rect 22560 22525 22569 22559
rect 22569 22525 22603 22559
rect 22603 22525 22612 22559
rect 22560 22516 22612 22525
rect 3240 22423 3292 22432
rect 3240 22389 3249 22423
rect 3249 22389 3283 22423
rect 3283 22389 3292 22423
rect 3240 22380 3292 22389
rect 13268 22423 13320 22432
rect 13268 22389 13277 22423
rect 13277 22389 13311 22423
rect 13311 22389 13320 22423
rect 13268 22380 13320 22389
rect 17960 22380 18012 22432
rect 28356 22720 28408 22772
rect 23664 22695 23716 22704
rect 23664 22661 23673 22695
rect 23673 22661 23707 22695
rect 23707 22661 23716 22695
rect 23664 22652 23716 22661
rect 24216 22695 24268 22704
rect 24216 22661 24225 22695
rect 24225 22661 24259 22695
rect 24259 22661 24268 22695
rect 24216 22652 24268 22661
rect 25872 22695 25924 22704
rect 25872 22661 25881 22695
rect 25881 22661 25915 22695
rect 25915 22661 25924 22695
rect 25872 22652 25924 22661
rect 27620 22652 27672 22704
rect 27896 22652 27948 22704
rect 27436 22584 27488 22636
rect 28448 22627 28500 22636
rect 25504 22516 25556 22568
rect 25780 22559 25832 22568
rect 25780 22525 25789 22559
rect 25789 22525 25823 22559
rect 25823 22525 25832 22559
rect 25780 22516 25832 22525
rect 28448 22593 28457 22627
rect 28457 22593 28491 22627
rect 28491 22593 28500 22627
rect 28448 22584 28500 22593
rect 32128 22584 32180 22636
rect 28632 22559 28684 22568
rect 28632 22525 28641 22559
rect 28641 22525 28675 22559
rect 28675 22525 28684 22559
rect 28632 22516 28684 22525
rect 30656 22559 30708 22568
rect 30656 22525 30665 22559
rect 30665 22525 30699 22559
rect 30699 22525 30708 22559
rect 30656 22516 30708 22525
rect 31116 22448 31168 22500
rect 29000 22423 29052 22432
rect 29000 22389 29009 22423
rect 29009 22389 29043 22423
rect 29043 22389 29052 22423
rect 29000 22380 29052 22389
rect 30380 22380 30432 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 8852 22176 8904 22228
rect 16028 22176 16080 22228
rect 27160 22176 27212 22228
rect 28632 22176 28684 22228
rect 30380 22219 30432 22228
rect 30380 22185 30389 22219
rect 30389 22185 30423 22219
rect 30423 22185 30432 22219
rect 30380 22176 30432 22185
rect 30656 22176 30708 22228
rect 5264 22108 5316 22160
rect 16120 22108 16172 22160
rect 17776 22108 17828 22160
rect 6368 22083 6420 22092
rect 6368 22049 6377 22083
rect 6377 22049 6411 22083
rect 6411 22049 6420 22083
rect 6368 22040 6420 22049
rect 9956 22040 10008 22092
rect 10140 22083 10192 22092
rect 10140 22049 10149 22083
rect 10149 22049 10183 22083
rect 10183 22049 10192 22083
rect 10140 22040 10192 22049
rect 11796 22040 11848 22092
rect 13084 22040 13136 22092
rect 5816 21972 5868 22024
rect 8668 21972 8720 22024
rect 7104 21947 7156 21956
rect 7104 21913 7113 21947
rect 7113 21913 7147 21947
rect 7147 21913 7156 21947
rect 7104 21904 7156 21913
rect 7288 21904 7340 21956
rect 10876 21972 10928 22024
rect 13268 22015 13320 22024
rect 13268 21981 13277 22015
rect 13277 21981 13311 22015
rect 13311 21981 13320 22015
rect 13268 21972 13320 21981
rect 17868 22040 17920 22092
rect 21088 22040 21140 22092
rect 21824 22040 21876 22092
rect 16764 22015 16816 22024
rect 16764 21981 16773 22015
rect 16773 21981 16807 22015
rect 16807 21981 16816 22015
rect 16764 21972 16816 21981
rect 16948 22015 17000 22024
rect 16948 21981 16957 22015
rect 16957 21981 16991 22015
rect 16991 21981 17000 22015
rect 16948 21972 17000 21981
rect 20536 21972 20588 22024
rect 20996 21972 21048 22024
rect 19340 21904 19392 21956
rect 19984 21904 20036 21956
rect 22008 21947 22060 21956
rect 22008 21913 22017 21947
rect 22017 21913 22051 21947
rect 22051 21913 22060 21947
rect 22008 21904 22060 21913
rect 22100 21947 22152 21956
rect 22100 21913 22109 21947
rect 22109 21913 22143 21947
rect 22143 21913 22152 21947
rect 23664 22040 23716 22092
rect 24676 22083 24728 22092
rect 24676 22049 24685 22083
rect 24685 22049 24719 22083
rect 24719 22049 24728 22083
rect 24676 22040 24728 22049
rect 25780 22040 25832 22092
rect 29736 22083 29788 22092
rect 29736 22049 29745 22083
rect 29745 22049 29779 22083
rect 29779 22049 29788 22083
rect 29736 22040 29788 22049
rect 22928 21972 22980 22024
rect 25688 21972 25740 22024
rect 26424 21972 26476 22024
rect 27804 21972 27856 22024
rect 29276 21972 29328 22024
rect 31024 22015 31076 22024
rect 31024 21981 31033 22015
rect 31033 21981 31067 22015
rect 31067 21981 31076 22015
rect 31024 21972 31076 21981
rect 37464 22015 37516 22024
rect 37464 21981 37473 22015
rect 37473 21981 37507 22015
rect 37507 21981 37516 22015
rect 37464 21972 37516 21981
rect 37740 22015 37792 22024
rect 37740 21981 37749 22015
rect 37749 21981 37783 22015
rect 37783 21981 37792 22015
rect 37740 21972 37792 21981
rect 22100 21904 22152 21913
rect 29736 21904 29788 21956
rect 8300 21879 8352 21888
rect 8300 21845 8309 21879
rect 8309 21845 8343 21879
rect 8343 21845 8352 21879
rect 8300 21836 8352 21845
rect 9956 21836 10008 21888
rect 12164 21836 12216 21888
rect 13084 21879 13136 21888
rect 13084 21845 13093 21879
rect 13093 21845 13127 21879
rect 13127 21845 13136 21879
rect 13084 21836 13136 21845
rect 20260 21879 20312 21888
rect 20260 21845 20269 21879
rect 20269 21845 20303 21879
rect 20303 21845 20312 21879
rect 20260 21836 20312 21845
rect 22192 21836 22244 21888
rect 28080 21879 28132 21888
rect 28080 21845 28089 21879
rect 28089 21845 28123 21879
rect 28123 21845 28132 21879
rect 28080 21836 28132 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 7104 21675 7156 21684
rect 7104 21641 7113 21675
rect 7113 21641 7147 21675
rect 7147 21641 7156 21675
rect 7104 21632 7156 21641
rect 8668 21675 8720 21684
rect 8668 21641 8677 21675
rect 8677 21641 8711 21675
rect 8711 21641 8720 21675
rect 8668 21632 8720 21641
rect 10876 21675 10928 21684
rect 9864 21607 9916 21616
rect 9864 21573 9873 21607
rect 9873 21573 9907 21607
rect 9907 21573 9916 21607
rect 9864 21564 9916 21573
rect 10876 21641 10885 21675
rect 10885 21641 10919 21675
rect 10919 21641 10928 21675
rect 10876 21632 10928 21641
rect 11888 21632 11940 21684
rect 12164 21632 12216 21684
rect 16212 21632 16264 21684
rect 15936 21564 15988 21616
rect 17960 21607 18012 21616
rect 17960 21573 17969 21607
rect 17969 21573 18003 21607
rect 18003 21573 18012 21607
rect 17960 21564 18012 21573
rect 20076 21564 20128 21616
rect 20628 21564 20680 21616
rect 7012 21496 7064 21548
rect 9588 21496 9640 21548
rect 11060 21539 11112 21548
rect 11060 21505 11069 21539
rect 11069 21505 11103 21539
rect 11103 21505 11112 21539
rect 11060 21496 11112 21505
rect 12256 21539 12308 21548
rect 12256 21505 12265 21539
rect 12265 21505 12299 21539
rect 12299 21505 12308 21539
rect 12256 21496 12308 21505
rect 15108 21496 15160 21548
rect 17592 21496 17644 21548
rect 7932 21471 7984 21480
rect 7932 21437 7941 21471
rect 7941 21437 7975 21471
rect 7975 21437 7984 21471
rect 7932 21428 7984 21437
rect 11152 21428 11204 21480
rect 13452 21471 13504 21480
rect 8668 21360 8720 21412
rect 13452 21437 13461 21471
rect 13461 21437 13495 21471
rect 13495 21437 13504 21471
rect 13452 21428 13504 21437
rect 17868 21471 17920 21480
rect 17868 21437 17877 21471
rect 17877 21437 17911 21471
rect 17911 21437 17920 21471
rect 17868 21428 17920 21437
rect 19800 21471 19852 21480
rect 15108 21360 15160 21412
rect 19800 21437 19809 21471
rect 19809 21437 19843 21471
rect 19843 21437 19852 21471
rect 19800 21428 19852 21437
rect 19800 21292 19852 21344
rect 20352 21292 20404 21344
rect 20536 21292 20588 21344
rect 22008 21632 22060 21684
rect 29000 21632 29052 21684
rect 29276 21675 29328 21684
rect 29276 21641 29285 21675
rect 29285 21641 29319 21675
rect 29319 21641 29328 21675
rect 29276 21632 29328 21641
rect 31024 21632 31076 21684
rect 22192 21607 22244 21616
rect 22192 21573 22201 21607
rect 22201 21573 22235 21607
rect 22235 21573 22244 21607
rect 22192 21564 22244 21573
rect 28080 21539 28132 21548
rect 28080 21505 28089 21539
rect 28089 21505 28123 21539
rect 28123 21505 28132 21539
rect 28080 21496 28132 21505
rect 29184 21539 29236 21548
rect 29184 21505 29193 21539
rect 29193 21505 29227 21539
rect 29227 21505 29236 21539
rect 29184 21496 29236 21505
rect 22100 21471 22152 21480
rect 22100 21437 22109 21471
rect 22109 21437 22143 21471
rect 22143 21437 22152 21471
rect 22100 21428 22152 21437
rect 28264 21471 28316 21480
rect 21824 21360 21876 21412
rect 28264 21437 28273 21471
rect 28273 21437 28307 21471
rect 28307 21437 28316 21471
rect 28264 21428 28316 21437
rect 25688 21292 25740 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 6000 21088 6052 21140
rect 7012 21131 7064 21140
rect 7012 21097 7021 21131
rect 7021 21097 7055 21131
rect 7055 21097 7064 21131
rect 7012 21088 7064 21097
rect 9220 21131 9272 21140
rect 9220 21097 9229 21131
rect 9229 21097 9263 21131
rect 9263 21097 9272 21131
rect 9220 21088 9272 21097
rect 9864 21131 9916 21140
rect 9864 21097 9873 21131
rect 9873 21097 9907 21131
rect 9907 21097 9916 21131
rect 9864 21088 9916 21097
rect 16948 21088 17000 21140
rect 17868 21088 17920 21140
rect 23480 21088 23532 21140
rect 28264 21131 28316 21140
rect 28264 21097 28273 21131
rect 28273 21097 28307 21131
rect 28307 21097 28316 21131
rect 28264 21088 28316 21097
rect 7932 20995 7984 21004
rect 7932 20961 7941 20995
rect 7941 20961 7975 20995
rect 7975 20961 7984 20995
rect 7932 20952 7984 20961
rect 17592 21020 17644 21072
rect 1768 20927 1820 20936
rect 1768 20893 1777 20927
rect 1777 20893 1811 20927
rect 1811 20893 1820 20927
rect 1768 20884 1820 20893
rect 3792 20884 3844 20936
rect 7656 20884 7708 20936
rect 10048 20927 10100 20936
rect 10048 20893 10057 20927
rect 10057 20893 10091 20927
rect 10091 20893 10100 20927
rect 10048 20884 10100 20893
rect 12440 20884 12492 20936
rect 12992 20927 13044 20936
rect 12992 20893 13001 20927
rect 13001 20893 13035 20927
rect 13035 20893 13044 20927
rect 12992 20884 13044 20893
rect 14556 20927 14608 20936
rect 14556 20893 14565 20927
rect 14565 20893 14599 20927
rect 14599 20893 14608 20927
rect 14556 20884 14608 20893
rect 14924 20884 14976 20936
rect 8300 20816 8352 20868
rect 5356 20748 5408 20800
rect 8116 20748 8168 20800
rect 15108 20816 15160 20868
rect 15200 20859 15252 20868
rect 15200 20825 15209 20859
rect 15209 20825 15243 20859
rect 15243 20825 15252 20859
rect 17408 20859 17460 20868
rect 15200 20816 15252 20825
rect 17408 20825 17417 20859
rect 17417 20825 17451 20859
rect 17451 20825 17460 20859
rect 17408 20816 17460 20825
rect 20628 20952 20680 21004
rect 19432 20927 19484 20936
rect 19432 20893 19441 20927
rect 19441 20893 19475 20927
rect 19475 20893 19484 20927
rect 19432 20884 19484 20893
rect 20260 20884 20312 20936
rect 25596 20927 25648 20936
rect 25596 20893 25605 20927
rect 25605 20893 25639 20927
rect 25639 20893 25648 20927
rect 25596 20884 25648 20893
rect 27804 20927 27856 20936
rect 27804 20893 27813 20927
rect 27813 20893 27847 20927
rect 27847 20893 27856 20927
rect 27804 20884 27856 20893
rect 29736 20927 29788 20936
rect 29736 20893 29745 20927
rect 29745 20893 29779 20927
rect 29779 20893 29788 20927
rect 29736 20884 29788 20893
rect 30380 20927 30432 20936
rect 30380 20893 30389 20927
rect 30389 20893 30423 20927
rect 30423 20893 30432 20927
rect 30380 20884 30432 20893
rect 38292 20927 38344 20936
rect 38292 20893 38301 20927
rect 38301 20893 38335 20927
rect 38335 20893 38344 20927
rect 38292 20884 38344 20893
rect 14648 20748 14700 20800
rect 24768 20816 24820 20868
rect 19800 20748 19852 20800
rect 20260 20748 20312 20800
rect 20352 20748 20404 20800
rect 25412 20791 25464 20800
rect 25412 20757 25421 20791
rect 25421 20757 25455 20791
rect 25455 20757 25464 20791
rect 25412 20748 25464 20757
rect 29000 20748 29052 20800
rect 31484 20748 31536 20800
rect 34520 20748 34572 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 5724 20544 5776 20596
rect 11060 20544 11112 20596
rect 19432 20544 19484 20596
rect 21272 20544 21324 20596
rect 25596 20544 25648 20596
rect 8116 20519 8168 20528
rect 8116 20485 8125 20519
rect 8125 20485 8159 20519
rect 8159 20485 8168 20519
rect 8116 20476 8168 20485
rect 9772 20476 9824 20528
rect 20444 20476 20496 20528
rect 20812 20476 20864 20528
rect 25412 20476 25464 20528
rect 3240 20408 3292 20460
rect 5816 20451 5868 20460
rect 5816 20417 5825 20451
rect 5825 20417 5859 20451
rect 5859 20417 5868 20451
rect 5816 20408 5868 20417
rect 7656 20408 7708 20460
rect 4620 20340 4672 20392
rect 5632 20340 5684 20392
rect 12348 20408 12400 20460
rect 13084 20408 13136 20460
rect 14648 20451 14700 20460
rect 14648 20417 14657 20451
rect 14657 20417 14691 20451
rect 14691 20417 14700 20451
rect 14648 20408 14700 20417
rect 25136 20451 25188 20460
rect 15844 20383 15896 20392
rect 15844 20349 15853 20383
rect 15853 20349 15887 20383
rect 15887 20349 15896 20383
rect 15844 20340 15896 20349
rect 16488 20340 16540 20392
rect 21364 20340 21416 20392
rect 8668 20315 8720 20324
rect 8668 20281 8677 20315
rect 8677 20281 8711 20315
rect 8711 20281 8720 20315
rect 8668 20272 8720 20281
rect 11152 20272 11204 20324
rect 25136 20417 25145 20451
rect 25145 20417 25179 20451
rect 25179 20417 25188 20451
rect 25136 20408 25188 20417
rect 23480 20383 23532 20392
rect 23480 20349 23489 20383
rect 23489 20349 23523 20383
rect 23523 20349 23532 20383
rect 23480 20340 23532 20349
rect 25688 20408 25740 20460
rect 28172 20408 28224 20460
rect 29000 20408 29052 20460
rect 5080 20204 5132 20256
rect 5172 20204 5224 20256
rect 9312 20204 9364 20256
rect 14372 20204 14424 20256
rect 15384 20204 15436 20256
rect 21180 20247 21232 20256
rect 21180 20213 21189 20247
rect 21189 20213 21223 20247
rect 21223 20213 21232 20247
rect 21180 20204 21232 20213
rect 22100 20204 22152 20256
rect 22744 20272 22796 20324
rect 24032 20315 24084 20324
rect 24032 20281 24041 20315
rect 24041 20281 24075 20315
rect 24075 20281 24084 20315
rect 24032 20272 24084 20281
rect 30472 20544 30524 20596
rect 29368 20519 29420 20528
rect 29368 20485 29377 20519
rect 29377 20485 29411 20519
rect 29411 20485 29420 20519
rect 29368 20476 29420 20485
rect 30748 20340 30800 20392
rect 29828 20315 29880 20324
rect 29828 20281 29837 20315
rect 29837 20281 29871 20315
rect 29871 20281 29880 20315
rect 29828 20272 29880 20281
rect 25872 20204 25924 20256
rect 27344 20204 27396 20256
rect 30104 20204 30156 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 10048 20000 10100 20052
rect 12256 20000 12308 20052
rect 13452 20000 13504 20052
rect 15200 20000 15252 20052
rect 15936 20000 15988 20052
rect 20076 20000 20128 20052
rect 21364 20043 21416 20052
rect 21364 20009 21373 20043
rect 21373 20009 21407 20043
rect 21407 20009 21416 20043
rect 21364 20000 21416 20009
rect 29368 20000 29420 20052
rect 30748 20043 30800 20052
rect 30748 20009 30757 20043
rect 30757 20009 30791 20043
rect 30791 20009 30800 20043
rect 30748 20000 30800 20009
rect 6092 19932 6144 19984
rect 14096 19932 14148 19984
rect 16580 19932 16632 19984
rect 20168 19932 20220 19984
rect 5080 19907 5132 19916
rect 5080 19873 5089 19907
rect 5089 19873 5123 19907
rect 5123 19873 5132 19907
rect 5080 19864 5132 19873
rect 7288 19864 7340 19916
rect 11980 19864 12032 19916
rect 15016 19864 15068 19916
rect 9312 19796 9364 19848
rect 9956 19839 10008 19848
rect 9956 19805 9965 19839
rect 9965 19805 9999 19839
rect 9999 19805 10008 19839
rect 9956 19796 10008 19805
rect 12072 19796 12124 19848
rect 12348 19796 12400 19848
rect 15108 19839 15160 19848
rect 5172 19771 5224 19780
rect 5172 19737 5181 19771
rect 5181 19737 5215 19771
rect 5215 19737 5224 19771
rect 10508 19771 10560 19780
rect 5172 19728 5224 19737
rect 10508 19737 10517 19771
rect 10517 19737 10551 19771
rect 10551 19737 10560 19771
rect 10508 19728 10560 19737
rect 12164 19728 12216 19780
rect 7288 19660 7340 19712
rect 15108 19805 15117 19839
rect 15117 19805 15151 19839
rect 15151 19805 15160 19839
rect 15108 19796 15160 19805
rect 15936 19796 15988 19848
rect 16764 19864 16816 19916
rect 18328 19864 18380 19916
rect 18880 19864 18932 19916
rect 22744 19864 22796 19916
rect 24768 19932 24820 19984
rect 29828 19932 29880 19984
rect 26332 19907 26384 19916
rect 26332 19873 26341 19907
rect 26341 19873 26375 19907
rect 26375 19873 26384 19907
rect 26332 19864 26384 19873
rect 27712 19864 27764 19916
rect 19340 19796 19392 19848
rect 20628 19796 20680 19848
rect 28172 19796 28224 19848
rect 16948 19728 17000 19780
rect 17224 19771 17276 19780
rect 17224 19737 17233 19771
rect 17233 19737 17267 19771
rect 17267 19737 17276 19771
rect 17224 19728 17276 19737
rect 17592 19728 17644 19780
rect 15660 19660 15712 19712
rect 19432 19660 19484 19712
rect 22652 19771 22704 19780
rect 22652 19737 22661 19771
rect 22661 19737 22695 19771
rect 22695 19737 22704 19771
rect 25688 19771 25740 19780
rect 22652 19728 22704 19737
rect 25688 19737 25697 19771
rect 25697 19737 25731 19771
rect 25731 19737 25740 19771
rect 25688 19728 25740 19737
rect 25872 19728 25924 19780
rect 27160 19728 27212 19780
rect 30472 19864 30524 19916
rect 29736 19796 29788 19848
rect 34520 19864 34572 19916
rect 31300 19703 31352 19712
rect 31300 19669 31309 19703
rect 31309 19669 31343 19703
rect 31343 19669 31352 19703
rect 31300 19660 31352 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 5080 19456 5132 19508
rect 9772 19499 9824 19508
rect 9772 19465 9781 19499
rect 9781 19465 9815 19499
rect 9815 19465 9824 19499
rect 9772 19456 9824 19465
rect 6828 19388 6880 19440
rect 12900 19456 12952 19508
rect 17224 19456 17276 19508
rect 17592 19456 17644 19508
rect 3424 19320 3476 19372
rect 5448 19320 5500 19372
rect 9956 19320 10008 19372
rect 10692 19320 10744 19372
rect 11520 19320 11572 19372
rect 13636 19388 13688 19440
rect 16488 19388 16540 19440
rect 17960 19431 18012 19440
rect 17960 19397 17969 19431
rect 17969 19397 18003 19431
rect 18003 19397 18012 19431
rect 17960 19388 18012 19397
rect 20720 19456 20772 19508
rect 21180 19456 21232 19508
rect 22652 19456 22704 19508
rect 27160 19499 27212 19508
rect 27160 19465 27169 19499
rect 27169 19465 27203 19499
rect 27203 19465 27212 19499
rect 27160 19456 27212 19465
rect 25688 19388 25740 19440
rect 32588 19388 32640 19440
rect 15200 19363 15252 19372
rect 15200 19329 15209 19363
rect 15209 19329 15243 19363
rect 15243 19329 15252 19363
rect 15200 19320 15252 19329
rect 17040 19320 17092 19372
rect 17316 19363 17368 19372
rect 17316 19329 17325 19363
rect 17325 19329 17359 19363
rect 17359 19329 17368 19363
rect 17316 19320 17368 19329
rect 19432 19363 19484 19372
rect 19432 19329 19441 19363
rect 19441 19329 19475 19363
rect 19475 19329 19484 19363
rect 19432 19320 19484 19329
rect 20536 19320 20588 19372
rect 22100 19320 22152 19372
rect 25136 19320 25188 19372
rect 27344 19363 27396 19372
rect 27344 19329 27353 19363
rect 27353 19329 27387 19363
rect 27387 19329 27396 19363
rect 27344 19320 27396 19329
rect 30104 19320 30156 19372
rect 14096 19295 14148 19304
rect 14096 19261 14105 19295
rect 14105 19261 14139 19295
rect 14139 19261 14148 19295
rect 14096 19252 14148 19261
rect 15384 19295 15436 19304
rect 15384 19261 15393 19295
rect 15393 19261 15427 19295
rect 15427 19261 15436 19295
rect 15384 19252 15436 19261
rect 19248 19252 19300 19304
rect 20168 19295 20220 19304
rect 20168 19261 20177 19295
rect 20177 19261 20211 19295
rect 20211 19261 20220 19295
rect 20168 19252 20220 19261
rect 20352 19295 20404 19304
rect 20352 19261 20361 19295
rect 20361 19261 20395 19295
rect 20395 19261 20404 19295
rect 20352 19252 20404 19261
rect 29828 19295 29880 19304
rect 29828 19261 29837 19295
rect 29837 19261 29871 19295
rect 29871 19261 29880 19295
rect 29828 19252 29880 19261
rect 31300 19252 31352 19304
rect 32680 19184 32732 19236
rect 1768 19159 1820 19168
rect 1768 19125 1777 19159
rect 1777 19125 1811 19159
rect 1811 19125 1820 19159
rect 1768 19116 1820 19125
rect 5816 19116 5868 19168
rect 14188 19116 14240 19168
rect 14832 19116 14884 19168
rect 18788 19116 18840 19168
rect 22100 19116 22152 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 4620 18912 4672 18964
rect 14188 18912 14240 18964
rect 15108 18912 15160 18964
rect 15844 18912 15896 18964
rect 16396 18912 16448 18964
rect 20168 18912 20220 18964
rect 22376 18955 22428 18964
rect 22376 18921 22385 18955
rect 22385 18921 22419 18955
rect 22419 18921 22428 18955
rect 22376 18912 22428 18921
rect 4988 18844 5040 18896
rect 5632 18776 5684 18828
rect 5908 18776 5960 18828
rect 6092 18819 6144 18828
rect 6092 18785 6101 18819
rect 6101 18785 6135 18819
rect 6135 18785 6144 18819
rect 6092 18776 6144 18785
rect 9404 18844 9456 18896
rect 23572 18844 23624 18896
rect 16856 18776 16908 18828
rect 17040 18776 17092 18828
rect 18512 18776 18564 18828
rect 30564 18844 30616 18896
rect 5080 18751 5132 18760
rect 5080 18717 5089 18751
rect 5089 18717 5123 18751
rect 5123 18717 5132 18751
rect 5080 18708 5132 18717
rect 6920 18751 6972 18760
rect 6920 18717 6929 18751
rect 6929 18717 6963 18751
rect 6963 18717 6972 18751
rect 6920 18708 6972 18717
rect 7104 18751 7156 18760
rect 7104 18717 7113 18751
rect 7113 18717 7147 18751
rect 7147 18717 7156 18751
rect 7104 18708 7156 18717
rect 8024 18751 8076 18760
rect 8024 18717 8033 18751
rect 8033 18717 8067 18751
rect 8067 18717 8076 18751
rect 8024 18708 8076 18717
rect 11520 18708 11572 18760
rect 14648 18708 14700 18760
rect 14832 18708 14884 18760
rect 20812 18708 20864 18760
rect 21548 18751 21600 18760
rect 21548 18717 21557 18751
rect 21557 18717 21591 18751
rect 21591 18717 21600 18751
rect 21548 18708 21600 18717
rect 29828 18776 29880 18828
rect 22284 18751 22336 18760
rect 22284 18717 22293 18751
rect 22293 18717 22327 18751
rect 22327 18717 22336 18751
rect 22284 18708 22336 18717
rect 24768 18751 24820 18760
rect 24768 18717 24777 18751
rect 24777 18717 24811 18751
rect 24811 18717 24820 18751
rect 24768 18708 24820 18717
rect 28448 18708 28500 18760
rect 4804 18640 4856 18692
rect 5172 18572 5224 18624
rect 11980 18683 12032 18692
rect 11980 18649 11990 18683
rect 11990 18649 12024 18683
rect 12024 18649 12032 18683
rect 11980 18640 12032 18649
rect 7564 18615 7616 18624
rect 7564 18581 7573 18615
rect 7573 18581 7607 18615
rect 7607 18581 7616 18615
rect 7564 18572 7616 18581
rect 9220 18615 9272 18624
rect 9220 18581 9229 18615
rect 9229 18581 9263 18615
rect 9263 18581 9272 18615
rect 9220 18572 9272 18581
rect 12716 18640 12768 18692
rect 14188 18640 14240 18692
rect 16396 18640 16448 18692
rect 16948 18640 17000 18692
rect 19248 18640 19300 18692
rect 22008 18640 22060 18692
rect 19432 18572 19484 18624
rect 21364 18615 21416 18624
rect 21364 18581 21373 18615
rect 21373 18581 21407 18615
rect 21407 18581 21416 18615
rect 21364 18572 21416 18581
rect 24584 18572 24636 18624
rect 28080 18615 28132 18624
rect 28080 18581 28089 18615
rect 28089 18581 28123 18615
rect 28123 18581 28132 18615
rect 28080 18572 28132 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 3792 18368 3844 18420
rect 6920 18368 6972 18420
rect 12164 18411 12216 18420
rect 12164 18377 12173 18411
rect 12173 18377 12207 18411
rect 12207 18377 12216 18411
rect 12164 18368 12216 18377
rect 7380 18300 7432 18352
rect 9404 18343 9456 18352
rect 9404 18309 9413 18343
rect 9413 18309 9447 18343
rect 9447 18309 9456 18343
rect 9404 18300 9456 18309
rect 10232 18300 10284 18352
rect 12808 18343 12860 18352
rect 12808 18309 12817 18343
rect 12817 18309 12851 18343
rect 12851 18309 12860 18343
rect 12808 18300 12860 18309
rect 12900 18343 12952 18352
rect 12900 18309 12909 18343
rect 12909 18309 12943 18343
rect 12943 18309 12952 18343
rect 14188 18343 14240 18352
rect 12900 18300 12952 18309
rect 14188 18309 14197 18343
rect 14197 18309 14231 18343
rect 14231 18309 14240 18343
rect 14188 18300 14240 18309
rect 1768 18275 1820 18284
rect 1768 18241 1777 18275
rect 1777 18241 1811 18275
rect 1811 18241 1820 18275
rect 1768 18232 1820 18241
rect 5356 18275 5408 18284
rect 5356 18241 5365 18275
rect 5365 18241 5399 18275
rect 5399 18241 5408 18275
rect 5356 18232 5408 18241
rect 7288 18275 7340 18284
rect 7288 18241 7297 18275
rect 7297 18241 7331 18275
rect 7331 18241 7340 18275
rect 7288 18232 7340 18241
rect 10048 18275 10100 18284
rect 10048 18241 10057 18275
rect 10057 18241 10091 18275
rect 10091 18241 10100 18275
rect 10048 18232 10100 18241
rect 12072 18275 12124 18284
rect 12072 18241 12081 18275
rect 12081 18241 12115 18275
rect 12115 18241 12124 18275
rect 12072 18232 12124 18241
rect 17316 18368 17368 18420
rect 16856 18300 16908 18352
rect 17408 18275 17460 18284
rect 17408 18241 17417 18275
rect 17417 18241 17451 18275
rect 17451 18241 17460 18275
rect 17408 18232 17460 18241
rect 20812 18368 20864 18420
rect 24768 18368 24820 18420
rect 28448 18411 28500 18420
rect 28448 18377 28457 18411
rect 28457 18377 28491 18411
rect 28491 18377 28500 18411
rect 28448 18368 28500 18377
rect 18696 18343 18748 18352
rect 18696 18309 18705 18343
rect 18705 18309 18739 18343
rect 18739 18309 18748 18343
rect 18696 18300 18748 18309
rect 24584 18343 24636 18352
rect 24584 18309 24593 18343
rect 24593 18309 24627 18343
rect 24627 18309 24636 18343
rect 24584 18300 24636 18309
rect 20168 18232 20220 18284
rect 21364 18232 21416 18284
rect 22008 18275 22060 18284
rect 22008 18241 22017 18275
rect 22017 18241 22051 18275
rect 22051 18241 22060 18275
rect 22008 18232 22060 18241
rect 25688 18275 25740 18284
rect 7564 18164 7616 18216
rect 11060 18164 11112 18216
rect 12808 18164 12860 18216
rect 6828 18096 6880 18148
rect 11980 18028 12032 18080
rect 14372 18164 14424 18216
rect 14832 18164 14884 18216
rect 18604 18207 18656 18216
rect 18604 18173 18613 18207
rect 18613 18173 18647 18207
rect 18647 18173 18656 18207
rect 18604 18164 18656 18173
rect 22192 18207 22244 18216
rect 15844 18096 15896 18148
rect 22192 18173 22201 18207
rect 22201 18173 22235 18207
rect 22235 18173 22244 18207
rect 22192 18164 22244 18173
rect 25688 18241 25697 18275
rect 25697 18241 25731 18275
rect 25731 18241 25740 18275
rect 25688 18232 25740 18241
rect 27712 18232 27764 18284
rect 31208 18275 31260 18284
rect 24860 18164 24912 18216
rect 25964 18164 26016 18216
rect 27528 18207 27580 18216
rect 27528 18173 27537 18207
rect 27537 18173 27571 18207
rect 27571 18173 27580 18207
rect 27528 18164 27580 18173
rect 27620 18164 27672 18216
rect 31208 18241 31217 18275
rect 31217 18241 31251 18275
rect 31251 18241 31260 18275
rect 31208 18232 31260 18241
rect 29092 18207 29144 18216
rect 29092 18173 29101 18207
rect 29101 18173 29135 18207
rect 29135 18173 29144 18207
rect 29092 18164 29144 18173
rect 24400 18096 24452 18148
rect 17132 18028 17184 18080
rect 28264 18028 28316 18080
rect 31024 18071 31076 18080
rect 31024 18037 31033 18071
rect 31033 18037 31067 18071
rect 31067 18037 31076 18071
rect 31024 18028 31076 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 5448 17867 5500 17876
rect 5448 17833 5457 17867
rect 5457 17833 5491 17867
rect 5491 17833 5500 17867
rect 5448 17824 5500 17833
rect 10048 17824 10100 17876
rect 11060 17867 11112 17876
rect 11060 17833 11069 17867
rect 11069 17833 11103 17867
rect 11103 17833 11112 17867
rect 11060 17824 11112 17833
rect 13636 17867 13688 17876
rect 13636 17833 13645 17867
rect 13645 17833 13679 17867
rect 13679 17833 13688 17867
rect 13636 17824 13688 17833
rect 14188 17824 14240 17876
rect 17132 17824 17184 17876
rect 21548 17824 21600 17876
rect 22192 17824 22244 17876
rect 27528 17824 27580 17876
rect 8300 17756 8352 17808
rect 2320 17663 2372 17672
rect 2320 17629 2329 17663
rect 2329 17629 2363 17663
rect 2363 17629 2372 17663
rect 2320 17620 2372 17629
rect 5632 17663 5684 17672
rect 5632 17629 5641 17663
rect 5641 17629 5675 17663
rect 5675 17629 5684 17663
rect 5632 17620 5684 17629
rect 5908 17620 5960 17672
rect 6276 17663 6328 17672
rect 6276 17629 6285 17663
rect 6285 17629 6319 17663
rect 6319 17629 6328 17663
rect 6276 17620 6328 17629
rect 7748 17620 7800 17672
rect 7932 17620 7984 17672
rect 10416 17756 10468 17808
rect 10508 17756 10560 17808
rect 24124 17756 24176 17808
rect 28264 17756 28316 17808
rect 9220 17731 9272 17740
rect 9220 17697 9229 17731
rect 9229 17697 9263 17731
rect 9263 17697 9272 17731
rect 9220 17688 9272 17697
rect 11060 17688 11112 17740
rect 11336 17688 11388 17740
rect 12624 17688 12676 17740
rect 16396 17731 16448 17740
rect 16396 17697 16405 17731
rect 16405 17697 16439 17731
rect 16439 17697 16448 17731
rect 16396 17688 16448 17697
rect 16580 17731 16632 17740
rect 16580 17697 16589 17731
rect 16589 17697 16623 17731
rect 16623 17697 16632 17731
rect 16580 17688 16632 17697
rect 18604 17688 18656 17740
rect 10876 17663 10928 17672
rect 10876 17629 10885 17663
rect 10885 17629 10919 17663
rect 10919 17629 10928 17663
rect 10876 17620 10928 17629
rect 8300 17552 8352 17604
rect 9864 17595 9916 17604
rect 9864 17561 9873 17595
rect 9873 17561 9907 17595
rect 9907 17561 9916 17595
rect 9864 17552 9916 17561
rect 11980 17595 12032 17604
rect 11980 17561 11989 17595
rect 11989 17561 12023 17595
rect 12023 17561 12032 17595
rect 11980 17552 12032 17561
rect 12532 17595 12584 17604
rect 12532 17561 12541 17595
rect 12541 17561 12575 17595
rect 12575 17561 12584 17595
rect 12532 17552 12584 17561
rect 4620 17527 4672 17536
rect 4620 17493 4629 17527
rect 4629 17493 4663 17527
rect 4663 17493 4672 17527
rect 4620 17484 4672 17493
rect 5448 17484 5500 17536
rect 11796 17484 11848 17536
rect 13820 17620 13872 17672
rect 15016 17620 15068 17672
rect 16672 17620 16724 17672
rect 14648 17484 14700 17536
rect 19248 17484 19300 17536
rect 19984 17552 20036 17604
rect 24860 17688 24912 17740
rect 28080 17688 28132 17740
rect 22468 17663 22520 17672
rect 22468 17629 22477 17663
rect 22477 17629 22511 17663
rect 22511 17629 22520 17663
rect 22468 17620 22520 17629
rect 24216 17552 24268 17604
rect 27620 17620 27672 17672
rect 29092 17620 29144 17672
rect 31024 17663 31076 17672
rect 31024 17629 31033 17663
rect 31033 17629 31067 17663
rect 31067 17629 31076 17663
rect 31024 17620 31076 17629
rect 31208 17552 31260 17604
rect 23480 17484 23532 17536
rect 25872 17484 25924 17536
rect 30380 17484 30432 17536
rect 32404 17484 32456 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 3240 17280 3292 17332
rect 4620 17212 4672 17264
rect 7104 17280 7156 17332
rect 10876 17280 10928 17332
rect 17040 17280 17092 17332
rect 18696 17280 18748 17332
rect 19248 17280 19300 17332
rect 20352 17280 20404 17332
rect 8300 17212 8352 17264
rect 9036 17212 9088 17264
rect 3884 17187 3936 17196
rect 3884 17153 3893 17187
rect 3893 17153 3927 17187
rect 3927 17153 3936 17187
rect 3884 17144 3936 17153
rect 4712 17187 4764 17196
rect 4712 17153 4721 17187
rect 4721 17153 4755 17187
rect 4755 17153 4764 17187
rect 4712 17144 4764 17153
rect 5356 17187 5408 17196
rect 5356 17153 5365 17187
rect 5365 17153 5399 17187
rect 5399 17153 5408 17187
rect 5356 17144 5408 17153
rect 6000 17144 6052 17196
rect 2044 17076 2096 17128
rect 3332 17076 3384 17128
rect 8392 17144 8444 17196
rect 6552 17008 6604 17060
rect 6828 16940 6880 16992
rect 12624 17212 12676 17264
rect 14832 17212 14884 17264
rect 17868 17212 17920 17264
rect 12348 17187 12400 17196
rect 12348 17153 12357 17187
rect 12357 17153 12391 17187
rect 12391 17153 12400 17187
rect 12348 17144 12400 17153
rect 12992 17187 13044 17196
rect 12992 17153 13001 17187
rect 13001 17153 13035 17187
rect 13035 17153 13044 17187
rect 12992 17144 13044 17153
rect 14556 17144 14608 17196
rect 18696 17187 18748 17196
rect 18696 17153 18705 17187
rect 18705 17153 18739 17187
rect 18739 17153 18748 17187
rect 18696 17144 18748 17153
rect 8024 17008 8076 17060
rect 9864 17076 9916 17128
rect 16672 17008 16724 17060
rect 8300 16940 8352 16992
rect 8392 16940 8444 16992
rect 10232 16940 10284 16992
rect 10876 16940 10928 16992
rect 11888 16940 11940 16992
rect 15108 16940 15160 16992
rect 21456 17280 21508 17332
rect 23572 17280 23624 17332
rect 25136 17280 25188 17332
rect 20720 17212 20772 17264
rect 21364 17212 21416 17264
rect 23664 17212 23716 17264
rect 27252 17255 27304 17264
rect 27252 17221 27261 17255
rect 27261 17221 27295 17255
rect 27295 17221 27304 17255
rect 27252 17212 27304 17221
rect 32404 17255 32456 17264
rect 32404 17221 32413 17255
rect 32413 17221 32447 17255
rect 32447 17221 32456 17255
rect 32404 17212 32456 17221
rect 32496 17255 32548 17264
rect 32496 17221 32505 17255
rect 32505 17221 32539 17255
rect 32539 17221 32548 17255
rect 32496 17212 32548 17221
rect 38292 17187 38344 17196
rect 38292 17153 38301 17187
rect 38301 17153 38335 17187
rect 38335 17153 38344 17187
rect 38292 17144 38344 17153
rect 17868 17008 17920 17060
rect 27896 17076 27948 17128
rect 30196 17119 30248 17128
rect 30196 17085 30205 17119
rect 30205 17085 30239 17119
rect 30239 17085 30248 17119
rect 30196 17076 30248 17085
rect 32220 17076 32272 17128
rect 32588 17076 32640 17128
rect 23848 17051 23900 17060
rect 21364 16940 21416 16992
rect 21456 16940 21508 16992
rect 22836 16940 22888 16992
rect 23848 17017 23857 17051
rect 23857 17017 23891 17051
rect 23891 17017 23900 17051
rect 23848 17008 23900 17017
rect 31116 17008 31168 17060
rect 30564 16940 30616 16992
rect 35900 16940 35952 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 2320 16779 2372 16788
rect 2320 16745 2329 16779
rect 2329 16745 2363 16779
rect 2363 16745 2372 16779
rect 2320 16736 2372 16745
rect 4712 16779 4764 16788
rect 4712 16745 4721 16779
rect 4721 16745 4755 16779
rect 4755 16745 4764 16779
rect 4712 16736 4764 16745
rect 5356 16779 5408 16788
rect 5356 16745 5365 16779
rect 5365 16745 5399 16779
rect 5399 16745 5408 16779
rect 5356 16736 5408 16745
rect 5632 16736 5684 16788
rect 3240 16575 3292 16584
rect 3240 16541 3249 16575
rect 3249 16541 3283 16575
rect 3283 16541 3292 16575
rect 3240 16532 3292 16541
rect 3332 16575 3384 16584
rect 3332 16541 3341 16575
rect 3341 16541 3375 16575
rect 3375 16541 3384 16575
rect 7932 16668 7984 16720
rect 3884 16600 3936 16652
rect 3332 16532 3384 16541
rect 4896 16575 4948 16584
rect 4896 16541 4905 16575
rect 4905 16541 4939 16575
rect 4939 16541 4948 16575
rect 4896 16532 4948 16541
rect 6368 16532 6420 16584
rect 8024 16600 8076 16652
rect 9036 16736 9088 16788
rect 12348 16736 12400 16788
rect 12624 16736 12676 16788
rect 12992 16668 13044 16720
rect 14372 16668 14424 16720
rect 14648 16668 14700 16720
rect 18696 16736 18748 16788
rect 20352 16736 20404 16788
rect 22468 16736 22520 16788
rect 23664 16779 23716 16788
rect 23664 16745 23673 16779
rect 23673 16745 23707 16779
rect 23707 16745 23716 16779
rect 23664 16736 23716 16745
rect 30564 16779 30616 16788
rect 30564 16745 30573 16779
rect 30573 16745 30607 16779
rect 30607 16745 30616 16779
rect 30564 16736 30616 16745
rect 32496 16736 32548 16788
rect 20720 16668 20772 16720
rect 7196 16575 7248 16584
rect 7196 16541 7205 16575
rect 7205 16541 7239 16575
rect 7239 16541 7248 16575
rect 7196 16532 7248 16541
rect 7380 16532 7432 16584
rect 16028 16600 16080 16652
rect 30196 16643 30248 16652
rect 12256 16575 12308 16584
rect 12256 16541 12265 16575
rect 12265 16541 12299 16575
rect 12299 16541 12308 16575
rect 12256 16532 12308 16541
rect 8116 16464 8168 16516
rect 14556 16464 14608 16516
rect 4712 16396 4764 16448
rect 9404 16396 9456 16448
rect 9496 16396 9548 16448
rect 15660 16396 15712 16448
rect 17408 16396 17460 16448
rect 17960 16575 18012 16584
rect 17960 16541 17969 16575
rect 17969 16541 18003 16575
rect 18003 16541 18012 16575
rect 18696 16575 18748 16584
rect 17960 16532 18012 16541
rect 18696 16541 18705 16575
rect 18705 16541 18739 16575
rect 18739 16541 18748 16575
rect 18696 16532 18748 16541
rect 30196 16609 30205 16643
rect 30205 16609 30239 16643
rect 30239 16609 30248 16643
rect 30196 16600 30248 16609
rect 30380 16643 30432 16652
rect 30380 16609 30389 16643
rect 30389 16609 30423 16643
rect 30423 16609 30432 16643
rect 30380 16600 30432 16609
rect 20628 16532 20680 16584
rect 23296 16532 23348 16584
rect 33232 16575 33284 16584
rect 18052 16464 18104 16516
rect 21364 16464 21416 16516
rect 17960 16396 18012 16448
rect 18420 16396 18472 16448
rect 20904 16396 20956 16448
rect 25688 16464 25740 16516
rect 27344 16396 27396 16448
rect 33232 16541 33241 16575
rect 33241 16541 33275 16575
rect 33275 16541 33284 16575
rect 33232 16532 33284 16541
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 4804 16235 4856 16244
rect 4804 16201 4813 16235
rect 4813 16201 4847 16235
rect 4847 16201 4856 16235
rect 4804 16192 4856 16201
rect 6276 16192 6328 16244
rect 8576 16192 8628 16244
rect 1584 16099 1636 16108
rect 1584 16065 1593 16099
rect 1593 16065 1627 16099
rect 1627 16065 1636 16099
rect 1584 16056 1636 16065
rect 8668 16124 8720 16176
rect 10508 16167 10560 16176
rect 10508 16133 10517 16167
rect 10517 16133 10551 16167
rect 10551 16133 10560 16167
rect 10508 16124 10560 16133
rect 11152 16124 11204 16176
rect 5724 16099 5776 16108
rect 5724 16065 5733 16099
rect 5733 16065 5767 16099
rect 5767 16065 5776 16099
rect 5724 16056 5776 16065
rect 6368 16056 6420 16108
rect 10324 16056 10376 16108
rect 11336 16192 11388 16244
rect 12624 16124 12676 16176
rect 18696 16124 18748 16176
rect 17960 16056 18012 16108
rect 19800 16056 19852 16108
rect 20168 16235 20220 16244
rect 20168 16201 20177 16235
rect 20177 16201 20211 16235
rect 20211 16201 20220 16235
rect 23296 16235 23348 16244
rect 20168 16192 20220 16201
rect 23296 16201 23305 16235
rect 23305 16201 23339 16235
rect 23339 16201 23348 16235
rect 23296 16192 23348 16201
rect 22284 16124 22336 16176
rect 30564 16192 30616 16244
rect 20444 16056 20496 16108
rect 20720 16056 20772 16108
rect 21180 16056 21232 16108
rect 7380 15988 7432 16040
rect 10968 15988 11020 16040
rect 17592 15988 17644 16040
rect 17868 15988 17920 16040
rect 18696 16031 18748 16040
rect 6276 15920 6328 15972
rect 9496 15920 9548 15972
rect 1768 15895 1820 15904
rect 1768 15861 1777 15895
rect 1777 15861 1811 15895
rect 1811 15861 1820 15895
rect 1768 15852 1820 15861
rect 2872 15895 2924 15904
rect 2872 15861 2881 15895
rect 2881 15861 2915 15895
rect 2915 15861 2924 15895
rect 2872 15852 2924 15861
rect 6736 15852 6788 15904
rect 12440 15920 12492 15972
rect 17960 15920 18012 15972
rect 18696 15997 18705 16031
rect 18705 15997 18739 16031
rect 18739 15997 18748 16031
rect 18696 15988 18748 15997
rect 18788 15988 18840 16040
rect 23572 16056 23624 16108
rect 28540 16167 28592 16176
rect 28540 16133 28549 16167
rect 28549 16133 28583 16167
rect 28583 16133 28592 16167
rect 28540 16124 28592 16133
rect 27344 16099 27396 16108
rect 27344 16065 27353 16099
rect 27353 16065 27387 16099
rect 27387 16065 27396 16099
rect 27344 16056 27396 16065
rect 23940 15988 23992 16040
rect 25504 16031 25556 16040
rect 25504 15997 25513 16031
rect 25513 15997 25547 16031
rect 25547 15997 25556 16031
rect 25504 15988 25556 15997
rect 25964 16031 26016 16040
rect 25964 15997 25973 16031
rect 25973 15997 26007 16031
rect 26007 15997 26016 16031
rect 25964 15988 26016 15997
rect 28632 15988 28684 16040
rect 29276 15988 29328 16040
rect 25780 15920 25832 15972
rect 10508 15852 10560 15904
rect 19248 15852 19300 15904
rect 20628 15852 20680 15904
rect 22560 15895 22612 15904
rect 22560 15861 22569 15895
rect 22569 15861 22603 15895
rect 22603 15861 22612 15895
rect 22560 15852 22612 15861
rect 31484 16099 31536 16108
rect 31484 16065 31493 16099
rect 31493 16065 31527 16099
rect 31527 16065 31536 16099
rect 31484 16056 31536 16065
rect 30380 16031 30432 16040
rect 30380 15997 30389 16031
rect 30389 15997 30423 16031
rect 30423 15997 30432 16031
rect 30380 15988 30432 15997
rect 30012 15852 30064 15904
rect 33508 15852 33560 15904
rect 38200 15895 38252 15904
rect 38200 15861 38209 15895
rect 38209 15861 38243 15895
rect 38243 15861 38252 15895
rect 38200 15852 38252 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 8576 15648 8628 15700
rect 8668 15648 8720 15700
rect 11336 15648 11388 15700
rect 6276 15623 6328 15632
rect 6276 15589 6285 15623
rect 6285 15589 6319 15623
rect 6319 15589 6328 15623
rect 6276 15580 6328 15589
rect 10784 15580 10836 15632
rect 8760 15512 8812 15564
rect 12164 15512 12216 15564
rect 8116 15444 8168 15496
rect 10508 15444 10560 15496
rect 19984 15648 20036 15700
rect 20444 15648 20496 15700
rect 22744 15648 22796 15700
rect 20812 15580 20864 15632
rect 23664 15580 23716 15632
rect 30380 15648 30432 15700
rect 33508 15691 33560 15700
rect 33508 15657 33517 15691
rect 33517 15657 33551 15691
rect 33551 15657 33560 15691
rect 33508 15648 33560 15657
rect 14464 15512 14516 15564
rect 17868 15512 17920 15564
rect 23848 15555 23900 15564
rect 23848 15521 23857 15555
rect 23857 15521 23891 15555
rect 23891 15521 23900 15555
rect 23848 15512 23900 15521
rect 18696 15487 18748 15496
rect 18696 15453 18705 15487
rect 18705 15453 18739 15487
rect 18739 15453 18748 15487
rect 18696 15444 18748 15453
rect 20720 15444 20772 15496
rect 22468 15444 22520 15496
rect 25044 15487 25096 15496
rect 25044 15453 25053 15487
rect 25053 15453 25087 15487
rect 25087 15453 25096 15487
rect 25044 15444 25096 15453
rect 27528 15487 27580 15496
rect 5540 15308 5592 15360
rect 6460 15308 6512 15360
rect 6736 15376 6788 15428
rect 8668 15308 8720 15360
rect 11520 15376 11572 15428
rect 15660 15376 15712 15428
rect 17132 15376 17184 15428
rect 19340 15376 19392 15428
rect 22008 15376 22060 15428
rect 15016 15308 15068 15360
rect 15108 15308 15160 15360
rect 18696 15308 18748 15360
rect 20444 15351 20496 15360
rect 20444 15317 20453 15351
rect 20453 15317 20487 15351
rect 20487 15317 20496 15351
rect 20444 15308 20496 15317
rect 21916 15351 21968 15360
rect 21916 15317 21925 15351
rect 21925 15317 21959 15351
rect 21959 15317 21968 15351
rect 21916 15308 21968 15317
rect 23480 15419 23532 15428
rect 23480 15385 23489 15419
rect 23489 15385 23523 15419
rect 23523 15385 23532 15419
rect 27528 15453 27537 15487
rect 27537 15453 27571 15487
rect 27571 15453 27580 15487
rect 27528 15444 27580 15453
rect 31024 15512 31076 15564
rect 23480 15376 23532 15385
rect 23756 15308 23808 15360
rect 25780 15376 25832 15428
rect 26516 15376 26568 15428
rect 31208 15444 31260 15496
rect 35900 15512 35952 15564
rect 34612 15444 34664 15496
rect 30012 15419 30064 15428
rect 30012 15385 30021 15419
rect 30021 15385 30055 15419
rect 30055 15385 30064 15419
rect 30012 15376 30064 15385
rect 27344 15351 27396 15360
rect 27344 15317 27353 15351
rect 27353 15317 27387 15351
rect 27387 15317 27396 15351
rect 27344 15308 27396 15317
rect 27436 15308 27488 15360
rect 32864 15351 32916 15360
rect 32864 15317 32873 15351
rect 32873 15317 32907 15351
rect 32907 15317 32916 15351
rect 32864 15308 32916 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 13360 15104 13412 15156
rect 15568 15104 15620 15156
rect 16488 15104 16540 15156
rect 18696 15104 18748 15156
rect 20628 15104 20680 15156
rect 20720 15104 20772 15156
rect 23480 15104 23532 15156
rect 8576 15036 8628 15088
rect 10968 15036 11020 15088
rect 17592 15036 17644 15088
rect 20444 15036 20496 15088
rect 1768 15011 1820 15020
rect 1768 14977 1777 15011
rect 1777 14977 1811 15011
rect 1811 14977 1820 15011
rect 1768 14968 1820 14977
rect 4988 14968 5040 15020
rect 8760 15011 8812 15020
rect 8760 14977 8769 15011
rect 8769 14977 8803 15011
rect 8803 14977 8812 15011
rect 8760 14968 8812 14977
rect 12164 15011 12216 15020
rect 12164 14977 12173 15011
rect 12173 14977 12207 15011
rect 12207 14977 12216 15011
rect 12164 14968 12216 14977
rect 14464 15011 14516 15020
rect 3516 14900 3568 14952
rect 5356 14943 5408 14952
rect 5356 14909 5365 14943
rect 5365 14909 5399 14943
rect 5399 14909 5408 14943
rect 5356 14900 5408 14909
rect 12440 14943 12492 14952
rect 12440 14909 12449 14943
rect 12449 14909 12483 14943
rect 12483 14909 12492 14943
rect 12440 14900 12492 14909
rect 14464 14977 14473 15011
rect 14473 14977 14507 15011
rect 14507 14977 14516 15011
rect 14464 14968 14516 14977
rect 17868 14968 17920 15020
rect 21824 14968 21876 15020
rect 22468 14968 22520 15020
rect 23480 14968 23532 15020
rect 24860 14968 24912 15020
rect 27988 15036 28040 15088
rect 29460 15011 29512 15020
rect 29460 14977 29469 15011
rect 29469 14977 29503 15011
rect 29503 14977 29512 15011
rect 29460 14968 29512 14977
rect 14280 14900 14332 14952
rect 5080 14764 5132 14816
rect 5356 14764 5408 14816
rect 5632 14764 5684 14816
rect 13820 14764 13872 14816
rect 19432 14900 19484 14952
rect 20168 14943 20220 14952
rect 20168 14909 20177 14943
rect 20177 14909 20211 14943
rect 20211 14909 20220 14943
rect 20168 14900 20220 14909
rect 29000 14900 29052 14952
rect 16212 14875 16264 14884
rect 16212 14841 16221 14875
rect 16221 14841 16255 14875
rect 16255 14841 16264 14875
rect 16212 14832 16264 14841
rect 19524 14832 19576 14884
rect 25320 14832 25372 14884
rect 18144 14764 18196 14816
rect 18512 14764 18564 14816
rect 25228 14764 25280 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 5632 14560 5684 14612
rect 5908 14560 5960 14612
rect 11152 14560 11204 14612
rect 12440 14560 12492 14612
rect 12624 14560 12676 14612
rect 13452 14560 13504 14612
rect 18144 14560 18196 14612
rect 19524 14560 19576 14612
rect 19984 14560 20036 14612
rect 23756 14560 23808 14612
rect 27528 14560 27580 14612
rect 29460 14560 29512 14612
rect 34612 14560 34664 14612
rect 26424 14492 26476 14544
rect 13728 14424 13780 14476
rect 14464 14424 14516 14476
rect 17868 14424 17920 14476
rect 2872 14356 2924 14408
rect 10324 14356 10376 14408
rect 13360 14356 13412 14408
rect 15752 14356 15804 14408
rect 17500 14356 17552 14408
rect 20444 14356 20496 14408
rect 22468 14424 22520 14476
rect 22836 14467 22888 14476
rect 22836 14433 22845 14467
rect 22845 14433 22879 14467
rect 22879 14433 22888 14467
rect 22836 14424 22888 14433
rect 23664 14424 23716 14476
rect 21824 14356 21876 14408
rect 23204 14356 23256 14408
rect 25044 14356 25096 14408
rect 25596 14356 25648 14408
rect 32864 14424 32916 14476
rect 27804 14356 27856 14408
rect 38292 14399 38344 14408
rect 38292 14365 38301 14399
rect 38301 14365 38335 14399
rect 38335 14365 38344 14399
rect 38292 14356 38344 14365
rect 7472 14288 7524 14340
rect 12256 14288 12308 14340
rect 1492 14220 1544 14272
rect 21916 14288 21968 14340
rect 31760 14288 31812 14340
rect 31944 14331 31996 14340
rect 31944 14297 31953 14331
rect 31953 14297 31987 14331
rect 31987 14297 31996 14331
rect 31944 14288 31996 14297
rect 17132 14220 17184 14272
rect 17592 14263 17644 14272
rect 17592 14229 17601 14263
rect 17601 14229 17635 14263
rect 17635 14229 17644 14263
rect 17592 14220 17644 14229
rect 17776 14220 17828 14272
rect 20168 14220 20220 14272
rect 20628 14220 20680 14272
rect 24032 14220 24084 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 1584 14016 1636 14068
rect 3424 14016 3476 14068
rect 5172 13948 5224 14000
rect 5908 13948 5960 14000
rect 6184 13948 6236 14000
rect 1952 13923 2004 13932
rect 1952 13889 1961 13923
rect 1961 13889 1995 13923
rect 1995 13889 2004 13923
rect 1952 13880 2004 13889
rect 2412 13923 2464 13932
rect 2412 13889 2421 13923
rect 2421 13889 2455 13923
rect 2455 13889 2464 13923
rect 2412 13880 2464 13889
rect 8760 14016 8812 14068
rect 20720 14016 20772 14068
rect 20812 14016 20864 14068
rect 23756 14016 23808 14068
rect 25504 14016 25556 14068
rect 31024 14059 31076 14068
rect 31024 14025 31033 14059
rect 31033 14025 31067 14059
rect 31067 14025 31076 14059
rect 31024 14016 31076 14025
rect 13728 13948 13780 14000
rect 18512 13948 18564 14000
rect 20628 13948 20680 14000
rect 15752 13880 15804 13932
rect 17776 13880 17828 13932
rect 17868 13880 17920 13932
rect 20352 13923 20404 13932
rect 20352 13889 20361 13923
rect 20361 13889 20395 13923
rect 20395 13889 20404 13923
rect 20352 13880 20404 13889
rect 20444 13880 20496 13932
rect 3516 13855 3568 13864
rect 3516 13821 3525 13855
rect 3525 13821 3559 13855
rect 3559 13821 3568 13855
rect 3516 13812 3568 13821
rect 3792 13855 3844 13864
rect 3792 13821 3801 13855
rect 3801 13821 3835 13855
rect 3835 13821 3844 13855
rect 3792 13812 3844 13821
rect 13176 13812 13228 13864
rect 13452 13812 13504 13864
rect 3976 13676 4028 13728
rect 11428 13744 11480 13796
rect 13544 13744 13596 13796
rect 17960 13812 18012 13864
rect 10140 13676 10192 13728
rect 13636 13676 13688 13728
rect 14004 13676 14056 13728
rect 15016 13676 15068 13728
rect 17592 13744 17644 13796
rect 20996 13744 21048 13796
rect 19064 13676 19116 13728
rect 21364 13812 21416 13864
rect 21732 13880 21784 13932
rect 22744 13880 22796 13932
rect 24032 13923 24084 13932
rect 24032 13889 24041 13923
rect 24041 13889 24075 13923
rect 24075 13889 24084 13923
rect 24032 13880 24084 13889
rect 25228 13923 25280 13932
rect 25228 13889 25237 13923
rect 25237 13889 25271 13923
rect 25271 13889 25280 13923
rect 25228 13880 25280 13889
rect 27712 13948 27764 14000
rect 28448 13991 28500 14000
rect 28448 13957 28457 13991
rect 28457 13957 28491 13991
rect 28491 13957 28500 13991
rect 28448 13948 28500 13957
rect 27344 13923 27396 13932
rect 27344 13889 27353 13923
rect 27353 13889 27387 13923
rect 27387 13889 27396 13923
rect 27344 13880 27396 13889
rect 38108 13880 38160 13932
rect 25044 13855 25096 13864
rect 25044 13821 25053 13855
rect 25053 13821 25087 13855
rect 25087 13821 25096 13855
rect 25044 13812 25096 13821
rect 27068 13812 27120 13864
rect 28356 13855 28408 13864
rect 28356 13821 28365 13855
rect 28365 13821 28399 13855
rect 28399 13821 28408 13855
rect 28356 13812 28408 13821
rect 29000 13812 29052 13864
rect 30196 13812 30248 13864
rect 21364 13676 21416 13728
rect 21456 13676 21508 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 4896 13472 4948 13524
rect 6736 13472 6788 13524
rect 13544 13472 13596 13524
rect 13820 13472 13872 13524
rect 14556 13515 14608 13524
rect 14556 13481 14580 13515
rect 14580 13481 14608 13515
rect 14556 13472 14608 13481
rect 15660 13472 15712 13524
rect 20996 13472 21048 13524
rect 12716 13404 12768 13456
rect 3884 13336 3936 13388
rect 10140 13336 10192 13388
rect 12072 13336 12124 13388
rect 13728 13336 13780 13388
rect 15568 13404 15620 13456
rect 26240 13404 26292 13456
rect 28540 13472 28592 13524
rect 31760 13472 31812 13524
rect 29184 13404 29236 13456
rect 30472 13404 30524 13456
rect 31208 13404 31260 13456
rect 21456 13336 21508 13388
rect 21548 13336 21600 13388
rect 25044 13336 25096 13388
rect 31852 13336 31904 13388
rect 1584 13268 1636 13320
rect 3976 13311 4028 13320
rect 3976 13277 3985 13311
rect 3985 13277 4019 13311
rect 4019 13277 4028 13311
rect 3976 13268 4028 13277
rect 7748 13268 7800 13320
rect 9128 13311 9180 13320
rect 9128 13277 9137 13311
rect 9137 13277 9171 13311
rect 9171 13277 9180 13311
rect 9128 13268 9180 13277
rect 12624 13268 12676 13320
rect 14188 13268 14240 13320
rect 18696 13268 18748 13320
rect 21364 13268 21416 13320
rect 6460 13132 6512 13184
rect 10784 13200 10836 13252
rect 12716 13132 12768 13184
rect 12900 13132 12952 13184
rect 21548 13200 21600 13252
rect 22008 13268 22060 13320
rect 27436 13268 27488 13320
rect 29644 13268 29696 13320
rect 29920 13311 29972 13320
rect 29920 13277 29929 13311
rect 29929 13277 29963 13311
rect 29963 13277 29972 13311
rect 29920 13268 29972 13277
rect 32128 13311 32180 13320
rect 32128 13277 32137 13311
rect 32137 13277 32171 13311
rect 32171 13277 32180 13311
rect 32128 13268 32180 13277
rect 22744 13200 22796 13252
rect 30656 13243 30708 13252
rect 30656 13209 30665 13243
rect 30665 13209 30699 13243
rect 30699 13209 30708 13243
rect 30656 13200 30708 13209
rect 16028 13175 16080 13184
rect 16028 13141 16037 13175
rect 16037 13141 16071 13175
rect 16071 13141 16080 13175
rect 16028 13132 16080 13141
rect 17500 13132 17552 13184
rect 19248 13132 19300 13184
rect 19340 13132 19392 13184
rect 21640 13132 21692 13184
rect 21916 13132 21968 13184
rect 22008 13132 22060 13184
rect 30932 13132 30984 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 1584 12971 1636 12980
rect 1584 12937 1593 12971
rect 1593 12937 1627 12971
rect 1627 12937 1636 12971
rect 1584 12928 1636 12937
rect 3792 12928 3844 12980
rect 6828 12903 6880 12912
rect 6828 12869 6837 12903
rect 6837 12869 6871 12903
rect 6871 12869 6880 12903
rect 6828 12860 6880 12869
rect 7380 12903 7432 12912
rect 7380 12869 7389 12903
rect 7389 12869 7423 12903
rect 7423 12869 7432 12903
rect 7380 12860 7432 12869
rect 9404 12860 9456 12912
rect 12164 12928 12216 12980
rect 12900 12928 12952 12980
rect 12624 12860 12676 12912
rect 14280 12903 14332 12912
rect 14280 12869 14289 12903
rect 14289 12869 14323 12903
rect 14323 12869 14332 12903
rect 14280 12860 14332 12869
rect 1768 12835 1820 12844
rect 1768 12801 1777 12835
rect 1777 12801 1811 12835
rect 1811 12801 1820 12835
rect 1768 12792 1820 12801
rect 8668 12835 8720 12844
rect 8668 12801 8677 12835
rect 8677 12801 8711 12835
rect 8711 12801 8720 12835
rect 8668 12792 8720 12801
rect 10232 12792 10284 12844
rect 10600 12792 10652 12844
rect 12072 12792 12124 12844
rect 15660 12792 15712 12844
rect 4620 12724 4672 12776
rect 1860 12656 1912 12708
rect 9036 12724 9088 12776
rect 11060 12724 11112 12776
rect 3884 12588 3936 12640
rect 9036 12588 9088 12640
rect 9128 12588 9180 12640
rect 11612 12588 11664 12640
rect 11704 12588 11756 12640
rect 15568 12724 15620 12776
rect 17868 12928 17920 12980
rect 19156 12971 19208 12980
rect 19156 12937 19165 12971
rect 19165 12937 19199 12971
rect 19199 12937 19208 12971
rect 19156 12928 19208 12937
rect 19248 12928 19300 12980
rect 17316 12792 17368 12844
rect 21088 12835 21140 12844
rect 21088 12801 21097 12835
rect 21097 12801 21131 12835
rect 21131 12801 21140 12835
rect 21088 12792 21140 12801
rect 21732 12792 21784 12844
rect 21824 12792 21876 12844
rect 25504 12928 25556 12980
rect 28448 12928 28500 12980
rect 25412 12860 25464 12912
rect 30932 12903 30984 12912
rect 30932 12869 30941 12903
rect 30941 12869 30975 12903
rect 30975 12869 30984 12903
rect 30932 12860 30984 12869
rect 26608 12792 26660 12844
rect 27804 12835 27856 12844
rect 27804 12801 27813 12835
rect 27813 12801 27847 12835
rect 27847 12801 27856 12835
rect 27804 12792 27856 12801
rect 27896 12792 27948 12844
rect 36728 12792 36780 12844
rect 14188 12656 14240 12708
rect 16212 12656 16264 12708
rect 18696 12656 18748 12708
rect 12624 12588 12676 12640
rect 15384 12588 15436 12640
rect 16488 12588 16540 12640
rect 17776 12588 17828 12640
rect 22192 12656 22244 12708
rect 22560 12724 22612 12776
rect 24952 12724 25004 12776
rect 30840 12767 30892 12776
rect 30840 12733 30849 12767
rect 30849 12733 30883 12767
rect 30883 12733 30892 12767
rect 30840 12724 30892 12733
rect 31116 12767 31168 12776
rect 31116 12733 31125 12767
rect 31125 12733 31159 12767
rect 31159 12733 31168 12767
rect 31116 12724 31168 12733
rect 31300 12724 31352 12776
rect 29920 12656 29972 12708
rect 38200 12631 38252 12640
rect 38200 12597 38209 12631
rect 38209 12597 38243 12631
rect 38243 12597 38252 12631
rect 38200 12588 38252 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 1952 12427 2004 12436
rect 1952 12393 1961 12427
rect 1961 12393 1995 12427
rect 1995 12393 2004 12427
rect 1952 12384 2004 12393
rect 7380 12384 7432 12436
rect 10508 12384 10560 12436
rect 17040 12384 17092 12436
rect 3976 12223 4028 12232
rect 3976 12189 3985 12223
rect 3985 12189 4019 12223
rect 4019 12189 4028 12223
rect 3976 12180 4028 12189
rect 5632 12248 5684 12300
rect 6368 12248 6420 12300
rect 9220 12248 9272 12300
rect 11060 12248 11112 12300
rect 12256 12291 12308 12300
rect 12256 12257 12265 12291
rect 12265 12257 12299 12291
rect 12299 12257 12308 12291
rect 12256 12248 12308 12257
rect 21364 12384 21416 12436
rect 24952 12427 25004 12436
rect 24952 12393 24961 12427
rect 24961 12393 24995 12427
rect 24995 12393 25004 12427
rect 24952 12384 25004 12393
rect 30656 12384 30708 12436
rect 32128 12384 32180 12436
rect 36728 12384 36780 12436
rect 17224 12316 17276 12368
rect 23296 12316 23348 12368
rect 26332 12359 26384 12368
rect 26332 12325 26341 12359
rect 26341 12325 26375 12359
rect 26375 12325 26384 12359
rect 26332 12316 26384 12325
rect 27068 12316 27120 12368
rect 31944 12316 31996 12368
rect 5816 12180 5868 12232
rect 6276 12180 6328 12232
rect 7196 12180 7248 12232
rect 9128 12112 9180 12164
rect 11244 12112 11296 12164
rect 6184 12044 6236 12096
rect 11520 12044 11572 12096
rect 14372 12180 14424 12232
rect 21824 12180 21876 12232
rect 11888 12155 11940 12164
rect 11888 12121 11897 12155
rect 11897 12121 11931 12155
rect 11931 12121 11940 12155
rect 11888 12112 11940 12121
rect 14556 12112 14608 12164
rect 21456 12112 21508 12164
rect 21548 12112 21600 12164
rect 24860 12223 24912 12232
rect 24860 12189 24869 12223
rect 24869 12189 24903 12223
rect 24903 12189 24912 12223
rect 24860 12180 24912 12189
rect 25504 12180 25556 12232
rect 26700 12180 26752 12232
rect 30840 12248 30892 12300
rect 33232 12248 33284 12300
rect 31852 12223 31904 12232
rect 22744 12112 22796 12164
rect 27712 12155 27764 12164
rect 27712 12121 27721 12155
rect 27721 12121 27755 12155
rect 27755 12121 27764 12155
rect 27712 12112 27764 12121
rect 28080 12112 28132 12164
rect 28724 12112 28776 12164
rect 31852 12189 31861 12223
rect 31861 12189 31895 12223
rect 31895 12189 31904 12223
rect 31852 12180 31904 12189
rect 32680 12180 32732 12232
rect 17224 12044 17276 12096
rect 20904 12044 20956 12096
rect 21088 12044 21140 12096
rect 21916 12044 21968 12096
rect 29184 12044 29236 12096
rect 32404 12044 32456 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 6184 11840 6236 11892
rect 8300 11840 8352 11892
rect 9312 11840 9364 11892
rect 7932 11772 7984 11824
rect 10508 11772 10560 11824
rect 12624 11840 12676 11892
rect 13728 11840 13780 11892
rect 18144 11840 18196 11892
rect 11888 11772 11940 11824
rect 14740 11815 14792 11824
rect 14740 11781 14749 11815
rect 14749 11781 14783 11815
rect 14783 11781 14792 11815
rect 14740 11772 14792 11781
rect 17776 11772 17828 11824
rect 17040 11704 17092 11756
rect 20444 11840 20496 11892
rect 20996 11840 21048 11892
rect 21456 11840 21508 11892
rect 28724 11840 28776 11892
rect 22008 11772 22060 11824
rect 29184 11815 29236 11824
rect 29184 11781 29193 11815
rect 29193 11781 29227 11815
rect 29227 11781 29236 11815
rect 29184 11772 29236 11781
rect 32220 11772 32272 11824
rect 32404 11815 32456 11824
rect 32404 11781 32413 11815
rect 32413 11781 32447 11815
rect 32447 11781 32456 11815
rect 32404 11772 32456 11781
rect 32496 11815 32548 11824
rect 32496 11781 32505 11815
rect 32505 11781 32539 11815
rect 32539 11781 32548 11815
rect 32496 11772 32548 11781
rect 20352 11704 20404 11756
rect 20720 11704 20772 11756
rect 20812 11704 20864 11756
rect 3976 11636 4028 11688
rect 5172 11636 5224 11688
rect 8300 11636 8352 11688
rect 9128 11679 9180 11688
rect 9128 11645 9137 11679
rect 9137 11645 9171 11679
rect 9171 11645 9180 11679
rect 9128 11636 9180 11645
rect 9220 11636 9272 11688
rect 17132 11636 17184 11688
rect 17316 11636 17368 11688
rect 8760 11568 8812 11620
rect 11152 11568 11204 11620
rect 21180 11636 21232 11688
rect 21548 11704 21600 11756
rect 25320 11747 25372 11756
rect 25320 11713 25329 11747
rect 25329 11713 25363 11747
rect 25363 11713 25372 11747
rect 25320 11704 25372 11713
rect 21732 11636 21784 11688
rect 29276 11636 29328 11688
rect 32680 11679 32732 11688
rect 32680 11645 32689 11679
rect 32689 11645 32723 11679
rect 32723 11645 32732 11679
rect 32680 11636 32732 11645
rect 8668 11500 8720 11552
rect 9128 11500 9180 11552
rect 9588 11500 9640 11552
rect 13728 11500 13780 11552
rect 22928 11568 22980 11620
rect 17040 11500 17092 11552
rect 23480 11500 23532 11552
rect 29092 11500 29144 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 5908 11296 5960 11348
rect 11428 11296 11480 11348
rect 1952 11228 2004 11280
rect 6184 11228 6236 11280
rect 7656 11228 7708 11280
rect 9588 11228 9640 11280
rect 20720 11296 20772 11348
rect 25412 11296 25464 11348
rect 26700 11339 26752 11348
rect 26700 11305 26709 11339
rect 26709 11305 26743 11339
rect 26743 11305 26752 11339
rect 26700 11296 26752 11305
rect 28080 11339 28132 11348
rect 28080 11305 28089 11339
rect 28089 11305 28123 11339
rect 28123 11305 28132 11339
rect 28080 11296 28132 11305
rect 32496 11296 32548 11348
rect 38108 11339 38160 11348
rect 38108 11305 38117 11339
rect 38117 11305 38151 11339
rect 38151 11305 38160 11339
rect 38108 11296 38160 11305
rect 1768 11135 1820 11144
rect 1768 11101 1777 11135
rect 1777 11101 1811 11135
rect 1811 11101 1820 11135
rect 1768 11092 1820 11101
rect 3976 11092 4028 11144
rect 11060 11160 11112 11212
rect 11152 11160 11204 11212
rect 17040 11160 17092 11212
rect 17776 11160 17828 11212
rect 5632 11092 5684 11144
rect 6184 11092 6236 11144
rect 8760 11092 8812 11144
rect 9128 11092 9180 11144
rect 9312 11024 9364 11076
rect 16580 11092 16632 11144
rect 17132 11135 17184 11144
rect 17132 11101 17141 11135
rect 17141 11101 17175 11135
rect 17175 11101 17184 11135
rect 17132 11092 17184 11101
rect 18972 11160 19024 11212
rect 19984 11160 20036 11212
rect 21180 11092 21232 11144
rect 21548 11135 21600 11144
rect 21548 11101 21557 11135
rect 21557 11101 21591 11135
rect 21591 11101 21600 11135
rect 21548 11092 21600 11101
rect 6736 10956 6788 11008
rect 17316 11024 17368 11076
rect 20168 11024 20220 11076
rect 21640 11024 21692 11076
rect 23296 11135 23348 11144
rect 23296 11101 23305 11135
rect 23305 11101 23339 11135
rect 23339 11101 23348 11135
rect 23296 11092 23348 11101
rect 24676 11092 24728 11144
rect 25044 11092 25096 11144
rect 26516 11092 26568 11144
rect 31852 11160 31904 11212
rect 29092 11135 29144 11144
rect 29092 11101 29101 11135
rect 29101 11101 29135 11135
rect 29135 11101 29144 11135
rect 29092 11092 29144 11101
rect 31300 11092 31352 11144
rect 38292 11135 38344 11144
rect 38292 11101 38301 11135
rect 38301 11101 38335 11135
rect 38335 11101 38344 11135
rect 38292 11092 38344 11101
rect 33048 11024 33100 11076
rect 12256 10956 12308 11008
rect 14924 10956 14976 11008
rect 15108 10956 15160 11008
rect 21456 10956 21508 11008
rect 24768 10956 24820 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 6552 10752 6604 10804
rect 5448 10727 5500 10736
rect 5448 10693 5457 10727
rect 5457 10693 5491 10727
rect 5491 10693 5500 10727
rect 5448 10684 5500 10693
rect 6092 10684 6144 10736
rect 6736 10727 6788 10736
rect 6736 10693 6745 10727
rect 6745 10693 6779 10727
rect 6779 10693 6788 10727
rect 6736 10684 6788 10693
rect 7932 10752 7984 10804
rect 15016 10752 15068 10804
rect 20720 10752 20772 10804
rect 22468 10752 22520 10804
rect 25044 10795 25096 10804
rect 25044 10761 25053 10795
rect 25053 10761 25087 10795
rect 25087 10761 25096 10795
rect 25044 10752 25096 10761
rect 13176 10684 13228 10736
rect 1584 10616 1636 10668
rect 11336 10616 11388 10668
rect 12624 10659 12676 10668
rect 12624 10625 12633 10659
rect 12633 10625 12667 10659
rect 12667 10625 12676 10659
rect 12624 10616 12676 10625
rect 14004 10616 14056 10668
rect 7012 10591 7064 10600
rect 7012 10557 7021 10591
rect 7021 10557 7055 10591
rect 7055 10557 7064 10591
rect 7012 10548 7064 10557
rect 8392 10548 8444 10600
rect 17408 10684 17460 10736
rect 21916 10684 21968 10736
rect 22376 10684 22428 10736
rect 23664 10727 23716 10736
rect 23664 10693 23673 10727
rect 23673 10693 23707 10727
rect 23707 10693 23716 10727
rect 23664 10684 23716 10693
rect 20812 10659 20864 10668
rect 20812 10625 20821 10659
rect 20821 10625 20855 10659
rect 20855 10625 20864 10659
rect 20812 10616 20864 10625
rect 21548 10616 21600 10668
rect 25228 10659 25280 10668
rect 25228 10625 25237 10659
rect 25237 10625 25271 10659
rect 25271 10625 25280 10659
rect 25228 10616 25280 10625
rect 28724 10659 28776 10668
rect 28724 10625 28733 10659
rect 28733 10625 28767 10659
rect 28767 10625 28776 10659
rect 28724 10616 28776 10625
rect 29368 10659 29420 10668
rect 29368 10625 29377 10659
rect 29377 10625 29411 10659
rect 29411 10625 29420 10659
rect 29368 10616 29420 10625
rect 30104 10616 30156 10668
rect 33048 10616 33100 10668
rect 16580 10548 16632 10600
rect 19156 10548 19208 10600
rect 20904 10548 20956 10600
rect 22836 10548 22888 10600
rect 6644 10480 6696 10532
rect 9864 10480 9916 10532
rect 13636 10412 13688 10464
rect 14372 10455 14424 10464
rect 14372 10421 14381 10455
rect 14381 10421 14415 10455
rect 14415 10421 14424 10455
rect 14372 10412 14424 10421
rect 21272 10480 21324 10532
rect 29920 10548 29972 10600
rect 30380 10480 30432 10532
rect 21364 10412 21416 10464
rect 21456 10412 21508 10464
rect 23940 10412 23992 10464
rect 24032 10412 24084 10464
rect 27804 10412 27856 10464
rect 30012 10412 30064 10464
rect 30564 10412 30616 10464
rect 34796 10412 34848 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 4620 10208 4672 10260
rect 12164 10208 12216 10260
rect 14004 10208 14056 10260
rect 25228 10208 25280 10260
rect 29920 10208 29972 10260
rect 10876 10140 10928 10192
rect 15200 10140 15252 10192
rect 17316 10140 17368 10192
rect 5264 10072 5316 10124
rect 1768 10047 1820 10056
rect 1768 10013 1777 10047
rect 1777 10013 1811 10047
rect 1811 10013 1820 10047
rect 1768 10004 1820 10013
rect 3976 10047 4028 10056
rect 3976 10013 3985 10047
rect 3985 10013 4019 10047
rect 4019 10013 4028 10047
rect 3976 10004 4028 10013
rect 14372 10072 14424 10124
rect 14556 10072 14608 10124
rect 24032 10140 24084 10192
rect 24216 10140 24268 10192
rect 24952 10140 25004 10192
rect 22100 10115 22152 10124
rect 22100 10081 22109 10115
rect 22109 10081 22143 10115
rect 22143 10081 22152 10115
rect 22100 10072 22152 10081
rect 25044 10072 25096 10124
rect 5908 9936 5960 9988
rect 6092 9936 6144 9988
rect 1860 9868 1912 9920
rect 4896 9868 4948 9920
rect 12532 9936 12584 9988
rect 13636 9936 13688 9988
rect 14924 9936 14976 9988
rect 20076 9936 20128 9988
rect 20720 10004 20772 10056
rect 21548 9936 21600 9988
rect 22376 10004 22428 10056
rect 23940 10004 23992 10056
rect 30012 10047 30064 10056
rect 30012 10013 30021 10047
rect 30021 10013 30055 10047
rect 30055 10013 30064 10047
rect 30012 10004 30064 10013
rect 22744 9936 22796 9988
rect 24768 9979 24820 9988
rect 24768 9945 24777 9979
rect 24777 9945 24811 9979
rect 24811 9945 24820 9979
rect 24768 9936 24820 9945
rect 9312 9868 9364 9920
rect 22100 9868 22152 9920
rect 25136 9868 25188 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 8116 9528 8168 9580
rect 20444 9664 20496 9716
rect 19984 9596 20036 9648
rect 20168 9596 20220 9648
rect 6552 9460 6604 9512
rect 7656 9460 7708 9512
rect 10508 9528 10560 9580
rect 18144 9528 18196 9580
rect 8300 9460 8352 9512
rect 9128 9503 9180 9512
rect 9128 9469 9137 9503
rect 9137 9469 9171 9503
rect 9171 9469 9180 9503
rect 9128 9460 9180 9469
rect 8024 9392 8076 9444
rect 12256 9392 12308 9444
rect 13912 9392 13964 9444
rect 11980 9324 12032 9376
rect 14280 9324 14332 9376
rect 17960 9460 18012 9512
rect 19156 9460 19208 9512
rect 19248 9460 19300 9512
rect 20076 9528 20128 9580
rect 20444 9528 20496 9580
rect 21088 9596 21140 9648
rect 21364 9664 21416 9716
rect 22836 9664 22888 9716
rect 23664 9707 23716 9716
rect 23664 9673 23673 9707
rect 23673 9673 23707 9707
rect 23707 9673 23716 9707
rect 23664 9664 23716 9673
rect 20812 9528 20864 9580
rect 22008 9528 22060 9580
rect 22560 9571 22612 9580
rect 22560 9537 22569 9571
rect 22569 9537 22603 9571
rect 22603 9537 22612 9571
rect 22560 9528 22612 9537
rect 21916 9392 21968 9444
rect 24768 9528 24820 9580
rect 30564 9528 30616 9580
rect 25228 9460 25280 9512
rect 28724 9460 28776 9512
rect 20536 9324 20588 9376
rect 21088 9324 21140 9376
rect 21640 9324 21692 9376
rect 22008 9324 22060 9376
rect 37740 9392 37792 9444
rect 23480 9324 23532 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 7012 9120 7064 9172
rect 8024 9120 8076 9172
rect 8116 9120 8168 9172
rect 21088 9120 21140 9172
rect 21180 9120 21232 9172
rect 28724 9163 28776 9172
rect 8484 9052 8536 9104
rect 14464 9052 14516 9104
rect 18144 9052 18196 9104
rect 25228 9095 25280 9104
rect 25228 9061 25237 9095
rect 25237 9061 25271 9095
rect 25271 9061 25280 9095
rect 25228 9052 25280 9061
rect 6644 9027 6696 9036
rect 6644 8993 6653 9027
rect 6653 8993 6687 9027
rect 6687 8993 6696 9027
rect 6644 8984 6696 8993
rect 11888 8984 11940 9036
rect 12256 8984 12308 9036
rect 18604 9027 18656 9036
rect 1860 8959 1912 8968
rect 1860 8925 1869 8959
rect 1869 8925 1903 8959
rect 1903 8925 1912 8959
rect 1860 8916 1912 8925
rect 11336 8959 11388 8968
rect 11336 8925 11345 8959
rect 11345 8925 11379 8959
rect 11379 8925 11388 8959
rect 11336 8916 11388 8925
rect 11520 8916 11572 8968
rect 12440 8916 12492 8968
rect 16580 8959 16632 8968
rect 16580 8925 16589 8959
rect 16589 8925 16623 8959
rect 16623 8925 16632 8959
rect 16580 8916 16632 8925
rect 6000 8891 6052 8900
rect 6000 8857 6009 8891
rect 6009 8857 6043 8891
rect 6043 8857 6052 8891
rect 6000 8848 6052 8857
rect 6460 8848 6512 8900
rect 8116 8848 8168 8900
rect 11244 8848 11296 8900
rect 8576 8780 8628 8832
rect 11980 8780 12032 8832
rect 16856 8891 16908 8900
rect 16856 8857 16865 8891
rect 16865 8857 16899 8891
rect 16899 8857 16908 8891
rect 16856 8848 16908 8857
rect 17868 8780 17920 8832
rect 18604 8993 18613 9027
rect 18613 8993 18647 9027
rect 18647 8993 18656 9027
rect 18604 8984 18656 8993
rect 18236 8916 18288 8968
rect 19340 8916 19392 8968
rect 20168 8916 20220 8968
rect 20628 8916 20680 8968
rect 21640 8959 21692 8968
rect 21640 8925 21649 8959
rect 21649 8925 21683 8959
rect 21683 8925 21692 8959
rect 21640 8916 21692 8925
rect 21916 8916 21968 8968
rect 22560 8959 22612 8968
rect 22560 8925 22569 8959
rect 22569 8925 22603 8959
rect 22603 8925 22612 8959
rect 22560 8916 22612 8925
rect 23572 8916 23624 8968
rect 28724 9129 28733 9163
rect 28733 9129 28767 9163
rect 28767 9129 28776 9163
rect 28724 9120 28776 9129
rect 27988 8916 28040 8968
rect 28632 8959 28684 8968
rect 28632 8925 28641 8959
rect 28641 8925 28675 8959
rect 28675 8925 28684 8959
rect 28632 8916 28684 8925
rect 29368 8916 29420 8968
rect 30564 8959 30616 8968
rect 30564 8925 30573 8959
rect 30573 8925 30607 8959
rect 30607 8925 30616 8959
rect 30564 8916 30616 8925
rect 34796 8916 34848 8968
rect 22652 8848 22704 8900
rect 20076 8780 20128 8832
rect 20628 8823 20680 8832
rect 20628 8789 20637 8823
rect 20637 8789 20671 8823
rect 20671 8789 20680 8823
rect 20628 8780 20680 8789
rect 20720 8780 20772 8832
rect 21824 8780 21876 8832
rect 23756 8848 23808 8900
rect 24216 8780 24268 8832
rect 27160 8780 27212 8832
rect 28448 8780 28500 8832
rect 32496 8780 32548 8832
rect 38200 8823 38252 8832
rect 38200 8789 38209 8823
rect 38209 8789 38243 8823
rect 38243 8789 38252 8823
rect 38200 8780 38252 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 2044 8619 2096 8628
rect 2044 8585 2053 8619
rect 2053 8585 2087 8619
rect 2087 8585 2096 8619
rect 2044 8576 2096 8585
rect 8116 8508 8168 8560
rect 2320 8440 2372 8492
rect 6368 8440 6420 8492
rect 8300 8576 8352 8628
rect 9220 8576 9272 8628
rect 10140 8576 10192 8628
rect 10508 8576 10560 8628
rect 15476 8576 15528 8628
rect 8484 8551 8536 8560
rect 8484 8517 8493 8551
rect 8493 8517 8527 8551
rect 8527 8517 8536 8551
rect 8484 8508 8536 8517
rect 11980 8551 12032 8560
rect 11980 8517 11989 8551
rect 11989 8517 12023 8551
rect 12023 8517 12032 8551
rect 11980 8508 12032 8517
rect 15844 8508 15896 8560
rect 16856 8576 16908 8628
rect 18972 8576 19024 8628
rect 19708 8576 19760 8628
rect 20444 8576 20496 8628
rect 20904 8576 20956 8628
rect 21088 8619 21140 8628
rect 21088 8585 21097 8619
rect 21097 8585 21131 8619
rect 21131 8585 21140 8619
rect 21088 8576 21140 8585
rect 18236 8508 18288 8560
rect 19616 8508 19668 8560
rect 9588 8440 9640 8492
rect 5816 8372 5868 8424
rect 8576 8372 8628 8424
rect 19800 8440 19852 8492
rect 20352 8440 20404 8492
rect 20812 8440 20864 8492
rect 11336 8304 11388 8356
rect 17868 8372 17920 8424
rect 17960 8372 18012 8424
rect 13912 8304 13964 8356
rect 14464 8304 14516 8356
rect 16120 8304 16172 8356
rect 22192 8551 22244 8560
rect 22192 8517 22201 8551
rect 22201 8517 22235 8551
rect 22235 8517 22244 8551
rect 22192 8508 22244 8517
rect 22652 8508 22704 8560
rect 23388 8576 23440 8628
rect 23848 8576 23900 8628
rect 24860 8508 24912 8560
rect 23572 8483 23624 8492
rect 23572 8449 23581 8483
rect 23581 8449 23615 8483
rect 23615 8449 23624 8483
rect 23572 8440 23624 8449
rect 24032 8440 24084 8492
rect 25964 8508 26016 8560
rect 26148 8508 26200 8560
rect 26240 8508 26292 8560
rect 29368 8508 29420 8560
rect 27160 8483 27212 8492
rect 27160 8449 27169 8483
rect 27169 8449 27203 8483
rect 27203 8449 27212 8483
rect 27160 8440 27212 8449
rect 28448 8483 28500 8492
rect 28448 8449 28457 8483
rect 28457 8449 28491 8483
rect 28491 8449 28500 8483
rect 28448 8440 28500 8449
rect 30564 8551 30616 8560
rect 30564 8517 30573 8551
rect 30573 8517 30607 8551
rect 30607 8517 30616 8551
rect 30564 8508 30616 8517
rect 31208 8508 31260 8560
rect 24676 8415 24728 8424
rect 24676 8381 24685 8415
rect 24685 8381 24719 8415
rect 24719 8381 24728 8415
rect 24676 8372 24728 8381
rect 24860 8415 24912 8424
rect 24860 8381 24869 8415
rect 24869 8381 24903 8415
rect 24903 8381 24912 8415
rect 24860 8372 24912 8381
rect 26332 8372 26384 8424
rect 3976 8236 4028 8288
rect 11060 8236 11112 8288
rect 11796 8236 11848 8288
rect 13820 8236 13872 8288
rect 14004 8236 14056 8288
rect 19800 8279 19852 8288
rect 19800 8245 19809 8279
rect 19809 8245 19843 8279
rect 19843 8245 19852 8279
rect 20168 8304 20220 8356
rect 19800 8236 19852 8245
rect 21272 8236 21324 8288
rect 23572 8304 23624 8356
rect 25044 8347 25096 8356
rect 25044 8313 25053 8347
rect 25053 8313 25087 8347
rect 25087 8313 25096 8347
rect 25044 8304 25096 8313
rect 26516 8347 26568 8356
rect 26516 8313 26525 8347
rect 26525 8313 26559 8347
rect 26559 8313 26568 8347
rect 32496 8483 32548 8492
rect 32496 8449 32505 8483
rect 32505 8449 32539 8483
rect 32539 8449 32548 8483
rect 32496 8440 32548 8449
rect 31760 8372 31812 8424
rect 26516 8304 26568 8313
rect 34428 8304 34480 8356
rect 23664 8279 23716 8288
rect 23664 8245 23673 8279
rect 23673 8245 23707 8279
rect 23707 8245 23716 8279
rect 23664 8236 23716 8245
rect 28448 8236 28500 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 2412 8032 2464 8084
rect 5724 8075 5776 8084
rect 5724 8041 5733 8075
rect 5733 8041 5767 8075
rect 5767 8041 5776 8075
rect 5724 8032 5776 8041
rect 10048 8032 10100 8084
rect 10324 8032 10376 8084
rect 18696 8032 18748 8084
rect 19340 8032 19392 8084
rect 20076 8032 20128 8084
rect 22100 8032 22152 8084
rect 22468 8075 22520 8084
rect 6000 7896 6052 7948
rect 13728 7964 13780 8016
rect 11060 7896 11112 7948
rect 1860 7828 1912 7880
rect 2780 7871 2832 7880
rect 2780 7837 2789 7871
rect 2789 7837 2823 7871
rect 2823 7837 2832 7871
rect 3976 7871 4028 7880
rect 2780 7828 2832 7837
rect 3976 7837 3985 7871
rect 3985 7837 4019 7871
rect 4019 7837 4028 7871
rect 3976 7828 4028 7837
rect 6552 7871 6604 7880
rect 6552 7837 6561 7871
rect 6561 7837 6595 7871
rect 6595 7837 6604 7871
rect 6552 7828 6604 7837
rect 11152 7871 11204 7880
rect 11152 7837 11161 7871
rect 11161 7837 11195 7871
rect 11195 7837 11204 7871
rect 11152 7828 11204 7837
rect 17960 7896 18012 7948
rect 20812 7964 20864 8016
rect 20996 7964 21048 8016
rect 22468 8041 22477 8075
rect 22477 8041 22511 8075
rect 22511 8041 22520 8075
rect 22468 8032 22520 8041
rect 24860 8032 24912 8084
rect 26148 8032 26200 8084
rect 29644 8032 29696 8084
rect 30564 8032 30616 8084
rect 31760 8075 31812 8084
rect 31760 8041 31769 8075
rect 31769 8041 31803 8075
rect 31803 8041 31812 8075
rect 31760 8032 31812 8041
rect 22560 7964 22612 8016
rect 20720 7896 20772 7948
rect 28264 7964 28316 8016
rect 14280 7871 14332 7880
rect 14280 7837 14289 7871
rect 14289 7837 14323 7871
rect 14323 7837 14332 7871
rect 14280 7828 14332 7837
rect 18052 7828 18104 7880
rect 18696 7871 18748 7880
rect 18696 7837 18705 7871
rect 18705 7837 18739 7871
rect 18739 7837 18748 7871
rect 18696 7828 18748 7837
rect 21916 7828 21968 7880
rect 22008 7828 22060 7880
rect 22284 7828 22336 7880
rect 22468 7828 22520 7880
rect 4528 7760 4580 7812
rect 8484 7760 8536 7812
rect 11336 7760 11388 7812
rect 8668 7692 8720 7744
rect 10600 7692 10652 7744
rect 15200 7760 15252 7812
rect 18236 7760 18288 7812
rect 13820 7692 13872 7744
rect 18328 7692 18380 7744
rect 18512 7692 18564 7744
rect 19340 7760 19392 7812
rect 19616 7760 19668 7812
rect 19800 7760 19852 7812
rect 23664 7760 23716 7812
rect 23848 7871 23900 7880
rect 23848 7837 23857 7871
rect 23857 7837 23891 7871
rect 23891 7837 23900 7871
rect 24768 7871 24820 7880
rect 23848 7828 23900 7837
rect 24768 7837 24777 7871
rect 24777 7837 24811 7871
rect 24811 7837 24820 7871
rect 24768 7828 24820 7837
rect 28632 7939 28684 7948
rect 28632 7905 28641 7939
rect 28641 7905 28675 7939
rect 28675 7905 28684 7939
rect 28632 7896 28684 7905
rect 28448 7803 28500 7812
rect 28448 7769 28457 7803
rect 28457 7769 28491 7803
rect 28491 7769 28500 7803
rect 28448 7760 28500 7769
rect 28724 7760 28776 7812
rect 30380 7828 30432 7880
rect 33048 7828 33100 7880
rect 38292 7871 38344 7880
rect 38292 7837 38301 7871
rect 38301 7837 38335 7871
rect 38335 7837 38344 7871
rect 38292 7828 38344 7837
rect 22376 7692 22428 7744
rect 23572 7692 23624 7744
rect 27344 7692 27396 7744
rect 37280 7692 37332 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 6092 7488 6144 7540
rect 8208 7488 8260 7540
rect 8484 7488 8536 7540
rect 14004 7488 14056 7540
rect 6552 7420 6604 7472
rect 1676 7352 1728 7404
rect 9312 7420 9364 7472
rect 9404 7420 9456 7472
rect 13912 7420 13964 7472
rect 7840 7327 7892 7336
rect 7840 7293 7849 7327
rect 7849 7293 7883 7327
rect 7883 7293 7892 7327
rect 7840 7284 7892 7293
rect 9588 7284 9640 7336
rect 18328 7488 18380 7540
rect 14556 7463 14608 7472
rect 14556 7429 14565 7463
rect 14565 7429 14599 7463
rect 14599 7429 14608 7463
rect 14556 7420 14608 7429
rect 21456 7420 21508 7472
rect 23572 7420 23624 7472
rect 24400 7420 24452 7472
rect 29184 7463 29236 7472
rect 29184 7429 29193 7463
rect 29193 7429 29227 7463
rect 29227 7429 29236 7463
rect 29184 7420 29236 7429
rect 14280 7327 14332 7336
rect 14280 7293 14289 7327
rect 14289 7293 14323 7327
rect 14323 7293 14332 7327
rect 14280 7284 14332 7293
rect 13820 7216 13872 7268
rect 15108 7284 15160 7336
rect 15568 7284 15620 7336
rect 16304 7327 16356 7336
rect 16304 7293 16313 7327
rect 16313 7293 16347 7327
rect 16347 7293 16356 7327
rect 16304 7284 16356 7293
rect 17960 7327 18012 7336
rect 17960 7293 17969 7327
rect 17969 7293 18003 7327
rect 18003 7293 18012 7327
rect 17960 7284 18012 7293
rect 18236 7327 18288 7336
rect 18236 7293 18245 7327
rect 18245 7293 18279 7327
rect 18279 7293 18288 7327
rect 18236 7284 18288 7293
rect 18328 7284 18380 7336
rect 19892 7284 19944 7336
rect 21088 7352 21140 7404
rect 21732 7352 21784 7404
rect 22008 7395 22060 7404
rect 22008 7361 22017 7395
rect 22017 7361 22051 7395
rect 22051 7361 22060 7395
rect 22008 7352 22060 7361
rect 23664 7352 23716 7404
rect 24032 7352 24084 7404
rect 27344 7395 27396 7404
rect 27344 7361 27353 7395
rect 27353 7361 27387 7395
rect 27387 7361 27396 7395
rect 27344 7352 27396 7361
rect 30196 7395 30248 7404
rect 30196 7361 30205 7395
rect 30205 7361 30239 7395
rect 30239 7361 30248 7395
rect 30196 7352 30248 7361
rect 21640 7284 21692 7336
rect 11060 7148 11112 7200
rect 12072 7148 12124 7200
rect 23480 7216 23532 7268
rect 26516 7284 26568 7336
rect 29092 7327 29144 7336
rect 29092 7293 29101 7327
rect 29101 7293 29135 7327
rect 29135 7293 29144 7327
rect 29092 7284 29144 7293
rect 29368 7327 29420 7336
rect 29368 7293 29377 7327
rect 29377 7293 29411 7327
rect 29411 7293 29420 7327
rect 29368 7284 29420 7293
rect 27252 7216 27304 7268
rect 24768 7148 24820 7200
rect 31208 7148 31260 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 9404 6944 9456 6996
rect 19892 6944 19944 6996
rect 21640 6944 21692 6996
rect 21732 6944 21784 6996
rect 25596 6944 25648 6996
rect 11336 6876 11388 6928
rect 13820 6876 13872 6928
rect 13912 6876 13964 6928
rect 14648 6876 14700 6928
rect 16580 6876 16632 6928
rect 20628 6876 20680 6928
rect 21548 6919 21600 6928
rect 21548 6885 21557 6919
rect 21557 6885 21591 6919
rect 21591 6885 21600 6919
rect 21548 6876 21600 6885
rect 2872 6604 2924 6656
rect 6460 6808 6512 6860
rect 10508 6808 10560 6860
rect 11704 6808 11756 6860
rect 17224 6808 17276 6860
rect 23296 6876 23348 6928
rect 9220 6740 9272 6792
rect 11428 6740 11480 6792
rect 18236 6740 18288 6792
rect 19064 6740 19116 6792
rect 21916 6740 21968 6792
rect 29184 6808 29236 6860
rect 23204 6740 23256 6792
rect 23388 6740 23440 6792
rect 28724 6783 28776 6792
rect 28724 6749 28733 6783
rect 28733 6749 28767 6783
rect 28767 6749 28776 6783
rect 28724 6740 28776 6749
rect 9588 6672 9640 6724
rect 7840 6647 7892 6656
rect 7840 6613 7849 6647
rect 7849 6613 7883 6647
rect 7883 6613 7892 6647
rect 7840 6604 7892 6613
rect 7932 6604 7984 6656
rect 17224 6604 17276 6656
rect 17776 6604 17828 6656
rect 20812 6604 20864 6656
rect 22192 6604 22244 6656
rect 25688 6604 25740 6656
rect 25964 6604 26016 6656
rect 28908 6604 28960 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 7932 6400 7984 6452
rect 10416 6443 10468 6452
rect 10416 6409 10425 6443
rect 10425 6409 10459 6443
rect 10459 6409 10468 6443
rect 10416 6400 10468 6409
rect 10508 6400 10560 6452
rect 16580 6400 16632 6452
rect 16672 6400 16724 6452
rect 19340 6400 19392 6452
rect 19984 6443 20036 6452
rect 19984 6409 19993 6443
rect 19993 6409 20027 6443
rect 20027 6409 20036 6443
rect 19984 6400 20036 6409
rect 20260 6400 20312 6452
rect 23020 6400 23072 6452
rect 23204 6375 23256 6384
rect 23204 6341 23213 6375
rect 23213 6341 23247 6375
rect 23247 6341 23256 6375
rect 23204 6332 23256 6341
rect 23572 6332 23624 6384
rect 24124 6332 24176 6384
rect 25320 6375 25372 6384
rect 25320 6341 25329 6375
rect 25329 6341 25363 6375
rect 25363 6341 25372 6375
rect 25320 6332 25372 6341
rect 25964 6332 26016 6384
rect 30840 6400 30892 6452
rect 27620 6332 27672 6384
rect 28816 6332 28868 6384
rect 28908 6332 28960 6384
rect 30380 6332 30432 6384
rect 1952 6307 2004 6316
rect 1952 6273 1961 6307
rect 1961 6273 1995 6307
rect 1995 6273 2004 6307
rect 1952 6264 2004 6273
rect 5356 6264 5408 6316
rect 3976 6239 4028 6248
rect 3976 6205 3985 6239
rect 3985 6205 4019 6239
rect 4019 6205 4028 6239
rect 3976 6196 4028 6205
rect 5908 6196 5960 6248
rect 5724 6171 5776 6180
rect 5724 6137 5733 6171
rect 5733 6137 5767 6171
rect 5767 6137 5776 6171
rect 5724 6128 5776 6137
rect 7196 6128 7248 6180
rect 9496 6196 9548 6248
rect 9588 6196 9640 6248
rect 12808 6196 12860 6248
rect 15292 6196 15344 6248
rect 10692 6128 10744 6180
rect 16672 6128 16724 6180
rect 9128 6060 9180 6112
rect 9312 6060 9364 6112
rect 19248 6264 19300 6316
rect 19892 6307 19944 6316
rect 19892 6273 19901 6307
rect 19901 6273 19935 6307
rect 19935 6273 19944 6307
rect 19892 6264 19944 6273
rect 21456 6264 21508 6316
rect 22008 6307 22060 6316
rect 22008 6273 22017 6307
rect 22017 6273 22051 6307
rect 22051 6273 22060 6307
rect 22008 6264 22060 6273
rect 24216 6307 24268 6316
rect 24216 6273 24225 6307
rect 24225 6273 24259 6307
rect 24259 6273 24268 6307
rect 24216 6264 24268 6273
rect 30012 6264 30064 6316
rect 38292 6307 38344 6316
rect 38292 6273 38301 6307
rect 38301 6273 38335 6307
rect 38335 6273 38344 6307
rect 38292 6264 38344 6273
rect 20904 6196 20956 6248
rect 22928 6196 22980 6248
rect 21456 6128 21508 6180
rect 24952 6196 25004 6248
rect 28172 6196 28224 6248
rect 30656 6239 30708 6248
rect 24676 6128 24728 6180
rect 27804 6171 27856 6180
rect 27804 6137 27813 6171
rect 27813 6137 27847 6171
rect 27847 6137 27856 6171
rect 27804 6128 27856 6137
rect 28632 6128 28684 6180
rect 18604 6103 18656 6112
rect 18604 6069 18613 6103
rect 18613 6069 18647 6103
rect 18647 6069 18656 6103
rect 18604 6060 18656 6069
rect 18696 6060 18748 6112
rect 21180 6060 21232 6112
rect 21548 6060 21600 6112
rect 23020 6060 23072 6112
rect 30656 6205 30665 6239
rect 30665 6205 30699 6239
rect 30699 6205 30708 6239
rect 30656 6196 30708 6205
rect 38108 6103 38160 6112
rect 38108 6069 38117 6103
rect 38117 6069 38151 6103
rect 38151 6069 38160 6103
rect 38108 6060 38160 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 1584 5899 1636 5908
rect 1584 5865 1593 5899
rect 1593 5865 1627 5899
rect 1627 5865 1636 5899
rect 1584 5856 1636 5865
rect 6184 5856 6236 5908
rect 12164 5856 12216 5908
rect 16028 5856 16080 5908
rect 1768 5695 1820 5704
rect 1768 5661 1777 5695
rect 1777 5661 1811 5695
rect 1811 5661 1820 5695
rect 1768 5652 1820 5661
rect 3976 5695 4028 5704
rect 3976 5661 3985 5695
rect 3985 5661 4019 5695
rect 4019 5661 4028 5695
rect 3976 5652 4028 5661
rect 9312 5788 9364 5840
rect 8668 5720 8720 5772
rect 18604 5788 18656 5840
rect 21456 5788 21508 5840
rect 22100 5899 22152 5908
rect 22100 5865 22109 5899
rect 22109 5865 22143 5899
rect 22143 5865 22152 5899
rect 22100 5856 22152 5865
rect 20996 5720 21048 5772
rect 21640 5720 21692 5772
rect 23204 5856 23256 5908
rect 25872 5856 25924 5908
rect 27620 5899 27672 5908
rect 27620 5865 27629 5899
rect 27629 5865 27663 5899
rect 27663 5865 27672 5899
rect 27620 5856 27672 5865
rect 28816 5899 28868 5908
rect 28816 5865 28825 5899
rect 28825 5865 28859 5899
rect 28859 5865 28868 5899
rect 28816 5856 28868 5865
rect 30012 5899 30064 5908
rect 30012 5865 30021 5899
rect 30021 5865 30055 5899
rect 30055 5865 30064 5899
rect 30012 5856 30064 5865
rect 30656 5856 30708 5908
rect 23296 5788 23348 5840
rect 9220 5652 9272 5704
rect 11152 5652 11204 5704
rect 11612 5584 11664 5636
rect 11980 5584 12032 5636
rect 13636 5584 13688 5636
rect 14280 5584 14332 5636
rect 16304 5516 16356 5568
rect 17224 5516 17276 5568
rect 21732 5652 21784 5704
rect 22376 5652 22428 5704
rect 22652 5695 22704 5704
rect 22652 5661 22661 5695
rect 22661 5661 22695 5695
rect 22695 5661 22704 5695
rect 22652 5652 22704 5661
rect 23480 5652 23532 5704
rect 23848 5652 23900 5704
rect 25412 5695 25464 5704
rect 25412 5661 25421 5695
rect 25421 5661 25455 5695
rect 25455 5661 25464 5695
rect 25412 5652 25464 5661
rect 27436 5652 27488 5704
rect 27988 5720 28040 5772
rect 28172 5763 28224 5772
rect 28172 5729 28181 5763
rect 28181 5729 28215 5763
rect 28215 5729 28224 5763
rect 28172 5720 28224 5729
rect 29000 5695 29052 5704
rect 29000 5661 29009 5695
rect 29009 5661 29043 5695
rect 29043 5661 29052 5695
rect 29000 5652 29052 5661
rect 30196 5695 30248 5704
rect 30196 5661 30205 5695
rect 30205 5661 30239 5695
rect 30239 5661 30248 5695
rect 30196 5652 30248 5661
rect 38108 5652 38160 5704
rect 18144 5627 18196 5636
rect 18144 5593 18153 5627
rect 18153 5593 18187 5627
rect 18187 5593 18196 5627
rect 20904 5627 20956 5636
rect 18144 5584 18196 5593
rect 20904 5593 20913 5627
rect 20913 5593 20947 5627
rect 20947 5593 20956 5627
rect 20904 5584 20956 5593
rect 21364 5584 21416 5636
rect 21548 5627 21600 5636
rect 21548 5593 21557 5627
rect 21557 5593 21591 5627
rect 21591 5593 21600 5627
rect 21548 5584 21600 5593
rect 20168 5516 20220 5568
rect 20628 5516 20680 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 1492 5176 1544 5228
rect 7012 5312 7064 5364
rect 3976 5244 4028 5296
rect 11152 5244 11204 5296
rect 9220 5219 9272 5228
rect 9220 5185 9229 5219
rect 9229 5185 9263 5219
rect 9263 5185 9272 5219
rect 9220 5176 9272 5185
rect 5448 5083 5500 5092
rect 5448 5049 5457 5083
rect 5457 5049 5491 5083
rect 5491 5049 5500 5083
rect 5448 5040 5500 5049
rect 1768 5015 1820 5024
rect 1768 4981 1777 5015
rect 1777 4981 1811 5015
rect 1811 4981 1820 5015
rect 1768 4972 1820 4981
rect 2504 4972 2556 5024
rect 6276 5040 6328 5092
rect 10784 5108 10836 5160
rect 14004 5312 14056 5364
rect 14188 5244 14240 5296
rect 18512 5244 18564 5296
rect 20628 5244 20680 5296
rect 17132 5219 17184 5228
rect 17132 5185 17141 5219
rect 17141 5185 17175 5219
rect 17175 5185 17184 5219
rect 17132 5176 17184 5185
rect 17040 5108 17092 5160
rect 17224 5108 17276 5160
rect 17960 5151 18012 5160
rect 17960 5117 17969 5151
rect 17969 5117 18003 5151
rect 18003 5117 18012 5151
rect 17960 5108 18012 5117
rect 18328 5108 18380 5160
rect 18604 5108 18656 5160
rect 20628 5108 20680 5160
rect 21272 5312 21324 5364
rect 22928 5312 22980 5364
rect 23480 5312 23532 5364
rect 24584 5312 24636 5364
rect 25412 5312 25464 5364
rect 29000 5312 29052 5364
rect 29092 5312 29144 5364
rect 22376 5244 22428 5296
rect 22652 5244 22704 5296
rect 22468 5176 22520 5228
rect 24032 5176 24084 5228
rect 24584 5219 24636 5228
rect 24584 5185 24593 5219
rect 24593 5185 24627 5219
rect 24627 5185 24636 5219
rect 24584 5176 24636 5185
rect 24676 5176 24728 5228
rect 25872 5176 25924 5228
rect 26516 5244 26568 5296
rect 27988 5219 28040 5228
rect 19340 5040 19392 5092
rect 23388 5108 23440 5160
rect 26516 5040 26568 5092
rect 10692 4972 10744 5024
rect 11060 4972 11112 5024
rect 13912 4972 13964 5024
rect 15752 5015 15804 5024
rect 15752 4981 15761 5015
rect 15761 4981 15795 5015
rect 15795 4981 15804 5015
rect 15752 4972 15804 4981
rect 19432 4972 19484 5024
rect 19524 4972 19576 5024
rect 20076 4972 20128 5024
rect 21732 4972 21784 5024
rect 23940 4972 23992 5024
rect 24676 5015 24728 5024
rect 24676 4981 24685 5015
rect 24685 4981 24719 5015
rect 24719 4981 24728 5015
rect 24676 4972 24728 4981
rect 24768 4972 24820 5024
rect 27988 5185 27997 5219
rect 27997 5185 28031 5219
rect 28031 5185 28040 5219
rect 27988 5176 28040 5185
rect 36728 5244 36780 5296
rect 31208 5219 31260 5228
rect 31208 5185 31217 5219
rect 31217 5185 31251 5219
rect 31251 5185 31260 5219
rect 31208 5176 31260 5185
rect 33324 5040 33376 5092
rect 28080 4972 28132 5024
rect 32956 4972 33008 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 5724 4632 5776 4684
rect 11336 4768 11388 4820
rect 11980 4768 12032 4820
rect 12256 4811 12308 4820
rect 12256 4777 12265 4811
rect 12265 4777 12299 4811
rect 12299 4777 12308 4811
rect 12256 4768 12308 4777
rect 12348 4768 12400 4820
rect 14004 4768 14056 4820
rect 17040 4768 17092 4820
rect 24676 4768 24728 4820
rect 27988 4768 28040 4820
rect 16028 4743 16080 4752
rect 9680 4632 9732 4684
rect 16028 4709 16037 4743
rect 16037 4709 16071 4743
rect 16071 4709 16080 4743
rect 16028 4700 16080 4709
rect 16856 4700 16908 4752
rect 18144 4700 18196 4752
rect 18236 4743 18288 4752
rect 18236 4709 18245 4743
rect 18245 4709 18279 4743
rect 18279 4709 18288 4743
rect 18236 4700 18288 4709
rect 18420 4700 18472 4752
rect 19984 4700 20036 4752
rect 20628 4700 20680 4752
rect 24032 4743 24084 4752
rect 24032 4709 24041 4743
rect 24041 4709 24075 4743
rect 24075 4709 24084 4743
rect 24032 4700 24084 4709
rect 27712 4700 27764 4752
rect 3976 4607 4028 4616
rect 3976 4573 3985 4607
rect 3985 4573 4019 4607
rect 4019 4573 4028 4607
rect 3976 4564 4028 4573
rect 10508 4607 10560 4616
rect 10508 4573 10517 4607
rect 10517 4573 10551 4607
rect 10551 4573 10560 4607
rect 10508 4564 10560 4573
rect 19340 4632 19392 4684
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 17040 4564 17092 4616
rect 18052 4564 18104 4616
rect 19248 4564 19300 4616
rect 20076 4564 20128 4616
rect 22468 4632 22520 4684
rect 23388 4675 23440 4684
rect 23388 4641 23397 4675
rect 23397 4641 23431 4675
rect 23431 4641 23440 4675
rect 23388 4632 23440 4641
rect 24676 4632 24728 4684
rect 28080 4675 28132 4684
rect 22376 4564 22428 4616
rect 5908 4496 5960 4548
rect 11060 4496 11112 4548
rect 7288 4428 7340 4480
rect 12348 4496 12400 4548
rect 14464 4496 14516 4548
rect 24768 4564 24820 4616
rect 25228 4607 25280 4616
rect 25228 4573 25237 4607
rect 25237 4573 25271 4607
rect 25271 4573 25280 4607
rect 28080 4641 28089 4675
rect 28089 4641 28123 4675
rect 28123 4641 28132 4675
rect 28080 4632 28132 4641
rect 26516 4607 26568 4616
rect 25228 4564 25280 4573
rect 26516 4573 26525 4607
rect 26525 4573 26559 4607
rect 26559 4573 26568 4607
rect 26516 4564 26568 4573
rect 27896 4607 27948 4616
rect 12256 4428 12308 4480
rect 17224 4428 17276 4480
rect 17592 4471 17644 4480
rect 17592 4437 17601 4471
rect 17601 4437 17635 4471
rect 17635 4437 17644 4471
rect 17592 4428 17644 4437
rect 17684 4428 17736 4480
rect 25320 4496 25372 4548
rect 27896 4573 27905 4607
rect 27905 4573 27939 4607
rect 27939 4573 27948 4607
rect 27896 4564 27948 4573
rect 32864 4564 32916 4616
rect 34428 4564 34480 4616
rect 29736 4496 29788 4548
rect 25780 4428 25832 4480
rect 25872 4428 25924 4480
rect 38200 4471 38252 4480
rect 38200 4437 38209 4471
rect 38209 4437 38243 4471
rect 38243 4437 38252 4471
rect 38200 4428 38252 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 5908 4224 5960 4276
rect 13912 4224 13964 4276
rect 14004 4224 14056 4276
rect 16856 4224 16908 4276
rect 17132 4224 17184 4276
rect 17224 4224 17276 4276
rect 17592 4156 17644 4208
rect 2780 4088 2832 4140
rect 5816 4088 5868 4140
rect 7288 4088 7340 4140
rect 7380 4088 7432 4140
rect 8392 4131 8444 4140
rect 8392 4097 8401 4131
rect 8401 4097 8435 4131
rect 8435 4097 8444 4131
rect 8392 4088 8444 4097
rect 17684 4088 17736 4140
rect 17960 4156 18012 4208
rect 18328 4156 18380 4208
rect 18512 4156 18564 4208
rect 19984 4224 20036 4276
rect 24768 4224 24820 4276
rect 25780 4267 25832 4276
rect 25780 4233 25789 4267
rect 25789 4233 25823 4267
rect 25823 4233 25832 4267
rect 25780 4224 25832 4233
rect 27896 4224 27948 4276
rect 20076 4131 20128 4140
rect 20076 4097 20085 4131
rect 20085 4097 20119 4131
rect 20119 4097 20128 4131
rect 20076 4088 20128 4097
rect 20168 4131 20220 4140
rect 20168 4097 20177 4131
rect 20177 4097 20211 4131
rect 20211 4097 20220 4131
rect 21272 4131 21324 4140
rect 20168 4088 20220 4097
rect 21272 4097 21281 4131
rect 21281 4097 21315 4131
rect 21315 4097 21324 4131
rect 21272 4088 21324 4097
rect 21916 4088 21968 4140
rect 22652 4131 22704 4140
rect 22652 4097 22661 4131
rect 22661 4097 22695 4131
rect 22695 4097 22704 4131
rect 22652 4088 22704 4097
rect 23204 4088 23256 4140
rect 23480 4088 23532 4140
rect 24492 4131 24544 4140
rect 24492 4097 24501 4131
rect 24501 4097 24535 4131
rect 24535 4097 24544 4131
rect 24492 4088 24544 4097
rect 24676 4088 24728 4140
rect 10508 4020 10560 4072
rect 11612 4020 11664 4072
rect 12992 4063 13044 4072
rect 1676 3952 1728 4004
rect 12992 4029 13001 4063
rect 13001 4029 13035 4063
rect 13035 4029 13044 4063
rect 12992 4020 13044 4029
rect 13452 4020 13504 4072
rect 19064 4020 19116 4072
rect 14280 3884 14332 3936
rect 14648 3884 14700 3936
rect 14740 3884 14792 3936
rect 17776 3884 17828 3936
rect 24400 4020 24452 4072
rect 26148 4088 26200 4140
rect 23480 3952 23532 4004
rect 25412 3952 25464 4004
rect 20720 3884 20772 3936
rect 22192 3884 22244 3936
rect 22836 3884 22888 3936
rect 23848 3884 23900 3936
rect 28172 4131 28224 4140
rect 28172 4097 28181 4131
rect 28181 4097 28215 4131
rect 28215 4097 28224 4131
rect 28172 4088 28224 4097
rect 29276 4088 29328 4140
rect 30196 4088 30248 4140
rect 30748 4063 30800 4072
rect 30748 4029 30757 4063
rect 30757 4029 30791 4063
rect 30791 4029 30800 4063
rect 30748 4020 30800 4029
rect 31668 3952 31720 4004
rect 27068 3884 27120 3936
rect 28724 3884 28776 3936
rect 29368 3927 29420 3936
rect 29368 3893 29377 3927
rect 29377 3893 29411 3927
rect 29411 3893 29420 3927
rect 29368 3884 29420 3893
rect 30656 3884 30708 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 1860 3680 1912 3732
rect 7472 3680 7524 3732
rect 9036 3680 9088 3732
rect 10140 3680 10192 3732
rect 11060 3680 11112 3732
rect 15384 3680 15436 3732
rect 18512 3680 18564 3732
rect 18604 3680 18656 3732
rect 24492 3680 24544 3732
rect 11428 3612 11480 3664
rect 12992 3612 13044 3664
rect 14740 3612 14792 3664
rect 17316 3612 17368 3664
rect 25596 3680 25648 3732
rect 25688 3680 25740 3732
rect 26608 3680 26660 3732
rect 30840 3723 30892 3732
rect 30840 3689 30849 3723
rect 30849 3689 30883 3723
rect 30883 3689 30892 3723
rect 30840 3680 30892 3689
rect 33048 3680 33100 3732
rect 28172 3612 28224 3664
rect 37280 3612 37332 3664
rect 4068 3544 4120 3596
rect 7196 3544 7248 3596
rect 1768 3519 1820 3528
rect 1768 3485 1777 3519
rect 1777 3485 1811 3519
rect 1811 3485 1820 3519
rect 1768 3476 1820 3485
rect 14188 3544 14240 3596
rect 15292 3544 15344 3596
rect 15384 3544 15436 3596
rect 20352 3544 20404 3596
rect 7840 3408 7892 3460
rect 14372 3476 14424 3528
rect 15016 3519 15068 3528
rect 15016 3485 15025 3519
rect 15025 3485 15059 3519
rect 15059 3485 15068 3519
rect 15016 3476 15068 3485
rect 17040 3476 17092 3528
rect 18052 3476 18104 3528
rect 18696 3515 18748 3528
rect 18696 3481 18705 3515
rect 18705 3481 18739 3515
rect 18739 3481 18748 3515
rect 18696 3476 18748 3481
rect 18880 3476 18932 3528
rect 20444 3476 20496 3528
rect 29368 3544 29420 3596
rect 30656 3587 30708 3596
rect 30656 3553 30665 3587
rect 30665 3553 30699 3587
rect 30699 3553 30708 3587
rect 30656 3544 30708 3553
rect 21088 3476 21140 3528
rect 22468 3476 22520 3528
rect 23204 3476 23256 3528
rect 24584 3519 24636 3528
rect 24584 3485 24593 3519
rect 24593 3485 24627 3519
rect 24627 3485 24636 3519
rect 24584 3476 24636 3485
rect 25780 3476 25832 3528
rect 26424 3476 26476 3528
rect 27804 3476 27856 3528
rect 28080 3519 28132 3528
rect 28080 3485 28089 3519
rect 28089 3485 28123 3519
rect 28123 3485 28132 3519
rect 28080 3476 28132 3485
rect 9036 3408 9088 3460
rect 14464 3408 14516 3460
rect 18972 3408 19024 3460
rect 23388 3451 23440 3460
rect 23388 3417 23397 3451
rect 23397 3417 23431 3451
rect 23431 3417 23440 3451
rect 23388 3408 23440 3417
rect 23480 3451 23532 3460
rect 23480 3417 23489 3451
rect 23489 3417 23523 3451
rect 23523 3417 23532 3451
rect 24032 3451 24084 3460
rect 23480 3408 23532 3417
rect 24032 3417 24041 3451
rect 24041 3417 24075 3451
rect 24075 3417 24084 3451
rect 24032 3408 24084 3417
rect 24400 3408 24452 3460
rect 11520 3340 11572 3392
rect 14372 3340 14424 3392
rect 15752 3340 15804 3392
rect 17224 3383 17276 3392
rect 17224 3349 17233 3383
rect 17233 3349 17267 3383
rect 17267 3349 17276 3383
rect 17224 3340 17276 3349
rect 18144 3340 18196 3392
rect 19984 3383 20036 3392
rect 19984 3349 19993 3383
rect 19993 3349 20027 3383
rect 20027 3349 20036 3383
rect 19984 3340 20036 3349
rect 20168 3340 20220 3392
rect 21364 3340 21416 3392
rect 23848 3340 23900 3392
rect 24124 3340 24176 3392
rect 25596 3408 25648 3460
rect 31024 3476 31076 3528
rect 33692 3476 33744 3528
rect 38292 3519 38344 3528
rect 38292 3485 38301 3519
rect 38301 3485 38335 3519
rect 38335 3485 38344 3519
rect 38292 3476 38344 3485
rect 27068 3340 27120 3392
rect 27344 3383 27396 3392
rect 27344 3349 27353 3383
rect 27353 3349 27387 3383
rect 27387 3349 27396 3383
rect 27344 3340 27396 3349
rect 27896 3383 27948 3392
rect 27896 3349 27905 3383
rect 27905 3349 27939 3383
rect 27939 3349 27948 3383
rect 27896 3340 27948 3349
rect 28540 3383 28592 3392
rect 28540 3349 28549 3383
rect 28549 3349 28583 3383
rect 28583 3349 28592 3383
rect 28540 3340 28592 3349
rect 28816 3340 28868 3392
rect 31208 3340 31260 3392
rect 31576 3383 31628 3392
rect 31576 3349 31585 3383
rect 31585 3349 31619 3383
rect 31619 3349 31628 3383
rect 31576 3340 31628 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 5816 3136 5868 3188
rect 13452 3179 13504 3188
rect 13452 3145 13461 3179
rect 13461 3145 13495 3179
rect 13495 3145 13504 3179
rect 13452 3136 13504 3145
rect 6644 3068 6696 3120
rect 7472 3068 7524 3120
rect 9680 3068 9732 3120
rect 11520 3068 11572 3120
rect 12072 3068 12124 3120
rect 17224 3136 17276 3188
rect 2504 3043 2556 3052
rect 2504 3009 2513 3043
rect 2513 3009 2547 3043
rect 2547 3009 2556 3043
rect 2504 3000 2556 3009
rect 3332 3043 3384 3052
rect 3332 3009 3341 3043
rect 3341 3009 3375 3043
rect 3375 3009 3384 3043
rect 3332 3000 3384 3009
rect 4068 3000 4120 3052
rect 9128 3043 9180 3052
rect 5448 2932 5500 2984
rect 9128 3009 9137 3043
rect 9137 3009 9171 3043
rect 9171 3009 9180 3043
rect 9128 3000 9180 3009
rect 14280 3068 14332 3120
rect 14372 3111 14424 3120
rect 14372 3077 14381 3111
rect 14381 3077 14415 3111
rect 14415 3077 14424 3111
rect 14372 3068 14424 3077
rect 17868 3068 17920 3120
rect 7196 2932 7248 2984
rect 10048 2932 10100 2984
rect 20 2796 72 2848
rect 5816 2796 5868 2848
rect 10140 2796 10192 2848
rect 21272 3136 21324 3188
rect 23388 3136 23440 3188
rect 20812 3068 20864 3120
rect 22192 3111 22244 3120
rect 22192 3077 22201 3111
rect 22201 3077 22235 3111
rect 22235 3077 22244 3111
rect 22192 3068 22244 3077
rect 23572 3068 23624 3120
rect 14464 2932 14516 2984
rect 18052 3000 18104 3052
rect 16120 2975 16172 2984
rect 16120 2941 16129 2975
rect 16129 2941 16163 2975
rect 16163 2941 16172 2975
rect 18328 3000 18380 3052
rect 21916 3000 21968 3052
rect 24124 3043 24176 3052
rect 16120 2932 16172 2941
rect 18788 2932 18840 2984
rect 19156 2975 19208 2984
rect 19156 2941 19165 2975
rect 19165 2941 19199 2975
rect 19199 2941 19208 2975
rect 19156 2932 19208 2941
rect 22100 2975 22152 2984
rect 22100 2941 22109 2975
rect 22109 2941 22143 2975
rect 22143 2941 22152 2975
rect 24124 3009 24133 3043
rect 24133 3009 24167 3043
rect 24167 3009 24176 3043
rect 24124 3000 24176 3009
rect 31024 3179 31076 3188
rect 31024 3145 31033 3179
rect 31033 3145 31067 3179
rect 31067 3145 31076 3179
rect 31024 3136 31076 3145
rect 36728 3179 36780 3188
rect 36728 3145 36737 3179
rect 36737 3145 36771 3179
rect 36771 3145 36780 3179
rect 36728 3136 36780 3145
rect 26148 3068 26200 3120
rect 28540 3068 28592 3120
rect 28816 3111 28868 3120
rect 28816 3077 28825 3111
rect 28825 3077 28859 3111
rect 28859 3077 28868 3111
rect 28816 3068 28868 3077
rect 31576 3068 31628 3120
rect 32956 3068 33008 3120
rect 22100 2932 22152 2941
rect 15752 2864 15804 2916
rect 18604 2864 18656 2916
rect 20720 2864 20772 2916
rect 20168 2796 20220 2848
rect 20536 2796 20588 2848
rect 24032 2932 24084 2984
rect 27896 3000 27948 3052
rect 27988 3000 28040 3052
rect 31208 3043 31260 3052
rect 31208 3009 31217 3043
rect 31217 3009 31251 3043
rect 31251 3009 31260 3043
rect 31208 3000 31260 3009
rect 32496 3043 32548 3052
rect 32496 3009 32505 3043
rect 32505 3009 32539 3043
rect 32539 3009 32548 3043
rect 32496 3000 32548 3009
rect 25688 2864 25740 2916
rect 27068 2796 27120 2848
rect 27252 2864 27304 2916
rect 30748 2932 30800 2984
rect 39304 2932 39356 2984
rect 27804 2796 27856 2848
rect 29920 2796 29972 2848
rect 30288 2796 30340 2848
rect 31760 2796 31812 2848
rect 32312 2839 32364 2848
rect 32312 2805 32321 2839
rect 32321 2805 32355 2839
rect 32355 2805 32364 2839
rect 32312 2796 32364 2805
rect 38200 2839 38252 2848
rect 38200 2805 38209 2839
rect 38209 2805 38243 2839
rect 38243 2805 38252 2839
rect 38200 2796 38252 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 2412 2592 2464 2644
rect 7380 2592 7432 2644
rect 7472 2592 7524 2644
rect 10324 2592 10376 2644
rect 15016 2592 15068 2644
rect 7012 2524 7064 2576
rect 17960 2592 18012 2644
rect 18052 2592 18104 2644
rect 22100 2592 22152 2644
rect 23756 2592 23808 2644
rect 25504 2592 25556 2644
rect 2872 2456 2924 2508
rect 3976 2499 4028 2508
rect 3976 2465 3985 2499
rect 3985 2465 4019 2499
rect 4019 2465 4028 2499
rect 3976 2456 4028 2465
rect 7196 2456 7248 2508
rect 2596 2388 2648 2440
rect 1308 2252 1360 2304
rect 5816 2388 5868 2440
rect 6644 2388 6696 2440
rect 16672 2524 16724 2576
rect 20720 2524 20772 2576
rect 19984 2456 20036 2508
rect 7748 2431 7800 2440
rect 7748 2397 7757 2431
rect 7757 2397 7791 2431
rect 7791 2397 7800 2431
rect 7748 2388 7800 2397
rect 10784 2388 10836 2440
rect 11612 2388 11664 2440
rect 13544 2388 13596 2440
rect 14832 2388 14884 2440
rect 16764 2388 16816 2440
rect 18144 2431 18196 2440
rect 18144 2397 18153 2431
rect 18153 2397 18187 2431
rect 18187 2397 18196 2431
rect 18144 2388 18196 2397
rect 19340 2388 19392 2440
rect 20168 2431 20220 2440
rect 20168 2397 20177 2431
rect 20177 2397 20211 2431
rect 20211 2397 20220 2431
rect 20168 2388 20220 2397
rect 21272 2388 21324 2440
rect 4528 2252 4580 2304
rect 5816 2252 5868 2304
rect 9036 2252 9088 2304
rect 10324 2252 10376 2304
rect 11704 2295 11756 2304
rect 11704 2261 11713 2295
rect 11713 2261 11747 2295
rect 11747 2261 11756 2295
rect 11704 2252 11756 2261
rect 16672 2252 16724 2304
rect 22560 2320 22612 2372
rect 25412 2388 25464 2440
rect 28080 2592 28132 2644
rect 29736 2635 29788 2644
rect 29736 2601 29745 2635
rect 29745 2601 29779 2635
rect 29779 2601 29788 2635
rect 29736 2592 29788 2601
rect 32496 2592 32548 2644
rect 32864 2592 32916 2644
rect 33692 2635 33744 2644
rect 28724 2431 28776 2440
rect 27068 2320 27120 2372
rect 28724 2397 28733 2431
rect 28733 2397 28767 2431
rect 28767 2397 28776 2431
rect 28724 2388 28776 2397
rect 29920 2431 29972 2440
rect 29920 2397 29929 2431
rect 29929 2397 29963 2431
rect 29963 2397 29972 2431
rect 29920 2388 29972 2397
rect 30380 2431 30432 2440
rect 30380 2397 30389 2431
rect 30389 2397 30423 2431
rect 30423 2397 30432 2431
rect 30380 2388 30432 2397
rect 29000 2320 29052 2372
rect 31668 2524 31720 2576
rect 33692 2601 33701 2635
rect 33701 2601 33735 2635
rect 33735 2601 33744 2635
rect 33692 2592 33744 2601
rect 31760 2456 31812 2508
rect 32312 2431 32364 2440
rect 32312 2397 32321 2431
rect 32321 2397 32355 2431
rect 32355 2397 32364 2431
rect 32312 2388 32364 2397
rect 33324 2456 33376 2508
rect 33508 2388 33560 2440
rect 34796 2388 34848 2440
rect 36084 2388 36136 2440
rect 18052 2252 18104 2304
rect 19340 2252 19392 2304
rect 21180 2252 21232 2304
rect 23848 2252 23900 2304
rect 26148 2252 26200 2304
rect 27436 2252 27488 2304
rect 31576 2252 31628 2304
rect 38016 2252 38068 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 7012 2048 7064 2100
rect 11980 2048 12032 2100
rect 17960 2048 18012 2100
rect 22836 2048 22888 2100
rect 11704 1980 11756 2032
rect 26424 1980 26476 2032
rect 7748 1912 7800 1964
rect 23940 1912 23992 1964
rect 19248 1844 19300 1896
rect 21180 1844 21232 1896
<< metal2 >>
rect 18 39200 74 39800
rect 1306 39200 1362 39800
rect 3238 39200 3294 39800
rect 4526 39200 4582 39800
rect 5814 39200 5870 39800
rect 7746 39200 7802 39800
rect 9034 39200 9090 39800
rect 10322 39200 10378 39800
rect 12254 39200 12310 39800
rect 13542 39200 13598 39800
rect 15474 39200 15530 39800
rect 16762 39200 16818 39800
rect 18050 39200 18106 39800
rect 19982 39200 20038 39800
rect 21270 39200 21326 39800
rect 22558 39200 22614 39800
rect 24490 39200 24546 39800
rect 25778 39200 25834 39800
rect 27710 39200 27766 39800
rect 28998 39200 29054 39800
rect 30286 39200 30342 39800
rect 32218 39200 32274 39800
rect 33506 39200 33562 39800
rect 34794 39200 34850 39800
rect 36726 39200 36782 39800
rect 38014 39200 38070 39800
rect 39302 39200 39358 39800
rect 32 36922 60 39200
rect 1320 37126 1348 39200
rect 3146 38176 3202 38185
rect 3146 38111 3202 38120
rect 3160 37262 3188 38111
rect 3252 37262 3280 39200
rect 4540 37754 4568 39200
rect 4540 37726 4660 37754
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4632 37262 4660 37726
rect 2780 37256 2832 37262
rect 2780 37198 2832 37204
rect 3148 37256 3200 37262
rect 3148 37198 3200 37204
rect 3240 37256 3292 37262
rect 3240 37198 3292 37204
rect 4620 37256 4672 37262
rect 4620 37198 4672 37204
rect 1308 37120 1360 37126
rect 1308 37062 1360 37068
rect 2320 37120 2372 37126
rect 2320 37062 2372 37068
rect 20 36916 72 36922
rect 20 36858 72 36864
rect 2332 36854 2360 37062
rect 2320 36848 2372 36854
rect 2792 36825 2820 37198
rect 4068 37188 4120 37194
rect 4068 37130 4120 37136
rect 2964 37120 3016 37126
rect 2964 37062 3016 37068
rect 3976 37120 4028 37126
rect 3976 37062 4028 37068
rect 2320 36790 2372 36796
rect 2778 36816 2834 36825
rect 2778 36751 2834 36760
rect 1768 33516 1820 33522
rect 1768 33458 1820 33464
rect 1780 33425 1808 33458
rect 1766 33416 1822 33425
rect 1766 33351 1822 33360
rect 1768 32428 1820 32434
rect 1768 32370 1820 32376
rect 1780 32065 1808 32370
rect 1766 32056 1822 32065
rect 1766 31991 1822 32000
rect 1584 30728 1636 30734
rect 1582 30696 1584 30705
rect 1860 30728 1912 30734
rect 1636 30696 1638 30705
rect 1860 30670 1912 30676
rect 1582 30631 1638 30640
rect 1768 29164 1820 29170
rect 1768 29106 1820 29112
rect 1780 28665 1808 29106
rect 1766 28656 1822 28665
rect 1766 28591 1822 28600
rect 1768 27464 1820 27470
rect 1768 27406 1820 27412
rect 1780 27305 1808 27406
rect 1766 27296 1822 27305
rect 1766 27231 1822 27240
rect 1768 25288 1820 25294
rect 1766 25256 1768 25265
rect 1820 25256 1822 25265
rect 1766 25191 1822 25200
rect 1584 24200 1636 24206
rect 1584 24142 1636 24148
rect 1596 23866 1624 24142
rect 1768 24064 1820 24070
rect 1768 24006 1820 24012
rect 1780 23905 1808 24006
rect 1766 23896 1822 23905
rect 1584 23860 1636 23866
rect 1766 23831 1822 23840
rect 1584 23802 1636 23808
rect 1768 22636 1820 22642
rect 1768 22578 1820 22584
rect 1780 22545 1808 22578
rect 1766 22536 1822 22545
rect 1766 22471 1822 22480
rect 1768 20936 1820 20942
rect 1768 20878 1820 20884
rect 1780 20505 1808 20878
rect 1766 20496 1822 20505
rect 1766 20431 1822 20440
rect 1768 19168 1820 19174
rect 1766 19136 1768 19145
rect 1820 19136 1822 19145
rect 1766 19071 1822 19080
rect 1768 18284 1820 18290
rect 1768 18226 1820 18232
rect 1780 17785 1808 18226
rect 1766 17776 1822 17785
rect 1766 17711 1822 17720
rect 1584 16108 1636 16114
rect 1584 16050 1636 16056
rect 1492 14272 1544 14278
rect 1492 14214 1544 14220
rect 1504 5234 1532 14214
rect 1596 14074 1624 16050
rect 1768 15904 1820 15910
rect 1768 15846 1820 15852
rect 1780 15745 1808 15846
rect 1766 15736 1822 15745
rect 1766 15671 1822 15680
rect 1768 15020 1820 15026
rect 1768 14962 1820 14968
rect 1780 14385 1808 14962
rect 1766 14376 1822 14385
rect 1766 14311 1822 14320
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 1584 13320 1636 13326
rect 1584 13262 1636 13268
rect 1596 12986 1624 13262
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 1768 12844 1820 12850
rect 1768 12786 1820 12792
rect 1780 12345 1808 12786
rect 1872 12714 1900 30670
rect 2976 29646 3004 37062
rect 2964 29640 3016 29646
rect 2964 29582 3016 29588
rect 3988 28082 4016 37062
rect 4080 35290 4108 37130
rect 5828 37126 5856 39200
rect 7760 37126 7788 39200
rect 9048 37262 9076 39200
rect 7840 37256 7892 37262
rect 7840 37198 7892 37204
rect 9036 37256 9088 37262
rect 9036 37198 9088 37204
rect 4620 37120 4672 37126
rect 4620 37062 4672 37068
rect 5816 37120 5868 37126
rect 5816 37062 5868 37068
rect 7748 37120 7800 37126
rect 7748 37062 7800 37068
rect 4632 36922 4660 37062
rect 4620 36916 4672 36922
rect 4620 36858 4672 36864
rect 7656 36848 7708 36854
rect 7656 36790 7708 36796
rect 4620 36780 4672 36786
rect 4620 36722 4672 36728
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4068 35284 4120 35290
rect 4068 35226 4120 35232
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4632 32570 4660 36722
rect 7196 33312 7248 33318
rect 7196 33254 7248 33260
rect 4620 32564 4672 32570
rect 4620 32506 4672 32512
rect 4620 32428 4672 32434
rect 4620 32370 4672 32376
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 3976 28076 4028 28082
rect 3976 28018 4028 28024
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 3148 25152 3200 25158
rect 3148 25094 3200 25100
rect 3160 22642 3188 25094
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4632 24410 4660 32370
rect 6276 32224 6328 32230
rect 6276 32166 6328 32172
rect 5172 30184 5224 30190
rect 5172 30126 5224 30132
rect 5184 29850 5212 30126
rect 5172 29844 5224 29850
rect 5172 29786 5224 29792
rect 5724 29028 5776 29034
rect 5724 28970 5776 28976
rect 5736 27470 5764 28970
rect 5908 27668 5960 27674
rect 5908 27610 5960 27616
rect 5724 27464 5776 27470
rect 5724 27406 5776 27412
rect 5356 27328 5408 27334
rect 5356 27270 5408 27276
rect 5816 27328 5868 27334
rect 5816 27270 5868 27276
rect 5368 24818 5396 27270
rect 5828 26994 5856 27270
rect 5816 26988 5868 26994
rect 5816 26930 5868 26936
rect 5356 24812 5408 24818
rect 5356 24754 5408 24760
rect 5356 24608 5408 24614
rect 5356 24550 5408 24556
rect 4620 24404 4672 24410
rect 4620 24346 4672 24352
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 5368 22710 5396 24550
rect 5356 22704 5408 22710
rect 5356 22646 5408 22652
rect 5724 22704 5776 22710
rect 5724 22646 5776 22652
rect 3148 22636 3200 22642
rect 3148 22578 3200 22584
rect 3240 22432 3292 22438
rect 3240 22374 3292 22380
rect 3252 20466 3280 22374
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 5264 22160 5316 22166
rect 5264 22102 5316 22108
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 3792 20936 3844 20942
rect 3792 20878 3844 20884
rect 3240 20460 3292 20466
rect 3240 20402 3292 20408
rect 3424 19372 3476 19378
rect 3424 19314 3476 19320
rect 2320 17672 2372 17678
rect 2320 17614 2372 17620
rect 2044 17128 2096 17134
rect 2044 17070 2096 17076
rect 1952 13932 2004 13938
rect 1952 13874 2004 13880
rect 1860 12708 1912 12714
rect 1860 12650 1912 12656
rect 1964 12442 1992 13874
rect 1952 12436 2004 12442
rect 1952 12378 2004 12384
rect 1766 12336 1822 12345
rect 1766 12271 1822 12280
rect 1952 11280 2004 11286
rect 1952 11222 2004 11228
rect 1768 11144 1820 11150
rect 1768 11086 1820 11092
rect 1780 10985 1808 11086
rect 1766 10976 1822 10985
rect 1766 10911 1822 10920
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 1596 5914 1624 10610
rect 1768 10056 1820 10062
rect 1768 9998 1820 10004
rect 1780 9625 1808 9998
rect 1860 9920 1912 9926
rect 1860 9862 1912 9868
rect 1766 9616 1822 9625
rect 1766 9551 1822 9560
rect 1872 8974 1900 9862
rect 1860 8968 1912 8974
rect 1860 8910 1912 8916
rect 1860 7880 1912 7886
rect 1860 7822 1912 7828
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1584 5908 1636 5914
rect 1584 5850 1636 5856
rect 1492 5228 1544 5234
rect 1492 5170 1544 5176
rect 1688 4010 1716 7346
rect 1766 6216 1822 6225
rect 1766 6151 1822 6160
rect 1780 5710 1808 6151
rect 1768 5704 1820 5710
rect 1768 5646 1820 5652
rect 1768 5024 1820 5030
rect 1768 4966 1820 4972
rect 1780 4865 1808 4966
rect 1766 4856 1822 4865
rect 1766 4791 1822 4800
rect 1676 4004 1728 4010
rect 1676 3946 1728 3952
rect 1872 3738 1900 7822
rect 1964 6322 1992 11222
rect 2056 8634 2084 17070
rect 2332 16794 2360 17614
rect 3240 17332 3292 17338
rect 3240 17274 3292 17280
rect 2320 16788 2372 16794
rect 2320 16730 2372 16736
rect 3252 16590 3280 17274
rect 3332 17128 3384 17134
rect 3332 17070 3384 17076
rect 3344 16590 3372 17070
rect 3240 16584 3292 16590
rect 3240 16526 3292 16532
rect 3332 16584 3384 16590
rect 3332 16526 3384 16532
rect 2872 15904 2924 15910
rect 2872 15846 2924 15852
rect 2884 14414 2912 15846
rect 2872 14408 2924 14414
rect 2872 14350 2924 14356
rect 3436 14074 3464 19314
rect 3804 18426 3832 20878
rect 4620 20392 4672 20398
rect 4620 20334 4672 20340
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4632 18970 4660 20334
rect 5080 20256 5132 20262
rect 5080 20198 5132 20204
rect 5172 20256 5224 20262
rect 5172 20198 5224 20204
rect 5092 19922 5120 20198
rect 5080 19916 5132 19922
rect 5080 19858 5132 19864
rect 5092 19514 5120 19858
rect 5184 19786 5212 20198
rect 5172 19780 5224 19786
rect 5172 19722 5224 19728
rect 5080 19508 5132 19514
rect 5080 19450 5132 19456
rect 4620 18964 4672 18970
rect 4620 18906 4672 18912
rect 4988 18896 5040 18902
rect 4988 18838 5040 18844
rect 4804 18692 4856 18698
rect 4804 18634 4856 18640
rect 3792 18420 3844 18426
rect 3792 18362 3844 18368
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4620 17536 4672 17542
rect 4620 17478 4672 17484
rect 4632 17270 4660 17478
rect 4620 17264 4672 17270
rect 4620 17206 4672 17212
rect 3884 17196 3936 17202
rect 3884 17138 3936 17144
rect 3896 16658 3924 17138
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 3884 16652 3936 16658
rect 3884 16594 3936 16600
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 3516 14952 3568 14958
rect 3516 14894 3568 14900
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 2412 13932 2464 13938
rect 2412 13874 2464 13880
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 2320 8492 2372 8498
rect 2320 8434 2372 8440
rect 2332 6914 2360 8434
rect 2424 8090 2452 13874
rect 3528 13870 3556 14894
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 3516 13864 3568 13870
rect 3516 13806 3568 13812
rect 3792 13864 3844 13870
rect 3792 13806 3844 13812
rect 3804 12986 3832 13806
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 3884 13388 3936 13394
rect 3884 13330 3936 13336
rect 3792 12980 3844 12986
rect 3792 12922 3844 12928
rect 3896 12646 3924 13330
rect 3988 13326 4016 13670
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 3976 13320 4028 13326
rect 3976 13262 4028 13268
rect 3884 12640 3936 12646
rect 3884 12582 3936 12588
rect 3988 12238 4016 13262
rect 4632 12782 4660 17206
rect 4712 17196 4764 17202
rect 4712 17138 4764 17144
rect 4724 16794 4752 17138
rect 4712 16788 4764 16794
rect 4712 16730 4764 16736
rect 4712 16448 4764 16454
rect 4712 16390 4764 16396
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4724 12434 4752 16390
rect 4816 16250 4844 18634
rect 4896 16584 4948 16590
rect 4896 16526 4948 16532
rect 4804 16244 4856 16250
rect 4804 16186 4856 16192
rect 4908 13530 4936 16526
rect 5000 15026 5028 18838
rect 5080 18760 5132 18766
rect 5080 18702 5132 18708
rect 4988 15020 5040 15026
rect 4988 14962 5040 14968
rect 5092 14822 5120 18702
rect 5172 18624 5224 18630
rect 5172 18566 5224 18572
rect 5080 14816 5132 14822
rect 5080 14758 5132 14764
rect 5184 14006 5212 18566
rect 5276 16402 5304 22102
rect 5356 20800 5408 20806
rect 5356 20742 5408 20748
rect 5368 18290 5396 20742
rect 5736 20602 5764 22646
rect 5816 22500 5868 22506
rect 5816 22442 5868 22448
rect 5828 22030 5856 22442
rect 5816 22024 5868 22030
rect 5816 21966 5868 21972
rect 5724 20596 5776 20602
rect 5724 20538 5776 20544
rect 5816 20460 5868 20466
rect 5816 20402 5868 20408
rect 5632 20392 5684 20398
rect 5632 20334 5684 20340
rect 5448 19372 5500 19378
rect 5448 19314 5500 19320
rect 5356 18284 5408 18290
rect 5356 18226 5408 18232
rect 5460 17882 5488 19314
rect 5644 18834 5672 20334
rect 5828 19174 5856 20402
rect 5816 19168 5868 19174
rect 5816 19110 5868 19116
rect 5632 18828 5684 18834
rect 5632 18770 5684 18776
rect 5448 17876 5500 17882
rect 5448 17818 5500 17824
rect 5644 17678 5672 18770
rect 5632 17672 5684 17678
rect 5632 17614 5684 17620
rect 5448 17536 5500 17542
rect 5448 17478 5500 17484
rect 5356 17196 5408 17202
rect 5356 17138 5408 17144
rect 5368 16794 5396 17138
rect 5356 16788 5408 16794
rect 5356 16730 5408 16736
rect 5276 16374 5396 16402
rect 5368 14958 5396 16374
rect 5356 14952 5408 14958
rect 5276 14900 5356 14906
rect 5276 14894 5408 14900
rect 5276 14878 5396 14894
rect 5172 14000 5224 14006
rect 5172 13942 5224 13948
rect 4896 13524 4948 13530
rect 4896 13466 4948 13472
rect 4724 12406 4936 12434
rect 3976 12232 4028 12238
rect 3976 12174 4028 12180
rect 3988 11694 4016 12174
rect 3976 11688 4028 11694
rect 3976 11630 4028 11636
rect 3988 11150 4016 11630
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 3988 10062 4016 11086
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 3988 8294 4016 9998
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 2412 8084 2464 8090
rect 2412 8026 2464 8032
rect 3988 7886 4016 8230
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 8072 4660 10202
rect 4908 9926 4936 12406
rect 5172 11688 5224 11694
rect 5172 11630 5224 11636
rect 4896 9920 4948 9926
rect 4896 9862 4948 9868
rect 4540 8044 4660 8072
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 2792 7585 2820 7822
rect 2778 7576 2834 7585
rect 2778 7511 2834 7520
rect 2332 6886 2452 6914
rect 1952 6316 2004 6322
rect 1952 6258 2004 6264
rect 1860 3732 1912 3738
rect 1860 3674 1912 3680
rect 1768 3528 1820 3534
rect 1768 3470 1820 3476
rect 20 2848 72 2854
rect 1780 2825 1808 3470
rect 20 2790 72 2796
rect 1766 2816 1822 2825
rect 32 800 60 2790
rect 1766 2751 1822 2760
rect 2424 2650 2452 6886
rect 2872 6656 2924 6662
rect 2872 6598 2924 6604
rect 2504 5024 2556 5030
rect 2504 4966 2556 4972
rect 2516 3058 2544 4966
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 2504 3052 2556 3058
rect 2504 2994 2556 3000
rect 2412 2644 2464 2650
rect 2412 2586 2464 2592
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 1308 2304 1360 2310
rect 1308 2246 1360 2252
rect 1320 800 1348 2246
rect 2608 800 2636 2382
rect 2792 1465 2820 4082
rect 2884 2514 2912 6598
rect 3988 6254 4016 7822
rect 4540 7818 4568 8044
rect 4528 7812 4580 7818
rect 4528 7754 4580 7760
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 3988 5710 4016 6190
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 3976 5704 4028 5710
rect 5184 5681 5212 11630
rect 5276 10130 5304 14878
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5264 10124 5316 10130
rect 5264 10066 5316 10072
rect 5368 6746 5396 14758
rect 5460 10742 5488 17478
rect 5632 16788 5684 16794
rect 5632 16730 5684 16736
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 5552 11234 5580 15302
rect 5644 14822 5672 16730
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 5632 14612 5684 14618
rect 5632 14554 5684 14560
rect 5644 12306 5672 14554
rect 5632 12300 5684 12306
rect 5632 12242 5684 12248
rect 5552 11206 5672 11234
rect 5644 11150 5672 11206
rect 5632 11144 5684 11150
rect 5632 11086 5684 11092
rect 5448 10736 5500 10742
rect 5448 10678 5500 10684
rect 5736 8090 5764 16050
rect 5828 12238 5856 19110
rect 5920 18834 5948 27610
rect 6184 25288 6236 25294
rect 6184 25230 6236 25236
rect 6000 22568 6052 22574
rect 6000 22510 6052 22516
rect 6012 21146 6040 22510
rect 6000 21140 6052 21146
rect 6000 21082 6052 21088
rect 6092 19984 6144 19990
rect 6092 19926 6144 19932
rect 6104 18834 6132 19926
rect 5908 18828 5960 18834
rect 5908 18770 5960 18776
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 5908 17672 5960 17678
rect 5908 17614 5960 17620
rect 5920 14618 5948 17614
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 5908 14612 5960 14618
rect 5908 14554 5960 14560
rect 5908 14000 5960 14006
rect 5908 13942 5960 13948
rect 5816 12232 5868 12238
rect 5816 12174 5868 12180
rect 5920 11354 5948 13942
rect 5908 11348 5960 11354
rect 5908 11290 5960 11296
rect 5908 9988 5960 9994
rect 6012 9976 6040 17138
rect 6104 10742 6132 18770
rect 6196 14006 6224 25230
rect 6288 24818 6316 32166
rect 6828 27872 6880 27878
rect 6828 27814 6880 27820
rect 6840 27674 6868 27814
rect 6828 27668 6880 27674
rect 6828 27610 6880 27616
rect 7208 27470 7236 33254
rect 7288 30184 7340 30190
rect 7288 30126 7340 30132
rect 7300 29850 7328 30126
rect 7288 29844 7340 29850
rect 7288 29786 7340 29792
rect 7668 28558 7696 36790
rect 7852 32026 7880 37198
rect 10336 37126 10364 39200
rect 11244 37256 11296 37262
rect 11244 37198 11296 37204
rect 11704 37256 11756 37262
rect 11704 37198 11756 37204
rect 8944 37120 8996 37126
rect 8944 37062 8996 37068
rect 10324 37120 10376 37126
rect 10324 37062 10376 37068
rect 7840 32020 7892 32026
rect 7840 31962 7892 31968
rect 8668 30048 8720 30054
rect 8668 29990 8720 29996
rect 8484 29640 8536 29646
rect 8484 29582 8536 29588
rect 8024 29096 8076 29102
rect 8024 29038 8076 29044
rect 8208 29096 8260 29102
rect 8208 29038 8260 29044
rect 8036 28694 8064 29038
rect 8024 28688 8076 28694
rect 8024 28630 8076 28636
rect 7656 28552 7708 28558
rect 7656 28494 7708 28500
rect 8220 28218 8248 29038
rect 8496 28558 8524 29582
rect 8680 29578 8708 29990
rect 8668 29572 8720 29578
rect 8668 29514 8720 29520
rect 8680 29306 8708 29514
rect 8668 29300 8720 29306
rect 8668 29242 8720 29248
rect 8484 28552 8536 28558
rect 8484 28494 8536 28500
rect 8392 28416 8444 28422
rect 8392 28358 8444 28364
rect 8208 28212 8260 28218
rect 8208 28154 8260 28160
rect 8404 28082 8432 28358
rect 8392 28076 8444 28082
rect 8392 28018 8444 28024
rect 6736 27464 6788 27470
rect 6736 27406 6788 27412
rect 7196 27464 7248 27470
rect 7196 27406 7248 27412
rect 6748 27062 6776 27406
rect 7840 27328 7892 27334
rect 7840 27270 7892 27276
rect 6736 27056 6788 27062
rect 6736 26998 6788 27004
rect 6748 25294 6776 26998
rect 7748 26784 7800 26790
rect 7748 26726 7800 26732
rect 7760 26450 7788 26726
rect 7748 26444 7800 26450
rect 7748 26386 7800 26392
rect 7288 26240 7340 26246
rect 7288 26182 7340 26188
rect 7300 25906 7328 26182
rect 7760 26042 7788 26386
rect 7748 26036 7800 26042
rect 7748 25978 7800 25984
rect 7852 25906 7880 27270
rect 8300 26920 8352 26926
rect 8300 26862 8352 26868
rect 7288 25900 7340 25906
rect 7288 25842 7340 25848
rect 7840 25900 7892 25906
rect 7840 25842 7892 25848
rect 8312 25498 8340 26862
rect 8300 25492 8352 25498
rect 8300 25434 8352 25440
rect 6736 25288 6788 25294
rect 6736 25230 6788 25236
rect 6276 24812 6328 24818
rect 6276 24754 6328 24760
rect 8392 24608 8444 24614
rect 8392 24550 8444 24556
rect 6368 24200 6420 24206
rect 6368 24142 6420 24148
rect 7748 24200 7800 24206
rect 7748 24142 7800 24148
rect 6380 22098 6408 24142
rect 7288 24132 7340 24138
rect 7288 24074 7340 24080
rect 6460 23112 6512 23118
rect 6460 23054 6512 23060
rect 6368 22092 6420 22098
rect 6368 22034 6420 22040
rect 6276 17672 6328 17678
rect 6276 17614 6328 17620
rect 6288 16250 6316 17614
rect 6368 16584 6420 16590
rect 6368 16526 6420 16532
rect 6276 16244 6328 16250
rect 6276 16186 6328 16192
rect 6380 16114 6408 16526
rect 6368 16108 6420 16114
rect 6368 16050 6420 16056
rect 6276 15972 6328 15978
rect 6276 15914 6328 15920
rect 6288 15638 6316 15914
rect 6276 15632 6328 15638
rect 6276 15574 6328 15580
rect 6472 15366 6500 23054
rect 7300 21962 7328 24074
rect 7760 23322 7788 24142
rect 8208 24064 8260 24070
rect 8208 24006 8260 24012
rect 8220 23866 8248 24006
rect 8208 23860 8260 23866
rect 8208 23802 8260 23808
rect 7748 23316 7800 23322
rect 7748 23258 7800 23264
rect 8116 22500 8168 22506
rect 8116 22442 8168 22448
rect 7104 21956 7156 21962
rect 7104 21898 7156 21904
rect 7288 21956 7340 21962
rect 7288 21898 7340 21904
rect 7116 21690 7144 21898
rect 7104 21684 7156 21690
rect 7104 21626 7156 21632
rect 7012 21548 7064 21554
rect 7012 21490 7064 21496
rect 7024 21146 7052 21490
rect 7012 21140 7064 21146
rect 7012 21082 7064 21088
rect 7300 19922 7328 21898
rect 7932 21480 7984 21486
rect 7932 21422 7984 21428
rect 7944 21010 7972 21422
rect 7932 21004 7984 21010
rect 7932 20946 7984 20952
rect 7656 20936 7708 20942
rect 7656 20878 7708 20884
rect 7668 20466 7696 20878
rect 8128 20806 8156 22442
rect 8300 21888 8352 21894
rect 8300 21830 8352 21836
rect 8312 20874 8340 21830
rect 8300 20868 8352 20874
rect 8300 20810 8352 20816
rect 8116 20800 8168 20806
rect 8116 20742 8168 20748
rect 8128 20534 8156 20742
rect 8116 20528 8168 20534
rect 8116 20470 8168 20476
rect 7656 20460 7708 20466
rect 7656 20402 7708 20408
rect 7288 19916 7340 19922
rect 7288 19858 7340 19864
rect 7288 19712 7340 19718
rect 7288 19654 7340 19660
rect 6828 19440 6880 19446
rect 6828 19382 6880 19388
rect 6840 18154 6868 19382
rect 6920 18760 6972 18766
rect 6920 18702 6972 18708
rect 7104 18760 7156 18766
rect 7104 18702 7156 18708
rect 6932 18426 6960 18702
rect 6920 18420 6972 18426
rect 6920 18362 6972 18368
rect 6828 18148 6880 18154
rect 6828 18090 6880 18096
rect 7116 17338 7144 18702
rect 7300 18290 7328 19654
rect 7564 18624 7616 18630
rect 7564 18566 7616 18572
rect 7380 18352 7432 18358
rect 7380 18294 7432 18300
rect 7288 18284 7340 18290
rect 7288 18226 7340 18232
rect 7104 17332 7156 17338
rect 7104 17274 7156 17280
rect 6552 17060 6604 17066
rect 6552 17002 6604 17008
rect 6460 15360 6512 15366
rect 6460 15302 6512 15308
rect 6184 14000 6236 14006
rect 6184 13942 6236 13948
rect 6460 13184 6512 13190
rect 6460 13126 6512 13132
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 6276 12232 6328 12238
rect 6276 12174 6328 12180
rect 6184 12096 6236 12102
rect 6184 12038 6236 12044
rect 6196 11898 6224 12038
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 6184 11280 6236 11286
rect 6184 11222 6236 11228
rect 6196 11150 6224 11222
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 6092 10736 6144 10742
rect 6092 10678 6144 10684
rect 5960 9948 6040 9976
rect 6092 9988 6144 9994
rect 5908 9930 5960 9936
rect 6092 9930 6144 9936
rect 5920 9081 5948 9930
rect 5906 9072 5962 9081
rect 5906 9007 5962 9016
rect 5816 8424 5868 8430
rect 5816 8366 5868 8372
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5368 6718 5488 6746
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 3976 5646 4028 5652
rect 5170 5672 5226 5681
rect 3988 5302 4016 5646
rect 5170 5607 5226 5616
rect 3976 5296 4028 5302
rect 3976 5238 4028 5244
rect 3988 4622 4016 5238
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 5368 4865 5396 6258
rect 5460 5098 5488 6718
rect 5724 6180 5776 6186
rect 5724 6122 5776 6128
rect 5448 5092 5500 5098
rect 5448 5034 5500 5040
rect 5354 4856 5410 4865
rect 5354 4791 5410 4800
rect 3976 4616 4028 4622
rect 4028 4564 4108 4570
rect 3976 4558 4108 4564
rect 3988 4542 4108 4558
rect 4080 3602 4108 4542
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 4080 3058 4108 3538
rect 3332 3052 3384 3058
rect 3332 2994 3384 3000
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 3344 2961 3372 2994
rect 3330 2952 3386 2961
rect 3330 2887 3386 2896
rect 4080 2774 4108 2994
rect 5460 2990 5488 5034
rect 5736 4690 5764 6122
rect 5724 4684 5776 4690
rect 5724 4626 5776 4632
rect 5828 4146 5856 8366
rect 5920 6254 5948 9007
rect 6000 8900 6052 8906
rect 6000 8842 6052 8848
rect 6012 7954 6040 8842
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 6104 7546 6132 9930
rect 6092 7540 6144 7546
rect 6092 7482 6144 7488
rect 5908 6248 5960 6254
rect 5908 6190 5960 6196
rect 6196 5914 6224 11086
rect 6184 5908 6236 5914
rect 6184 5850 6236 5856
rect 6288 5098 6316 12174
rect 6380 8498 6408 12242
rect 6472 8906 6500 13126
rect 6564 10810 6592 17002
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 6736 15904 6788 15910
rect 6736 15846 6788 15852
rect 6748 15434 6776 15846
rect 6736 15428 6788 15434
rect 6736 15370 6788 15376
rect 6748 13530 6776 15370
rect 6736 13524 6788 13530
rect 6736 13466 6788 13472
rect 6840 12918 6868 16934
rect 7392 16590 7420 18294
rect 7576 18222 7604 18566
rect 7564 18216 7616 18222
rect 7564 18158 7616 18164
rect 7196 16584 7248 16590
rect 7196 16526 7248 16532
rect 7380 16584 7432 16590
rect 7380 16526 7432 16532
rect 6828 12912 6880 12918
rect 6828 12854 6880 12860
rect 7208 12238 7236 16526
rect 7380 16040 7432 16046
rect 7380 15982 7432 15988
rect 7392 12918 7420 15982
rect 7472 14340 7524 14346
rect 7472 14282 7524 14288
rect 7380 12912 7432 12918
rect 7380 12854 7432 12860
rect 7392 12442 7420 12854
rect 7380 12436 7432 12442
rect 7380 12378 7432 12384
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 6736 11008 6788 11014
rect 6736 10950 6788 10956
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 6748 10742 6776 10950
rect 6736 10736 6788 10742
rect 6736 10678 6788 10684
rect 7012 10600 7064 10606
rect 7012 10542 7064 10548
rect 6644 10532 6696 10538
rect 6644 10474 6696 10480
rect 6552 9512 6604 9518
rect 6552 9454 6604 9460
rect 6460 8900 6512 8906
rect 6460 8842 6512 8848
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 6564 7886 6592 9454
rect 6656 9042 6684 10474
rect 7024 9178 7052 10542
rect 7012 9172 7064 9178
rect 7012 9114 7064 9120
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6564 7478 6592 7822
rect 6552 7472 6604 7478
rect 6552 7414 6604 7420
rect 6564 6882 6592 7414
rect 6472 6866 6592 6882
rect 6460 6860 6592 6866
rect 6512 6854 6592 6860
rect 6460 6802 6512 6808
rect 7024 5370 7052 9114
rect 7208 6186 7236 12174
rect 7196 6180 7248 6186
rect 7196 6122 7248 6128
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 6276 5092 6328 5098
rect 6276 5034 6328 5040
rect 5908 4548 5960 4554
rect 5908 4490 5960 4496
rect 5920 4282 5948 4490
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 5908 4276 5960 4282
rect 5908 4218 5960 4224
rect 7300 4146 7328 4422
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 5828 3194 5856 4082
rect 7196 3596 7248 3602
rect 7196 3538 7248 3544
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 6644 3120 6696 3126
rect 6644 3062 6696 3068
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 3988 2746 4108 2774
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 3988 2514 4016 2746
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 2872 2508 2924 2514
rect 2872 2450 2924 2456
rect 3976 2508 4028 2514
rect 3976 2450 4028 2456
rect 5828 2446 5856 2790
rect 6656 2446 6684 3062
rect 7208 2990 7236 3538
rect 7196 2984 7248 2990
rect 7196 2926 7248 2932
rect 7208 2774 7236 2926
rect 7116 2746 7236 2774
rect 7012 2576 7064 2582
rect 7012 2518 7064 2524
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 2778 1456 2834 1465
rect 2778 1391 2834 1400
rect 4540 800 4568 2246
rect 5828 800 5856 2246
rect 7024 2106 7052 2518
rect 7012 2100 7064 2106
rect 7012 2042 7064 2048
rect 7116 800 7144 2746
rect 7392 2650 7420 4082
rect 7484 3738 7512 14282
rect 7668 11286 7696 20402
rect 8024 18760 8076 18766
rect 8024 18702 8076 18708
rect 7748 17672 7800 17678
rect 7748 17614 7800 17620
rect 7932 17672 7984 17678
rect 7932 17614 7984 17620
rect 7760 13326 7788 17614
rect 7944 16726 7972 17614
rect 8036 17066 8064 18702
rect 8300 17808 8352 17814
rect 8300 17750 8352 17756
rect 8312 17610 8340 17750
rect 8300 17604 8352 17610
rect 8300 17546 8352 17552
rect 8300 17264 8352 17270
rect 8300 17206 8352 17212
rect 8312 17082 8340 17206
rect 8404 17202 8432 24550
rect 8392 17196 8444 17202
rect 8392 17138 8444 17144
rect 8024 17060 8076 17066
rect 8312 17054 8432 17082
rect 8024 17002 8076 17008
rect 7932 16720 7984 16726
rect 7932 16662 7984 16668
rect 8036 16658 8064 17002
rect 8404 16998 8432 17054
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 8392 16992 8444 16998
rect 8392 16934 8444 16940
rect 8024 16652 8076 16658
rect 8024 16594 8076 16600
rect 8116 16516 8168 16522
rect 8116 16458 8168 16464
rect 8128 15502 8156 16458
rect 8116 15496 8168 15502
rect 8116 15438 8168 15444
rect 7748 13320 7800 13326
rect 7748 13262 7800 13268
rect 8312 11898 8340 16934
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 7932 11824 7984 11830
rect 8496 11778 8524 28494
rect 8956 28082 8984 37062
rect 10692 36916 10744 36922
rect 10692 36858 10744 36864
rect 10600 31816 10652 31822
rect 10600 31758 10652 31764
rect 10612 30326 10640 31758
rect 10600 30320 10652 30326
rect 10600 30262 10652 30268
rect 10140 29572 10192 29578
rect 10140 29514 10192 29520
rect 10152 29306 10180 29514
rect 10140 29300 10192 29306
rect 10140 29242 10192 29248
rect 10704 28558 10732 36858
rect 11256 33114 11284 37198
rect 11244 33108 11296 33114
rect 11244 33050 11296 33056
rect 11716 32570 11744 37198
rect 12268 37108 12296 39200
rect 13556 37262 13584 39200
rect 13544 37256 13596 37262
rect 13544 37198 13596 37204
rect 13728 37188 13780 37194
rect 13728 37130 13780 37136
rect 12440 37120 12492 37126
rect 12268 37080 12440 37108
rect 12440 37062 12492 37068
rect 12532 32904 12584 32910
rect 12532 32846 12584 32852
rect 11704 32564 11756 32570
rect 11704 32506 11756 32512
rect 11888 32428 11940 32434
rect 11888 32370 11940 32376
rect 11244 30728 11296 30734
rect 11244 30670 11296 30676
rect 10784 29640 10836 29646
rect 10784 29582 10836 29588
rect 10232 28552 10284 28558
rect 10232 28494 10284 28500
rect 10692 28552 10744 28558
rect 10692 28494 10744 28500
rect 10048 28416 10100 28422
rect 10048 28358 10100 28364
rect 10060 28082 10088 28358
rect 8944 28076 8996 28082
rect 8944 28018 8996 28024
rect 10048 28076 10100 28082
rect 10048 28018 10100 28024
rect 9864 28008 9916 28014
rect 9864 27950 9916 27956
rect 9876 27674 9904 27950
rect 9864 27668 9916 27674
rect 9864 27610 9916 27616
rect 8944 27396 8996 27402
rect 8944 27338 8996 27344
rect 8956 25974 8984 27338
rect 9128 27328 9180 27334
rect 9128 27270 9180 27276
rect 9140 26994 9168 27270
rect 9128 26988 9180 26994
rect 9128 26930 9180 26936
rect 10244 26858 10272 28494
rect 10508 27872 10560 27878
rect 10508 27814 10560 27820
rect 10520 27606 10548 27814
rect 10508 27600 10560 27606
rect 10508 27542 10560 27548
rect 10796 27470 10824 29582
rect 11256 29170 11284 30670
rect 11900 29850 11928 32370
rect 11980 30592 12032 30598
rect 11980 30534 12032 30540
rect 11888 29844 11940 29850
rect 11888 29786 11940 29792
rect 11992 29578 12020 30534
rect 12544 30326 12572 32846
rect 13740 30938 13768 37130
rect 15488 37126 15516 39200
rect 15568 37256 15620 37262
rect 15568 37198 15620 37204
rect 14280 37120 14332 37126
rect 14280 37062 14332 37068
rect 15476 37120 15528 37126
rect 15476 37062 15528 37068
rect 14096 35080 14148 35086
rect 14096 35022 14148 35028
rect 13728 30932 13780 30938
rect 13728 30874 13780 30880
rect 14108 30326 14136 35022
rect 14292 31958 14320 37062
rect 15580 36922 15608 37198
rect 16776 37126 16804 39200
rect 18064 37262 18092 39200
rect 16856 37256 16908 37262
rect 16856 37198 16908 37204
rect 18052 37256 18104 37262
rect 18052 37198 18104 37204
rect 16764 37120 16816 37126
rect 16764 37062 16816 37068
rect 15568 36916 15620 36922
rect 15568 36858 15620 36864
rect 16868 32026 16896 37198
rect 17500 37188 17552 37194
rect 17500 37130 17552 37136
rect 17512 32570 17540 37130
rect 19996 37126 20024 39200
rect 21284 37126 21312 39200
rect 22572 37262 22600 39200
rect 24504 37262 24532 39200
rect 25792 37262 25820 39200
rect 22008 37256 22060 37262
rect 22008 37198 22060 37204
rect 22560 37256 22612 37262
rect 22560 37198 22612 37204
rect 24492 37256 24544 37262
rect 24492 37198 24544 37204
rect 25780 37256 25832 37262
rect 25780 37198 25832 37204
rect 17960 37120 18012 37126
rect 17960 37062 18012 37068
rect 19984 37120 20036 37126
rect 19984 37062 20036 37068
rect 21272 37120 21324 37126
rect 21272 37062 21324 37068
rect 17500 32564 17552 32570
rect 17500 32506 17552 32512
rect 16948 32428 17000 32434
rect 16948 32370 17000 32376
rect 16856 32020 16908 32026
rect 16856 31962 16908 31968
rect 14280 31952 14332 31958
rect 14280 31894 14332 31900
rect 15568 31340 15620 31346
rect 15568 31282 15620 31288
rect 15292 31136 15344 31142
rect 15292 31078 15344 31084
rect 14464 30728 14516 30734
rect 14464 30670 14516 30676
rect 14476 30394 14504 30670
rect 14464 30388 14516 30394
rect 14464 30330 14516 30336
rect 12532 30320 12584 30326
rect 12532 30262 12584 30268
rect 14096 30320 14148 30326
rect 14096 30262 14148 30268
rect 12256 30252 12308 30258
rect 12256 30194 12308 30200
rect 12440 30252 12492 30258
rect 12440 30194 12492 30200
rect 14188 30252 14240 30258
rect 14188 30194 14240 30200
rect 15016 30252 15068 30258
rect 15016 30194 15068 30200
rect 11888 29572 11940 29578
rect 11888 29514 11940 29520
rect 11980 29572 12032 29578
rect 11980 29514 12032 29520
rect 11900 29306 11928 29514
rect 11888 29300 11940 29306
rect 11888 29242 11940 29248
rect 11244 29164 11296 29170
rect 11244 29106 11296 29112
rect 10324 27464 10376 27470
rect 10324 27406 10376 27412
rect 10784 27464 10836 27470
rect 10784 27406 10836 27412
rect 10336 27062 10364 27406
rect 10324 27056 10376 27062
rect 10324 26998 10376 27004
rect 10232 26852 10284 26858
rect 10232 26794 10284 26800
rect 9312 26784 9364 26790
rect 9312 26726 9364 26732
rect 9324 26450 9352 26726
rect 10796 26586 10824 27406
rect 10784 26580 10836 26586
rect 10784 26522 10836 26528
rect 9312 26444 9364 26450
rect 9312 26386 9364 26392
rect 8944 25968 8996 25974
rect 8944 25910 8996 25916
rect 9772 25968 9824 25974
rect 9772 25910 9824 25916
rect 9784 25498 9812 25910
rect 10968 25696 11020 25702
rect 10968 25638 11020 25644
rect 9772 25492 9824 25498
rect 9772 25434 9824 25440
rect 9956 25288 10008 25294
rect 9956 25230 10008 25236
rect 9968 24954 9996 25230
rect 9956 24948 10008 24954
rect 9956 24890 10008 24896
rect 10784 24812 10836 24818
rect 10784 24754 10836 24760
rect 10796 24206 10824 24754
rect 10784 24200 10836 24206
rect 10784 24142 10836 24148
rect 10508 24064 10560 24070
rect 10508 24006 10560 24012
rect 10520 23730 10548 24006
rect 9220 23724 9272 23730
rect 9220 23666 9272 23672
rect 10508 23724 10560 23730
rect 10508 23666 10560 23672
rect 8852 22704 8904 22710
rect 8852 22646 8904 22652
rect 8864 22234 8892 22646
rect 8852 22228 8904 22234
rect 8852 22170 8904 22176
rect 8668 22024 8720 22030
rect 8668 21966 8720 21972
rect 8680 21690 8708 21966
rect 8668 21684 8720 21690
rect 8668 21626 8720 21632
rect 8668 21412 8720 21418
rect 8668 21354 8720 21360
rect 8680 20330 8708 21354
rect 9232 21146 9260 23666
rect 9404 23248 9456 23254
rect 9404 23190 9456 23196
rect 9416 22710 9444 23190
rect 9404 22704 9456 22710
rect 9404 22646 9456 22652
rect 10140 22568 10192 22574
rect 10140 22510 10192 22516
rect 10152 22098 10180 22510
rect 9956 22092 10008 22098
rect 9956 22034 10008 22040
rect 10140 22092 10192 22098
rect 10140 22034 10192 22040
rect 9968 21894 9996 22034
rect 9956 21888 10008 21894
rect 9956 21830 10008 21836
rect 9864 21616 9916 21622
rect 9864 21558 9916 21564
rect 9588 21548 9640 21554
rect 9588 21490 9640 21496
rect 9220 21140 9272 21146
rect 9220 21082 9272 21088
rect 8668 20324 8720 20330
rect 8668 20266 8720 20272
rect 8576 16244 8628 16250
rect 8576 16186 8628 16192
rect 8588 15706 8616 16186
rect 8680 16182 8708 20266
rect 9312 20256 9364 20262
rect 9312 20198 9364 20204
rect 9324 19854 9352 20198
rect 9312 19848 9364 19854
rect 9312 19790 9364 19796
rect 9404 18896 9456 18902
rect 9404 18838 9456 18844
rect 9220 18624 9272 18630
rect 9220 18566 9272 18572
rect 9232 17746 9260 18566
rect 9416 18358 9444 18838
rect 9404 18352 9456 18358
rect 9404 18294 9456 18300
rect 9220 17740 9272 17746
rect 9220 17682 9272 17688
rect 9036 17264 9088 17270
rect 9036 17206 9088 17212
rect 9048 16794 9076 17206
rect 9036 16788 9088 16794
rect 9036 16730 9088 16736
rect 9404 16448 9456 16454
rect 9404 16390 9456 16396
rect 9496 16448 9548 16454
rect 9496 16390 9548 16396
rect 8668 16176 8720 16182
rect 8668 16118 8720 16124
rect 8576 15700 8628 15706
rect 8576 15642 8628 15648
rect 8668 15700 8720 15706
rect 8668 15642 8720 15648
rect 8588 15094 8616 15642
rect 8680 15366 8708 15642
rect 8760 15564 8812 15570
rect 8760 15506 8812 15512
rect 8668 15360 8720 15366
rect 8668 15302 8720 15308
rect 8576 15088 8628 15094
rect 8576 15030 8628 15036
rect 8772 15026 8800 15506
rect 8760 15020 8812 15026
rect 8760 14962 8812 14968
rect 8772 14074 8800 14962
rect 8760 14068 8812 14074
rect 8760 14010 8812 14016
rect 8772 12866 8800 14010
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 8680 12850 8800 12866
rect 8668 12844 8800 12850
rect 8720 12838 8800 12844
rect 8668 12786 8720 12792
rect 8772 12458 8800 12838
rect 9036 12776 9088 12782
rect 9036 12718 9088 12724
rect 9048 12646 9076 12718
rect 9140 12646 9168 13262
rect 9416 12918 9444 16390
rect 9508 15978 9536 16390
rect 9496 15972 9548 15978
rect 9496 15914 9548 15920
rect 9404 12912 9456 12918
rect 9404 12854 9456 12860
rect 9036 12640 9088 12646
rect 9036 12582 9088 12588
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 7932 11766 7984 11772
rect 7656 11280 7708 11286
rect 7656 11222 7708 11228
rect 7668 9518 7696 11222
rect 7944 10810 7972 11766
rect 8312 11750 8524 11778
rect 8680 12430 8800 12458
rect 9600 12434 9628 21490
rect 9876 21146 9904 21558
rect 9864 21140 9916 21146
rect 9864 21082 9916 21088
rect 10048 20936 10100 20942
rect 10048 20878 10100 20884
rect 9772 20528 9824 20534
rect 9772 20470 9824 20476
rect 9784 19514 9812 20470
rect 10060 20058 10088 20878
rect 10048 20052 10100 20058
rect 10048 19994 10100 20000
rect 9956 19848 10008 19854
rect 9956 19790 10008 19796
rect 9772 19508 9824 19514
rect 9772 19450 9824 19456
rect 9968 19378 9996 19790
rect 10508 19780 10560 19786
rect 10508 19722 10560 19728
rect 9956 19372 10008 19378
rect 9956 19314 10008 19320
rect 10232 18352 10284 18358
rect 10232 18294 10284 18300
rect 10048 18284 10100 18290
rect 10048 18226 10100 18232
rect 10060 17882 10088 18226
rect 10048 17876 10100 17882
rect 10048 17818 10100 17824
rect 9864 17604 9916 17610
rect 9864 17546 9916 17552
rect 9876 17134 9904 17546
rect 9864 17128 9916 17134
rect 9864 17070 9916 17076
rect 8312 11694 8340 11750
rect 8300 11688 8352 11694
rect 8300 11630 8352 11636
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 8024 9444 8076 9450
rect 8024 9386 8076 9392
rect 8036 9178 8064 9386
rect 8128 9178 8156 9522
rect 8312 9518 8340 11630
rect 8680 11558 8708 12430
rect 9508 12406 9628 12434
rect 9220 12300 9272 12306
rect 9220 12242 9272 12248
rect 9128 12164 9180 12170
rect 9128 12106 9180 12112
rect 9140 11694 9168 12106
rect 9232 11694 9260 12242
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 9220 11688 9272 11694
rect 9220 11630 9272 11636
rect 8760 11620 8812 11626
rect 8760 11562 8812 11568
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8772 11150 8800 11562
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 9140 11150 9168 11494
rect 8760 11144 8812 11150
rect 8760 11086 8812 11092
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 8116 9172 8168 9178
rect 8116 9114 8168 9120
rect 8116 8900 8168 8906
rect 8116 8842 8168 8848
rect 8128 8566 8156 8842
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8116 8560 8168 8566
rect 8116 8502 8168 8508
rect 8312 7562 8340 8570
rect 8220 7546 8340 7562
rect 8208 7540 8340 7546
rect 8260 7534 8340 7540
rect 8208 7482 8260 7488
rect 7840 7336 7892 7342
rect 7840 7278 7892 7284
rect 7852 6662 7880 7278
rect 7840 6656 7892 6662
rect 7840 6598 7892 6604
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 7484 3126 7512 3674
rect 7852 3466 7880 6598
rect 7944 6458 7972 6598
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 8404 4146 8432 10542
rect 9140 9518 9168 11086
rect 9324 11082 9352 11834
rect 9312 11076 9364 11082
rect 9312 11018 9364 11024
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 8484 9104 8536 9110
rect 8484 9046 8536 9052
rect 8496 8566 8524 9046
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8484 8560 8536 8566
rect 8484 8502 8536 8508
rect 8588 8430 8616 8774
rect 9140 8650 9168 9454
rect 9140 8634 9260 8650
rect 9140 8628 9272 8634
rect 9140 8622 9220 8628
rect 9220 8570 9272 8576
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8484 7812 8536 7818
rect 8484 7754 8536 7760
rect 8496 7546 8524 7754
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8484 7540 8536 7546
rect 8484 7482 8536 7488
rect 8680 5778 8708 7686
rect 9232 6798 9260 8570
rect 9324 7478 9352 9862
rect 9312 7472 9364 7478
rect 9312 7414 9364 7420
rect 9404 7472 9456 7478
rect 9404 7414 9456 7420
rect 9416 7002 9444 7414
rect 9404 6996 9456 7002
rect 9404 6938 9456 6944
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9128 6112 9180 6118
rect 9232 6066 9260 6734
rect 9508 6254 9536 12406
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9600 11286 9628 11494
rect 9588 11280 9640 11286
rect 9588 11222 9640 11228
rect 9876 10538 9904 17070
rect 10244 16998 10272 18294
rect 10520 17814 10548 19722
rect 10692 19372 10744 19378
rect 10692 19314 10744 19320
rect 10416 17808 10468 17814
rect 10416 17750 10468 17756
rect 10508 17808 10560 17814
rect 10508 17750 10560 17756
rect 10232 16992 10284 16998
rect 10232 16934 10284 16940
rect 10140 13728 10192 13734
rect 10140 13670 10192 13676
rect 10152 13394 10180 13670
rect 10140 13388 10192 13394
rect 10140 13330 10192 13336
rect 9864 10532 9916 10538
rect 9864 10474 9916 10480
rect 10152 8634 10180 13330
rect 10244 12850 10272 16934
rect 10324 16108 10376 16114
rect 10324 16050 10376 16056
rect 10336 14414 10364 16050
rect 10324 14408 10376 14414
rect 10324 14350 10376 14356
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 9600 7342 9628 8434
rect 10336 8090 10364 14350
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 10324 8084 10376 8090
rect 10324 8026 10376 8032
rect 9588 7336 9640 7342
rect 9588 7278 9640 7284
rect 9588 6724 9640 6730
rect 9588 6666 9640 6672
rect 9600 6254 9628 6666
rect 9496 6248 9548 6254
rect 9496 6190 9548 6196
rect 9588 6248 9640 6254
rect 9588 6190 9640 6196
rect 9180 6060 9260 6066
rect 9128 6054 9260 6060
rect 9312 6112 9364 6118
rect 9312 6054 9364 6060
rect 9140 6038 9260 6054
rect 8668 5772 8720 5778
rect 8668 5714 8720 5720
rect 9232 5710 9260 6038
rect 9324 5846 9352 6054
rect 9312 5840 9364 5846
rect 9312 5782 9364 5788
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9232 5234 9260 5646
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 9048 3466 9076 3674
rect 7840 3460 7892 3466
rect 7840 3402 7892 3408
rect 9036 3460 9088 3466
rect 9036 3402 9088 3408
rect 7472 3120 7524 3126
rect 7472 3062 7524 3068
rect 9128 3052 9180 3058
rect 9232 3040 9260 5170
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9692 3126 9720 4626
rect 9680 3120 9732 3126
rect 9680 3062 9732 3068
rect 9180 3012 9260 3040
rect 9128 2994 9180 3000
rect 10060 2990 10088 8026
rect 10428 6458 10456 17750
rect 10508 16176 10560 16182
rect 10506 16144 10508 16153
rect 10560 16144 10562 16153
rect 10506 16079 10562 16088
rect 10508 15904 10560 15910
rect 10508 15846 10560 15852
rect 10520 15502 10548 15846
rect 10508 15496 10560 15502
rect 10508 15438 10560 15444
rect 10704 13138 10732 19314
rect 10796 15638 10824 24142
rect 10980 23730 11008 25638
rect 10968 23724 11020 23730
rect 10968 23666 11020 23672
rect 10876 22024 10928 22030
rect 10876 21966 10928 21972
rect 10888 21690 10916 21966
rect 10876 21684 10928 21690
rect 10876 21626 10928 21632
rect 11060 21548 11112 21554
rect 11060 21490 11112 21496
rect 11072 20602 11100 21490
rect 11152 21480 11204 21486
rect 11152 21422 11204 21428
rect 11060 20596 11112 20602
rect 11060 20538 11112 20544
rect 11164 20330 11192 21422
rect 11152 20324 11204 20330
rect 11152 20266 11204 20272
rect 11060 18216 11112 18222
rect 11060 18158 11112 18164
rect 11072 17882 11100 18158
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 11060 17740 11112 17746
rect 11060 17682 11112 17688
rect 10876 17672 10928 17678
rect 10876 17614 10928 17620
rect 10888 17338 10916 17614
rect 10876 17332 10928 17338
rect 10876 17274 10928 17280
rect 10876 16992 10928 16998
rect 10876 16934 10928 16940
rect 10784 15632 10836 15638
rect 10784 15574 10836 15580
rect 10796 13258 10824 15574
rect 10784 13252 10836 13258
rect 10784 13194 10836 13200
rect 10704 13110 10824 13138
rect 10600 12844 10652 12850
rect 10600 12786 10652 12792
rect 10508 12436 10560 12442
rect 10508 12378 10560 12384
rect 10520 11830 10548 12378
rect 10508 11824 10560 11830
rect 10508 11766 10560 11772
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10520 8634 10548 9522
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10612 7750 10640 12786
rect 10600 7744 10652 7750
rect 10600 7686 10652 7692
rect 10508 6860 10560 6866
rect 10508 6802 10560 6808
rect 10520 6458 10548 6802
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 10048 2984 10100 2990
rect 10048 2926 10100 2932
rect 10152 2854 10180 3674
rect 10140 2848 10192 2854
rect 10140 2790 10192 2796
rect 10428 2774 10456 6394
rect 10692 6180 10744 6186
rect 10692 6122 10744 6128
rect 10704 5030 10732 6122
rect 10796 5166 10824 13110
rect 10888 10198 10916 16934
rect 10966 16144 11022 16153
rect 10966 16079 11022 16088
rect 10980 16046 11008 16079
rect 10968 16040 11020 16046
rect 10968 15982 11020 15988
rect 10968 15088 11020 15094
rect 10968 15030 11020 15036
rect 10980 11234 11008 15030
rect 11072 12782 11100 17682
rect 11152 16176 11204 16182
rect 11152 16118 11204 16124
rect 11164 14618 11192 16118
rect 11152 14612 11204 14618
rect 11152 14554 11204 14560
rect 11060 12776 11112 12782
rect 11060 12718 11112 12724
rect 11072 12306 11100 12718
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 11256 12170 11284 29106
rect 11704 28416 11756 28422
rect 11704 28358 11756 28364
rect 11520 27532 11572 27538
rect 11520 27474 11572 27480
rect 11428 27464 11480 27470
rect 11428 27406 11480 27412
rect 11440 27130 11468 27406
rect 11428 27124 11480 27130
rect 11428 27066 11480 27072
rect 11532 26994 11560 27474
rect 11520 26988 11572 26994
rect 11520 26930 11572 26936
rect 11532 26234 11560 26930
rect 11440 26206 11560 26234
rect 11336 22976 11388 22982
rect 11336 22918 11388 22924
rect 11348 17746 11376 22918
rect 11336 17740 11388 17746
rect 11336 17682 11388 17688
rect 11336 16244 11388 16250
rect 11336 16186 11388 16192
rect 11348 15706 11376 16186
rect 11336 15700 11388 15706
rect 11336 15642 11388 15648
rect 11440 13802 11468 26206
rect 11716 25906 11744 28358
rect 11520 25900 11572 25906
rect 11520 25842 11572 25848
rect 11704 25900 11756 25906
rect 11704 25842 11756 25848
rect 11532 25498 11560 25842
rect 11520 25492 11572 25498
rect 11520 25434 11572 25440
rect 11704 25288 11756 25294
rect 11704 25230 11756 25236
rect 11716 23322 11744 25230
rect 12164 23656 12216 23662
rect 12164 23598 12216 23604
rect 11704 23316 11756 23322
rect 11704 23258 11756 23264
rect 11716 23118 11744 23258
rect 12176 23186 12204 23598
rect 12164 23180 12216 23186
rect 12164 23122 12216 23128
rect 11704 23112 11756 23118
rect 11704 23054 11756 23060
rect 11888 22704 11940 22710
rect 11888 22646 11940 22652
rect 11796 22568 11848 22574
rect 11796 22510 11848 22516
rect 11808 22098 11836 22510
rect 11796 22092 11848 22098
rect 11796 22034 11848 22040
rect 11900 21690 11928 22646
rect 12268 22574 12296 30194
rect 12452 28762 12480 30194
rect 14200 29850 14228 30194
rect 14188 29844 14240 29850
rect 14188 29786 14240 29792
rect 15028 29186 15056 30194
rect 15108 29844 15160 29850
rect 15108 29786 15160 29792
rect 15120 29306 15148 29786
rect 15304 29714 15332 31078
rect 15292 29708 15344 29714
rect 15292 29650 15344 29656
rect 15580 29646 15608 31282
rect 16960 30326 16988 32370
rect 17040 31816 17092 31822
rect 17040 31758 17092 31764
rect 17052 30938 17080 31758
rect 17040 30932 17092 30938
rect 17040 30874 17092 30880
rect 16948 30320 17000 30326
rect 16948 30262 17000 30268
rect 16856 30252 16908 30258
rect 16856 30194 16908 30200
rect 16868 29782 16896 30194
rect 16856 29776 16908 29782
rect 16856 29718 16908 29724
rect 15568 29640 15620 29646
rect 15568 29582 15620 29588
rect 15108 29300 15160 29306
rect 15108 29242 15160 29248
rect 15028 29158 15148 29186
rect 12440 28756 12492 28762
rect 12440 28698 12492 28704
rect 13268 28756 13320 28762
rect 13268 28698 13320 28704
rect 13452 28756 13504 28762
rect 13452 28698 13504 28704
rect 12900 28552 12952 28558
rect 12900 28494 12952 28500
rect 12912 28218 12940 28494
rect 13280 28218 13308 28698
rect 12900 28212 12952 28218
rect 12900 28154 12952 28160
rect 13268 28212 13320 28218
rect 13268 28154 13320 28160
rect 12624 28008 12676 28014
rect 12624 27950 12676 27956
rect 12636 27538 12664 27950
rect 12624 27532 12676 27538
rect 12624 27474 12676 27480
rect 13268 27328 13320 27334
rect 13268 27270 13320 27276
rect 13280 27062 13308 27270
rect 13268 27056 13320 27062
rect 13268 26998 13320 27004
rect 12900 26580 12952 26586
rect 12900 26522 12952 26528
rect 12716 25832 12768 25838
rect 12716 25774 12768 25780
rect 12728 25362 12756 25774
rect 12912 25362 12940 26522
rect 13084 26376 13136 26382
rect 13084 26318 13136 26324
rect 12716 25356 12768 25362
rect 12716 25298 12768 25304
rect 12900 25356 12952 25362
rect 12900 25298 12952 25304
rect 12900 24812 12952 24818
rect 12900 24754 12952 24760
rect 12624 24744 12676 24750
rect 12624 24686 12676 24692
rect 12348 24064 12400 24070
rect 12348 24006 12400 24012
rect 12360 23730 12388 24006
rect 12348 23724 12400 23730
rect 12348 23666 12400 23672
rect 11980 22568 12032 22574
rect 11980 22510 12032 22516
rect 12256 22568 12308 22574
rect 12256 22510 12308 22516
rect 11888 21684 11940 21690
rect 11888 21626 11940 21632
rect 11992 19922 12020 22510
rect 12164 21888 12216 21894
rect 12164 21830 12216 21836
rect 12176 21690 12204 21830
rect 12164 21684 12216 21690
rect 12164 21626 12216 21632
rect 12256 21548 12308 21554
rect 12256 21490 12308 21496
rect 12268 20058 12296 21490
rect 12440 20936 12492 20942
rect 12440 20878 12492 20884
rect 12348 20460 12400 20466
rect 12348 20402 12400 20408
rect 12256 20052 12308 20058
rect 12256 19994 12308 20000
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 12360 19854 12388 20402
rect 12072 19848 12124 19854
rect 12072 19790 12124 19796
rect 12348 19848 12400 19854
rect 12348 19790 12400 19796
rect 11520 19372 11572 19378
rect 11520 19314 11572 19320
rect 11532 18766 11560 19314
rect 11978 19000 12034 19009
rect 11978 18935 12034 18944
rect 11520 18760 11572 18766
rect 11520 18702 11572 18708
rect 11532 15434 11560 18702
rect 11992 18698 12020 18935
rect 11980 18692 12032 18698
rect 11980 18634 12032 18640
rect 12084 18290 12112 19790
rect 12164 19780 12216 19786
rect 12164 19722 12216 19728
rect 12176 18426 12204 19722
rect 12164 18420 12216 18426
rect 12164 18362 12216 18368
rect 12072 18284 12124 18290
rect 12072 18226 12124 18232
rect 11980 18080 12032 18086
rect 11980 18022 12032 18028
rect 11992 17610 12020 18022
rect 11980 17604 12032 17610
rect 11980 17546 12032 17552
rect 11796 17536 11848 17542
rect 11796 17478 11848 17484
rect 11520 15428 11572 15434
rect 11520 15370 11572 15376
rect 11428 13796 11480 13802
rect 11428 13738 11480 13744
rect 11244 12164 11296 12170
rect 11244 12106 11296 12112
rect 11152 11620 11204 11626
rect 11152 11562 11204 11568
rect 10980 11218 11100 11234
rect 11164 11218 11192 11562
rect 11440 11354 11468 13738
rect 11532 12102 11560 15370
rect 11612 12640 11664 12646
rect 11610 12608 11612 12617
rect 11704 12640 11756 12646
rect 11664 12608 11666 12617
rect 11704 12582 11756 12588
rect 11610 12543 11666 12552
rect 11520 12096 11572 12102
rect 11520 12038 11572 12044
rect 11428 11348 11480 11354
rect 11428 11290 11480 11296
rect 10980 11212 11112 11218
rect 10980 11206 11060 11212
rect 11060 11154 11112 11160
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 11336 10668 11388 10674
rect 11336 10610 11388 10616
rect 10876 10192 10928 10198
rect 10876 10134 10928 10140
rect 11348 8974 11376 10610
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 11244 8900 11296 8906
rect 11244 8842 11296 8848
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 11072 7954 11100 8230
rect 11256 7993 11284 8842
rect 11348 8362 11376 8910
rect 11336 8356 11388 8362
rect 11336 8298 11388 8304
rect 11242 7984 11298 7993
rect 11060 7948 11112 7954
rect 11242 7919 11298 7928
rect 11060 7890 11112 7896
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10520 4078 10548 4558
rect 10508 4072 10560 4078
rect 10508 4014 10560 4020
rect 10336 2746 10456 2774
rect 10336 2650 10364 2746
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 7472 2644 7524 2650
rect 7472 2586 7524 2592
rect 10324 2644 10376 2650
rect 10324 2586 10376 2592
rect 7484 2530 7512 2586
rect 7208 2514 7512 2530
rect 7196 2508 7512 2514
rect 7248 2502 7512 2508
rect 7196 2450 7248 2456
rect 10796 2446 10824 5102
rect 11072 5030 11100 7142
rect 11164 5710 11192 7822
rect 11336 7812 11388 7818
rect 11336 7754 11388 7760
rect 11348 6934 11376 7754
rect 11336 6928 11388 6934
rect 11336 6870 11388 6876
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 11152 5296 11204 5302
rect 11152 5238 11204 5244
rect 11060 5024 11112 5030
rect 11060 4966 11112 4972
rect 11164 4593 11192 5238
rect 11348 4826 11376 6870
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11150 4584 11206 4593
rect 11060 4548 11112 4554
rect 11150 4519 11206 4528
rect 11060 4490 11112 4496
rect 11072 3738 11100 4490
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 11440 3670 11468 6734
rect 11428 3664 11480 3670
rect 11428 3606 11480 3612
rect 11532 3398 11560 8910
rect 11716 6866 11744 12582
rect 11808 8294 11836 17478
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11900 12170 11928 16934
rect 12084 16810 12112 18226
rect 12348 17196 12400 17202
rect 12348 17138 12400 17144
rect 11992 16782 12112 16810
rect 12360 16794 12388 17138
rect 12348 16788 12400 16794
rect 11888 12164 11940 12170
rect 11888 12106 11940 12112
rect 11888 11824 11940 11830
rect 11888 11766 11940 11772
rect 11900 9042 11928 11766
rect 11992 9382 12020 16782
rect 12348 16730 12400 16736
rect 12256 16584 12308 16590
rect 12256 16526 12308 16532
rect 12164 15564 12216 15570
rect 12164 15506 12216 15512
rect 12176 15026 12204 15506
rect 12164 15020 12216 15026
rect 12164 14962 12216 14968
rect 12268 14346 12296 16526
rect 12452 15978 12480 20878
rect 12636 17746 12664 24686
rect 12808 24608 12860 24614
rect 12808 24550 12860 24556
rect 12820 23866 12848 24550
rect 12808 23860 12860 23866
rect 12808 23802 12860 23808
rect 12716 18692 12768 18698
rect 12716 18634 12768 18640
rect 12728 18204 12756 18634
rect 12820 18358 12848 23802
rect 12912 22094 12940 24754
rect 13096 22098 13124 26318
rect 13360 25764 13412 25770
rect 13360 25706 13412 25712
rect 13372 25226 13400 25706
rect 13360 25220 13412 25226
rect 13360 25162 13412 25168
rect 13464 24818 13492 28698
rect 14740 28688 14792 28694
rect 14740 28630 14792 28636
rect 14004 28620 14056 28626
rect 14004 28562 14056 28568
rect 14016 28082 14044 28562
rect 14464 28416 14516 28422
rect 14464 28358 14516 28364
rect 14476 28150 14504 28358
rect 14464 28144 14516 28150
rect 14464 28086 14516 28092
rect 14004 28076 14056 28082
rect 14004 28018 14056 28024
rect 13544 27056 13596 27062
rect 13544 26998 13596 27004
rect 13556 26586 13584 26998
rect 13544 26580 13596 26586
rect 13544 26522 13596 26528
rect 13636 25900 13688 25906
rect 13636 25842 13688 25848
rect 13648 24954 13676 25842
rect 13636 24948 13688 24954
rect 13636 24890 13688 24896
rect 13452 24812 13504 24818
rect 13452 24754 13504 24760
rect 13360 24744 13412 24750
rect 13360 24686 13412 24692
rect 13372 23866 13400 24686
rect 13636 24200 13688 24206
rect 13636 24142 13688 24148
rect 13360 23860 13412 23866
rect 13360 23802 13412 23808
rect 13648 23730 13676 24142
rect 13636 23724 13688 23730
rect 13636 23666 13688 23672
rect 13268 22432 13320 22438
rect 13268 22374 13320 22380
rect 12912 22066 13032 22094
rect 13004 20942 13032 22066
rect 13084 22092 13136 22098
rect 13084 22034 13136 22040
rect 13280 22030 13308 22374
rect 13268 22024 13320 22030
rect 13268 21966 13320 21972
rect 13084 21888 13136 21894
rect 13084 21830 13136 21836
rect 12992 20936 13044 20942
rect 12992 20878 13044 20884
rect 13096 20466 13124 21830
rect 13452 21480 13504 21486
rect 13452 21422 13504 21428
rect 13084 20460 13136 20466
rect 13084 20402 13136 20408
rect 13464 20058 13492 21422
rect 13452 20052 13504 20058
rect 13452 19994 13504 20000
rect 12900 19508 12952 19514
rect 12900 19450 12952 19456
rect 12912 18358 12940 19450
rect 13636 19440 13688 19446
rect 13636 19382 13688 19388
rect 12808 18352 12860 18358
rect 12808 18294 12860 18300
rect 12900 18352 12952 18358
rect 12900 18294 12952 18300
rect 12808 18216 12860 18222
rect 12728 18176 12808 18204
rect 12808 18158 12860 18164
rect 12624 17740 12676 17746
rect 12624 17682 12676 17688
rect 12532 17604 12584 17610
rect 12532 17546 12584 17552
rect 12440 15972 12492 15978
rect 12440 15914 12492 15920
rect 12440 14952 12492 14958
rect 12438 14920 12440 14929
rect 12492 14920 12494 14929
rect 12438 14855 12494 14864
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12256 14340 12308 14346
rect 12256 14282 12308 14288
rect 12072 13388 12124 13394
rect 12072 13330 12124 13336
rect 12084 12850 12112 13330
rect 12164 12980 12216 12986
rect 12164 12922 12216 12928
rect 12072 12844 12124 12850
rect 12072 12786 12124 12792
rect 12176 10266 12204 12922
rect 12256 12300 12308 12306
rect 12256 12242 12308 12248
rect 12268 11014 12296 12242
rect 12256 11008 12308 11014
rect 12256 10950 12308 10956
rect 12164 10260 12216 10266
rect 12164 10202 12216 10208
rect 12256 9444 12308 9450
rect 12256 9386 12308 9392
rect 11980 9376 12032 9382
rect 12032 9324 12204 9330
rect 11980 9318 12204 9324
rect 11992 9302 12204 9318
rect 11992 9253 12020 9302
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 11992 8566 12020 8774
rect 11980 8560 12032 8566
rect 11980 8502 12032 8508
rect 11796 8288 11848 8294
rect 11796 8230 11848 8236
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 11612 5636 11664 5642
rect 11612 5578 11664 5584
rect 11980 5636 12032 5642
rect 11980 5578 12032 5584
rect 11624 4078 11652 5578
rect 11992 4826 12020 5578
rect 11980 4820 12032 4826
rect 11980 4762 12032 4768
rect 11612 4072 11664 4078
rect 11612 4014 11664 4020
rect 11520 3392 11572 3398
rect 11520 3334 11572 3340
rect 11532 3126 11560 3334
rect 12084 3126 12112 7142
rect 12176 5914 12204 9302
rect 12268 9042 12296 9386
rect 12256 9036 12308 9042
rect 12256 8978 12308 8984
rect 12452 8974 12480 14554
rect 12544 9994 12572 17546
rect 12624 17264 12676 17270
rect 12624 17206 12676 17212
rect 12636 16794 12664 17206
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 12624 16176 12676 16182
rect 12624 16118 12676 16124
rect 12636 14618 12664 16118
rect 12624 14612 12676 14618
rect 12624 14554 12676 14560
rect 12716 13456 12768 13462
rect 12716 13398 12768 13404
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 12636 12918 12664 13262
rect 12728 13190 12756 13398
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12624 12912 12676 12918
rect 12624 12854 12676 12860
rect 12624 12640 12676 12646
rect 12622 12608 12624 12617
rect 12676 12608 12678 12617
rect 12622 12543 12678 12552
rect 12624 11892 12676 11898
rect 12624 11834 12676 11840
rect 12636 10674 12664 11834
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12532 9988 12584 9994
rect 12532 9930 12584 9936
rect 12440 8968 12492 8974
rect 12440 8910 12492 8916
rect 12820 6254 12848 18158
rect 13648 17882 13676 19382
rect 13636 17876 13688 17882
rect 13636 17818 13688 17824
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 13004 16726 13032 17138
rect 12992 16720 13044 16726
rect 12992 16662 13044 16668
rect 13832 15178 13860 17614
rect 13360 15156 13412 15162
rect 13360 15098 13412 15104
rect 13648 15150 13860 15178
rect 13372 14414 13400 15098
rect 13452 14612 13504 14618
rect 13452 14554 13504 14560
rect 13360 14408 13412 14414
rect 13360 14350 13412 14356
rect 13464 13870 13492 14554
rect 13176 13864 13228 13870
rect 13176 13806 13228 13812
rect 13452 13864 13504 13870
rect 13452 13806 13504 13812
rect 12900 13184 12952 13190
rect 12900 13126 12952 13132
rect 12912 12986 12940 13126
rect 12900 12980 12952 12986
rect 12900 12922 12952 12928
rect 13188 10742 13216 13806
rect 13544 13796 13596 13802
rect 13544 13738 13596 13744
rect 13556 13530 13584 13738
rect 13648 13734 13676 15150
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13728 14476 13780 14482
rect 13728 14418 13780 14424
rect 13740 14006 13768 14418
rect 13728 14000 13780 14006
rect 13728 13942 13780 13948
rect 13636 13728 13688 13734
rect 13636 13670 13688 13676
rect 13544 13524 13596 13530
rect 13544 13466 13596 13472
rect 13740 13394 13768 13942
rect 13832 13530 13860 14758
rect 14016 13734 14044 28018
rect 14752 26994 14780 28630
rect 15120 27946 15148 29158
rect 15292 28484 15344 28490
rect 15292 28426 15344 28432
rect 15200 28416 15252 28422
rect 15200 28358 15252 28364
rect 15212 28014 15240 28358
rect 15304 28014 15332 28426
rect 15200 28008 15252 28014
rect 15200 27950 15252 27956
rect 15292 28008 15344 28014
rect 15292 27950 15344 27956
rect 15108 27940 15160 27946
rect 15108 27882 15160 27888
rect 14740 26988 14792 26994
rect 14740 26930 14792 26936
rect 14372 26376 14424 26382
rect 14372 26318 14424 26324
rect 14648 26376 14700 26382
rect 14648 26318 14700 26324
rect 14384 26042 14412 26318
rect 14372 26036 14424 26042
rect 14372 25978 14424 25984
rect 14280 25900 14332 25906
rect 14280 25842 14332 25848
rect 14188 22704 14240 22710
rect 14188 22646 14240 22652
rect 14096 19984 14148 19990
rect 14096 19926 14148 19932
rect 14108 19310 14136 19926
rect 14096 19304 14148 19310
rect 14096 19246 14148 19252
rect 14200 19174 14228 22646
rect 14188 19168 14240 19174
rect 14188 19110 14240 19116
rect 14188 18964 14240 18970
rect 14188 18906 14240 18912
rect 14200 18698 14228 18906
rect 14188 18692 14240 18698
rect 14188 18634 14240 18640
rect 14188 18352 14240 18358
rect 14188 18294 14240 18300
rect 14200 17882 14228 18294
rect 14188 17876 14240 17882
rect 14188 17818 14240 17824
rect 14292 14958 14320 25842
rect 14556 24676 14608 24682
rect 14556 24618 14608 24624
rect 14372 23792 14424 23798
rect 14372 23734 14424 23740
rect 14384 23186 14412 23734
rect 14464 23520 14516 23526
rect 14464 23462 14516 23468
rect 14372 23180 14424 23186
rect 14372 23122 14424 23128
rect 14476 23050 14504 23462
rect 14464 23044 14516 23050
rect 14464 22986 14516 22992
rect 14568 22094 14596 24618
rect 14476 22066 14596 22094
rect 14660 22094 14688 26318
rect 14752 24834 14780 26930
rect 14924 26920 14976 26926
rect 14924 26862 14976 26868
rect 14936 26586 14964 26862
rect 14924 26580 14976 26586
rect 14924 26522 14976 26528
rect 14924 24880 14976 24886
rect 14752 24806 14872 24834
rect 14924 24822 14976 24828
rect 14844 24750 14872 24806
rect 14832 24744 14884 24750
rect 14832 24686 14884 24692
rect 14936 24410 14964 24822
rect 14924 24404 14976 24410
rect 14924 24346 14976 24352
rect 15016 23724 15068 23730
rect 15016 23666 15068 23672
rect 14924 23316 14976 23322
rect 14924 23258 14976 23264
rect 14660 22066 14780 22094
rect 14372 20256 14424 20262
rect 14372 20198 14424 20204
rect 14384 18222 14412 20198
rect 14372 18216 14424 18222
rect 14372 18158 14424 18164
rect 14372 16720 14424 16726
rect 14372 16662 14424 16668
rect 14280 14952 14332 14958
rect 14280 14894 14332 14900
rect 14004 13728 14056 13734
rect 14004 13670 14056 13676
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13728 13388 13780 13394
rect 13728 13330 13780 13336
rect 13740 11898 13768 13330
rect 14188 13320 14240 13326
rect 14188 13262 14240 13268
rect 14200 12714 14228 13262
rect 14292 12918 14320 14894
rect 14280 12912 14332 12918
rect 14280 12854 14332 12860
rect 14188 12708 14240 12714
rect 14188 12650 14240 12656
rect 14292 12322 14320 12854
rect 14384 12434 14412 16662
rect 14476 15570 14504 22066
rect 14556 20936 14608 20942
rect 14556 20878 14608 20884
rect 14568 17202 14596 20878
rect 14648 20800 14700 20806
rect 14648 20742 14700 20748
rect 14660 20466 14688 20742
rect 14648 20460 14700 20466
rect 14648 20402 14700 20408
rect 14648 18760 14700 18766
rect 14648 18702 14700 18708
rect 14660 17542 14688 18702
rect 14648 17536 14700 17542
rect 14648 17478 14700 17484
rect 14556 17196 14608 17202
rect 14556 17138 14608 17144
rect 14660 16726 14688 17478
rect 14648 16720 14700 16726
rect 14648 16662 14700 16668
rect 14554 16552 14610 16561
rect 14554 16487 14556 16496
rect 14608 16487 14610 16496
rect 14556 16458 14608 16464
rect 14464 15564 14516 15570
rect 14516 15524 14688 15552
rect 14464 15506 14516 15512
rect 14464 15020 14516 15026
rect 14464 14962 14516 14968
rect 14476 14482 14504 14962
rect 14660 14906 14688 15524
rect 14752 15042 14780 22066
rect 14936 20942 14964 23258
rect 15028 22778 15056 23666
rect 15016 22772 15068 22778
rect 15016 22714 15068 22720
rect 15120 21554 15148 27882
rect 15384 26784 15436 26790
rect 15384 26726 15436 26732
rect 15396 26518 15424 26726
rect 15384 26512 15436 26518
rect 15384 26454 15436 26460
rect 15476 25968 15528 25974
rect 15476 25910 15528 25916
rect 15200 25832 15252 25838
rect 15200 25774 15252 25780
rect 15212 25498 15240 25774
rect 15488 25498 15516 25910
rect 15200 25492 15252 25498
rect 15200 25434 15252 25440
rect 15476 25492 15528 25498
rect 15476 25434 15528 25440
rect 15476 24744 15528 24750
rect 15476 24686 15528 24692
rect 15108 21548 15160 21554
rect 15108 21490 15160 21496
rect 15108 21412 15160 21418
rect 15108 21354 15160 21360
rect 14924 20936 14976 20942
rect 14924 20878 14976 20884
rect 15120 20874 15148 21354
rect 15108 20868 15160 20874
rect 15108 20810 15160 20816
rect 15200 20868 15252 20874
rect 15200 20810 15252 20816
rect 15212 20058 15240 20810
rect 15384 20256 15436 20262
rect 15384 20198 15436 20204
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 15016 19916 15068 19922
rect 15016 19858 15068 19864
rect 14832 19168 14884 19174
rect 14832 19110 14884 19116
rect 14844 18766 14872 19110
rect 14832 18760 14884 18766
rect 14832 18702 14884 18708
rect 14832 18216 14884 18222
rect 14832 18158 14884 18164
rect 14844 17270 14872 18158
rect 15028 17678 15056 19858
rect 15108 19848 15160 19854
rect 15108 19790 15160 19796
rect 15120 18970 15148 19790
rect 15200 19372 15252 19378
rect 15200 19314 15252 19320
rect 15108 18964 15160 18970
rect 15108 18906 15160 18912
rect 15016 17672 15068 17678
rect 15016 17614 15068 17620
rect 14832 17264 14884 17270
rect 14832 17206 14884 17212
rect 15108 16992 15160 16998
rect 15108 16934 15160 16940
rect 15120 15366 15148 16934
rect 15016 15360 15068 15366
rect 15014 15328 15016 15337
rect 15108 15360 15160 15366
rect 15068 15328 15070 15337
rect 15108 15302 15160 15308
rect 15014 15263 15070 15272
rect 14752 15014 15148 15042
rect 14660 14878 14780 14906
rect 14464 14476 14516 14482
rect 14464 14418 14516 14424
rect 14556 13524 14608 13530
rect 14556 13466 14608 13472
rect 14384 12406 14504 12434
rect 14292 12294 14412 12322
rect 14384 12238 14412 12294
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 13728 11892 13780 11898
rect 13728 11834 13780 11840
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13176 10736 13228 10742
rect 13176 10678 13228 10684
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 13648 9994 13676 10406
rect 13636 9988 13688 9994
rect 13636 9930 13688 9936
rect 13740 8022 13768 11494
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 14016 10266 14044 10610
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 14004 10260 14056 10266
rect 14004 10202 14056 10208
rect 14384 10130 14412 10406
rect 14372 10124 14424 10130
rect 14372 10066 14424 10072
rect 13912 9444 13964 9450
rect 13912 9386 13964 9392
rect 13924 8362 13952 9386
rect 14280 9376 14332 9382
rect 14280 9318 14332 9324
rect 13912 8356 13964 8362
rect 13912 8298 13964 8304
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 14004 8288 14056 8294
rect 14004 8230 14056 8236
rect 13728 8016 13780 8022
rect 13728 7958 13780 7964
rect 13832 7750 13860 8230
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 14016 7546 14044 8230
rect 14292 7886 14320 9318
rect 14476 9110 14504 12406
rect 14568 12170 14596 13466
rect 14556 12164 14608 12170
rect 14556 12106 14608 12112
rect 14752 11830 14780 14878
rect 15016 13728 15068 13734
rect 15016 13670 15068 13676
rect 14740 11824 14792 11830
rect 14740 11766 14792 11772
rect 14924 11008 14976 11014
rect 14924 10950 14976 10956
rect 14556 10124 14608 10130
rect 14556 10066 14608 10072
rect 14464 9104 14516 9110
rect 14464 9046 14516 9052
rect 14464 8356 14516 8362
rect 14464 8298 14516 8304
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14004 7540 14056 7546
rect 14004 7482 14056 7488
rect 13912 7472 13964 7478
rect 13912 7414 13964 7420
rect 13820 7268 13872 7274
rect 13820 7210 13872 7216
rect 13832 6934 13860 7210
rect 13924 6934 13952 7414
rect 14292 7342 14320 7822
rect 14280 7336 14332 7342
rect 14280 7278 14332 7284
rect 13820 6928 13872 6934
rect 13820 6870 13872 6876
rect 13912 6928 13964 6934
rect 13912 6870 13964 6876
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 12164 5908 12216 5914
rect 12164 5850 12216 5856
rect 14292 5642 14320 7278
rect 14476 6905 14504 8298
rect 14568 7478 14596 10066
rect 14936 9994 14964 10950
rect 15028 10810 15056 13670
rect 15120 11014 15148 15014
rect 15212 12434 15240 19314
rect 15396 19310 15424 20198
rect 15384 19304 15436 19310
rect 15384 19246 15436 19252
rect 15384 12640 15436 12646
rect 15384 12582 15436 12588
rect 15212 12406 15332 12434
rect 15108 11008 15160 11014
rect 15108 10950 15160 10956
rect 15016 10804 15068 10810
rect 15016 10746 15068 10752
rect 14924 9988 14976 9994
rect 14924 9930 14976 9936
rect 14556 7472 14608 7478
rect 14556 7414 14608 7420
rect 15120 7342 15148 10950
rect 15200 10192 15252 10198
rect 15200 10134 15252 10140
rect 15212 7818 15240 10134
rect 15200 7812 15252 7818
rect 15200 7754 15252 7760
rect 15108 7336 15160 7342
rect 15108 7278 15160 7284
rect 14648 6928 14700 6934
rect 14462 6896 14518 6905
rect 14648 6870 14700 6876
rect 14462 6831 14518 6840
rect 13636 5636 13688 5642
rect 13636 5578 13688 5584
rect 14280 5636 14332 5642
rect 14280 5578 14332 5584
rect 13648 5273 13676 5578
rect 13924 5370 14044 5386
rect 13924 5364 14056 5370
rect 13924 5358 14004 5364
rect 13634 5264 13690 5273
rect 13634 5199 13690 5208
rect 13924 5030 13952 5358
rect 14004 5306 14056 5312
rect 14188 5296 14240 5302
rect 14292 5284 14320 5578
rect 14240 5256 14320 5284
rect 14188 5238 14240 5244
rect 13912 5024 13964 5030
rect 13912 4966 13964 4972
rect 12256 4820 12308 4826
rect 12256 4762 12308 4768
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 14004 4820 14056 4826
rect 14004 4762 14056 4768
rect 12268 4486 12296 4762
rect 12360 4554 12388 4762
rect 12348 4548 12400 4554
rect 12348 4490 12400 4496
rect 12256 4480 12308 4486
rect 12256 4422 12308 4428
rect 14016 4282 14044 4762
rect 14292 4622 14320 5256
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 13912 4276 13964 4282
rect 13912 4218 13964 4224
rect 14004 4276 14056 4282
rect 14004 4218 14056 4224
rect 13924 4185 13952 4218
rect 13910 4176 13966 4185
rect 13910 4111 13966 4120
rect 12992 4072 13044 4078
rect 12992 4014 13044 4020
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 13004 3670 13032 4014
rect 12992 3664 13044 3670
rect 12992 3606 13044 3612
rect 13464 3194 13492 4014
rect 14292 3942 14320 4558
rect 14476 4554 14504 6831
rect 14464 4548 14516 4554
rect 14464 4490 14516 4496
rect 14660 3942 14688 6870
rect 15304 6254 15332 12406
rect 15396 7324 15424 12582
rect 15488 8634 15516 24686
rect 15580 15162 15608 29582
rect 15844 29504 15896 29510
rect 15844 29446 15896 29452
rect 16580 29504 16632 29510
rect 16580 29446 16632 29452
rect 15856 29170 15884 29446
rect 15844 29164 15896 29170
rect 15844 29106 15896 29112
rect 16120 28144 16172 28150
rect 16120 28086 16172 28092
rect 16132 25498 16160 28086
rect 16488 26920 16540 26926
rect 16488 26862 16540 26868
rect 16500 26450 16528 26862
rect 16488 26444 16540 26450
rect 16488 26386 16540 26392
rect 16592 25906 16620 29446
rect 16764 27464 16816 27470
rect 16764 27406 16816 27412
rect 16776 27062 16804 27406
rect 17500 27396 17552 27402
rect 17500 27338 17552 27344
rect 17512 27130 17540 27338
rect 17500 27124 17552 27130
rect 17500 27066 17552 27072
rect 16764 27056 16816 27062
rect 16764 26998 16816 27004
rect 16672 26784 16724 26790
rect 16672 26726 16724 26732
rect 16684 26450 16712 26726
rect 16672 26444 16724 26450
rect 16672 26386 16724 26392
rect 16580 25900 16632 25906
rect 16580 25842 16632 25848
rect 16212 25832 16264 25838
rect 16212 25774 16264 25780
rect 16120 25492 16172 25498
rect 16120 25434 16172 25440
rect 16224 23322 16252 25774
rect 16592 23594 16620 25842
rect 16776 25378 16804 26998
rect 17972 26994 18000 37062
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 18052 36916 18104 36922
rect 18052 36858 18104 36864
rect 18064 30938 18092 36858
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19432 31340 19484 31346
rect 19432 31282 19484 31288
rect 18052 30932 18104 30938
rect 18052 30874 18104 30880
rect 18880 30660 18932 30666
rect 18880 30602 18932 30608
rect 18892 29578 18920 30602
rect 19444 30394 19472 31282
rect 19524 31272 19576 31278
rect 19524 31214 19576 31220
rect 19536 30802 19564 31214
rect 19708 31136 19760 31142
rect 19708 31078 19760 31084
rect 19720 30802 19748 31078
rect 19524 30796 19576 30802
rect 19524 30738 19576 30744
rect 19708 30796 19760 30802
rect 19708 30738 19760 30744
rect 19984 30728 20036 30734
rect 19984 30670 20036 30676
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19432 30388 19484 30394
rect 19432 30330 19484 30336
rect 19248 30252 19300 30258
rect 19248 30194 19300 30200
rect 18144 29572 18196 29578
rect 18144 29514 18196 29520
rect 18236 29572 18288 29578
rect 18236 29514 18288 29520
rect 18880 29572 18932 29578
rect 18880 29514 18932 29520
rect 18156 29306 18184 29514
rect 18144 29300 18196 29306
rect 18144 29242 18196 29248
rect 18144 27396 18196 27402
rect 18144 27338 18196 27344
rect 17592 26988 17644 26994
rect 17592 26930 17644 26936
rect 17960 26988 18012 26994
rect 17960 26930 18012 26936
rect 17604 26586 17632 26930
rect 17592 26580 17644 26586
rect 17592 26522 17644 26528
rect 18156 26518 18184 27338
rect 18248 27130 18276 29514
rect 18236 27124 18288 27130
rect 18236 27066 18288 27072
rect 18696 26920 18748 26926
rect 18696 26862 18748 26868
rect 18144 26512 18196 26518
rect 18144 26454 18196 26460
rect 16684 25350 16804 25378
rect 16684 24274 16712 25350
rect 16764 25288 16816 25294
rect 16764 25230 16816 25236
rect 16856 25288 16908 25294
rect 16856 25230 16908 25236
rect 16672 24268 16724 24274
rect 16672 24210 16724 24216
rect 16684 24177 16712 24210
rect 16670 24168 16726 24177
rect 16670 24103 16726 24112
rect 16672 23656 16724 23662
rect 16672 23598 16724 23604
rect 16580 23588 16632 23594
rect 16580 23530 16632 23536
rect 16212 23316 16264 23322
rect 16212 23258 16264 23264
rect 16684 23254 16712 23598
rect 16776 23322 16804 25230
rect 16764 23316 16816 23322
rect 16764 23258 16816 23264
rect 16672 23248 16724 23254
rect 16672 23190 16724 23196
rect 16028 23112 16080 23118
rect 16028 23054 16080 23060
rect 15660 22636 15712 22642
rect 15660 22578 15712 22584
rect 15672 19718 15700 22578
rect 16040 22234 16068 23054
rect 16868 22642 16896 25230
rect 17868 25220 17920 25226
rect 17868 25162 17920 25168
rect 16948 24200 17000 24206
rect 16948 24142 17000 24148
rect 16120 22636 16172 22642
rect 16120 22578 16172 22584
rect 16856 22636 16908 22642
rect 16856 22578 16908 22584
rect 16028 22228 16080 22234
rect 16028 22170 16080 22176
rect 16132 22166 16160 22578
rect 16960 22506 16988 24142
rect 17040 23792 17092 23798
rect 17040 23734 17092 23740
rect 17052 22778 17080 23734
rect 17040 22772 17092 22778
rect 17040 22714 17092 22720
rect 17776 22636 17828 22642
rect 17776 22578 17828 22584
rect 16948 22500 17000 22506
rect 16948 22442 17000 22448
rect 17788 22166 17816 22578
rect 16120 22160 16172 22166
rect 16120 22102 16172 22108
rect 17776 22160 17828 22166
rect 17776 22102 17828 22108
rect 16764 22024 16816 22030
rect 16764 21966 16816 21972
rect 16948 22024 17000 22030
rect 16948 21966 17000 21972
rect 16212 21684 16264 21690
rect 16212 21626 16264 21632
rect 15936 21616 15988 21622
rect 15936 21558 15988 21564
rect 15844 20392 15896 20398
rect 15844 20334 15896 20340
rect 15660 19712 15712 19718
rect 15660 19654 15712 19660
rect 15672 16454 15700 19654
rect 15856 18970 15884 20334
rect 15948 20058 15976 21558
rect 15936 20052 15988 20058
rect 15936 19994 15988 20000
rect 15948 19854 15976 19994
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 15844 18964 15896 18970
rect 15844 18906 15896 18912
rect 15844 18148 15896 18154
rect 15844 18090 15896 18096
rect 15660 16448 15712 16454
rect 15660 16390 15712 16396
rect 15672 15434 15700 16390
rect 15660 15428 15712 15434
rect 15660 15370 15712 15376
rect 15568 15156 15620 15162
rect 15568 15098 15620 15104
rect 15752 14408 15804 14414
rect 15752 14350 15804 14356
rect 15764 13938 15792 14350
rect 15752 13932 15804 13938
rect 15752 13874 15804 13880
rect 15660 13524 15712 13530
rect 15660 13466 15712 13472
rect 15568 13456 15620 13462
rect 15568 13398 15620 13404
rect 15580 12782 15608 13398
rect 15672 12850 15700 13466
rect 15660 12844 15712 12850
rect 15660 12786 15712 12792
rect 15568 12776 15620 12782
rect 15568 12718 15620 12724
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 15856 8566 15884 18090
rect 16028 16652 16080 16658
rect 16028 16594 16080 16600
rect 16040 15337 16068 16594
rect 16026 15328 16082 15337
rect 16026 15263 16082 15272
rect 16040 13190 16068 15263
rect 16224 14890 16252 21626
rect 16488 20392 16540 20398
rect 16488 20334 16540 20340
rect 16500 19446 16528 20334
rect 16580 19984 16632 19990
rect 16580 19926 16632 19932
rect 16488 19440 16540 19446
rect 16488 19382 16540 19388
rect 16396 18964 16448 18970
rect 16396 18906 16448 18912
rect 16408 18698 16436 18906
rect 16396 18692 16448 18698
rect 16396 18634 16448 18640
rect 16408 17746 16436 18634
rect 16592 17746 16620 19926
rect 16776 19922 16804 21966
rect 16960 21146 16988 21966
rect 17592 21548 17644 21554
rect 17592 21490 17644 21496
rect 16948 21140 17000 21146
rect 16948 21082 17000 21088
rect 17604 21078 17632 21490
rect 17592 21072 17644 21078
rect 17592 21014 17644 21020
rect 17408 20868 17460 20874
rect 17408 20810 17460 20816
rect 16764 19916 16816 19922
rect 16764 19858 16816 19864
rect 16948 19780 17000 19786
rect 16948 19722 17000 19728
rect 17224 19780 17276 19786
rect 17224 19722 17276 19728
rect 16856 18828 16908 18834
rect 16856 18770 16908 18776
rect 16868 18358 16896 18770
rect 16960 18698 16988 19722
rect 17236 19514 17264 19722
rect 17224 19508 17276 19514
rect 17224 19450 17276 19456
rect 17040 19372 17092 19378
rect 17040 19314 17092 19320
rect 17316 19372 17368 19378
rect 17316 19314 17368 19320
rect 17052 18834 17080 19314
rect 17040 18828 17092 18834
rect 17040 18770 17092 18776
rect 16948 18692 17000 18698
rect 16948 18634 17000 18640
rect 16856 18352 16908 18358
rect 16856 18294 16908 18300
rect 16396 17740 16448 17746
rect 16396 17682 16448 17688
rect 16580 17740 16632 17746
rect 16580 17682 16632 17688
rect 16672 17672 16724 17678
rect 16672 17614 16724 17620
rect 16684 17066 16712 17614
rect 17052 17338 17080 18770
rect 17328 18426 17356 19314
rect 17316 18420 17368 18426
rect 17420 18408 17448 20810
rect 17592 19780 17644 19786
rect 17592 19722 17644 19728
rect 17604 19514 17632 19722
rect 17592 19508 17644 19514
rect 17592 19450 17644 19456
rect 17420 18380 17540 18408
rect 17316 18362 17368 18368
rect 17408 18284 17460 18290
rect 17408 18226 17460 18232
rect 17132 18080 17184 18086
rect 17132 18022 17184 18028
rect 17144 17882 17172 18022
rect 17132 17876 17184 17882
rect 17132 17818 17184 17824
rect 17040 17332 17092 17338
rect 17040 17274 17092 17280
rect 16672 17060 16724 17066
rect 16672 17002 16724 17008
rect 17420 16454 17448 18226
rect 17408 16448 17460 16454
rect 17408 16390 17460 16396
rect 17132 15428 17184 15434
rect 17132 15370 17184 15376
rect 16488 15156 16540 15162
rect 16488 15098 16540 15104
rect 16212 14884 16264 14890
rect 16212 14826 16264 14832
rect 16028 13184 16080 13190
rect 16028 13126 16080 13132
rect 16224 12714 16252 14826
rect 16212 12708 16264 12714
rect 16212 12650 16264 12656
rect 16500 12646 16528 15098
rect 17144 14278 17172 15370
rect 17512 14414 17540 18380
rect 17604 16046 17632 19450
rect 17788 17218 17816 22102
rect 17880 22098 17908 25162
rect 17960 22432 18012 22438
rect 17960 22374 18012 22380
rect 17868 22092 17920 22098
rect 17868 22034 17920 22040
rect 17972 21622 18000 22374
rect 18156 22094 18184 26454
rect 18708 25294 18736 26862
rect 18420 25288 18472 25294
rect 18420 25230 18472 25236
rect 18696 25288 18748 25294
rect 18696 25230 18748 25236
rect 18328 24132 18380 24138
rect 18328 24074 18380 24080
rect 18340 23322 18368 24074
rect 18328 23316 18380 23322
rect 18328 23258 18380 23264
rect 18156 22066 18276 22094
rect 17960 21616 18012 21622
rect 17960 21558 18012 21564
rect 17868 21480 17920 21486
rect 17868 21422 17920 21428
rect 17880 21146 17908 21422
rect 17868 21140 17920 21146
rect 17868 21082 17920 21088
rect 17960 19440 18012 19446
rect 17960 19382 18012 19388
rect 17696 17190 17816 17218
rect 17868 17264 17920 17270
rect 17868 17206 17920 17212
rect 17592 16040 17644 16046
rect 17592 15982 17644 15988
rect 17590 15192 17646 15201
rect 17590 15127 17646 15136
rect 17604 15094 17632 15127
rect 17592 15088 17644 15094
rect 17592 15030 17644 15036
rect 17500 14408 17552 14414
rect 17500 14350 17552 14356
rect 17132 14272 17184 14278
rect 17132 14214 17184 14220
rect 17592 14272 17644 14278
rect 17592 14214 17644 14220
rect 17604 13802 17632 14214
rect 17592 13796 17644 13802
rect 17592 13738 17644 13744
rect 17500 13184 17552 13190
rect 17500 13126 17552 13132
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 16488 12640 16540 12646
rect 16488 12582 16540 12588
rect 17040 12436 17092 12442
rect 17040 12378 17092 12384
rect 17052 11762 17080 12378
rect 17224 12368 17276 12374
rect 17224 12310 17276 12316
rect 17236 12102 17264 12310
rect 17224 12096 17276 12102
rect 17224 12038 17276 12044
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 17328 11694 17356 12786
rect 17512 12434 17540 13126
rect 17420 12406 17540 12434
rect 17132 11688 17184 11694
rect 17132 11630 17184 11636
rect 17316 11688 17368 11694
rect 17316 11630 17368 11636
rect 17040 11552 17092 11558
rect 17040 11494 17092 11500
rect 17052 11218 17080 11494
rect 17040 11212 17092 11218
rect 17040 11154 17092 11160
rect 17144 11150 17172 11630
rect 16580 11144 16632 11150
rect 16580 11086 16632 11092
rect 17132 11144 17184 11150
rect 17132 11086 17184 11092
rect 16592 10606 16620 11086
rect 17316 11076 17368 11082
rect 17316 11018 17368 11024
rect 16580 10600 16632 10606
rect 16580 10542 16632 10548
rect 16592 8974 16620 10542
rect 17328 10198 17356 11018
rect 17420 10742 17448 12406
rect 17696 11506 17724 17190
rect 17880 17066 17908 17206
rect 17868 17060 17920 17066
rect 17868 17002 17920 17008
rect 17972 16590 18000 19382
rect 18248 19009 18276 22066
rect 18328 19916 18380 19922
rect 18328 19858 18380 19864
rect 18234 19000 18290 19009
rect 18234 18935 18290 18944
rect 17960 16584 18012 16590
rect 17960 16526 18012 16532
rect 18050 16552 18106 16561
rect 18050 16487 18052 16496
rect 18104 16487 18106 16496
rect 18052 16458 18104 16464
rect 17960 16448 18012 16454
rect 17960 16390 18012 16396
rect 17972 16114 18000 16390
rect 17960 16108 18012 16114
rect 17960 16050 18012 16056
rect 17868 16040 17920 16046
rect 17868 15982 17920 15988
rect 17880 15570 17908 15982
rect 17960 15972 18012 15978
rect 17960 15914 18012 15920
rect 17868 15564 17920 15570
rect 17868 15506 17920 15512
rect 17880 15026 17908 15506
rect 17868 15020 17920 15026
rect 17868 14962 17920 14968
rect 17880 14482 17908 14962
rect 17868 14476 17920 14482
rect 17868 14418 17920 14424
rect 17776 14272 17828 14278
rect 17776 14214 17828 14220
rect 17788 13938 17816 14214
rect 17880 13938 17908 14418
rect 17776 13932 17828 13938
rect 17776 13874 17828 13880
rect 17868 13932 17920 13938
rect 17868 13874 17920 13880
rect 17880 12986 17908 13874
rect 17972 13870 18000 15914
rect 18144 14816 18196 14822
rect 18144 14758 18196 14764
rect 18156 14618 18184 14758
rect 18144 14612 18196 14618
rect 18144 14554 18196 14560
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 17868 12980 17920 12986
rect 17868 12922 17920 12928
rect 17776 12640 17828 12646
rect 17776 12582 17828 12588
rect 17788 11830 17816 12582
rect 18156 11898 18184 14554
rect 18340 12434 18368 19858
rect 18432 16454 18460 25230
rect 18892 24274 18920 29514
rect 19260 29170 19288 30194
rect 19340 29640 19392 29646
rect 19340 29582 19392 29588
rect 19352 29306 19380 29582
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19996 29306 20024 30670
rect 20168 30592 20220 30598
rect 20168 30534 20220 30540
rect 20180 29782 20208 30534
rect 20168 29776 20220 29782
rect 20168 29718 20220 29724
rect 21088 29640 21140 29646
rect 21088 29582 21140 29588
rect 20996 29504 21048 29510
rect 20996 29446 21048 29452
rect 19340 29300 19392 29306
rect 19340 29242 19392 29248
rect 19984 29300 20036 29306
rect 19984 29242 20036 29248
rect 21008 29170 21036 29446
rect 19248 29164 19300 29170
rect 19248 29106 19300 29112
rect 20168 29164 20220 29170
rect 20168 29106 20220 29112
rect 20996 29164 21048 29170
rect 20996 29106 21048 29112
rect 19984 28416 20036 28422
rect 19984 28358 20036 28364
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19996 28218 20024 28358
rect 19984 28212 20036 28218
rect 19984 28154 20036 28160
rect 20076 28144 20128 28150
rect 20076 28086 20128 28092
rect 19432 27668 19484 27674
rect 19432 27610 19484 27616
rect 19340 26988 19392 26994
rect 19340 26930 19392 26936
rect 19352 26042 19380 26930
rect 19340 26036 19392 26042
rect 19340 25978 19392 25984
rect 19340 25900 19392 25906
rect 19340 25842 19392 25848
rect 18880 24268 18932 24274
rect 18880 24210 18932 24216
rect 19352 23186 19380 25842
rect 19444 23254 19472 27610
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 20088 26586 20116 28086
rect 20180 27946 20208 29106
rect 20904 28144 20956 28150
rect 20904 28086 20956 28092
rect 20168 27940 20220 27946
rect 20168 27882 20220 27888
rect 20628 27940 20680 27946
rect 20628 27882 20680 27888
rect 20076 26580 20128 26586
rect 20076 26522 20128 26528
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19984 25696 20036 25702
rect 19984 25638 20036 25644
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19616 24744 19668 24750
rect 19616 24686 19668 24692
rect 19628 24274 19656 24686
rect 19996 24274 20024 25638
rect 19616 24268 19668 24274
rect 19616 24210 19668 24216
rect 19984 24268 20036 24274
rect 19984 24210 20036 24216
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19996 23526 20024 24210
rect 19984 23520 20036 23526
rect 19984 23462 20036 23468
rect 19432 23248 19484 23254
rect 19432 23190 19484 23196
rect 19340 23180 19392 23186
rect 19340 23122 19392 23128
rect 19984 23112 20036 23118
rect 19984 23054 20036 23060
rect 18512 23044 18564 23050
rect 18512 22986 18564 22992
rect 19340 23044 19392 23050
rect 19340 22986 19392 22992
rect 18524 22778 18552 22986
rect 18512 22772 18564 22778
rect 18512 22714 18564 22720
rect 18524 18834 18552 22714
rect 19156 22636 19208 22642
rect 19156 22578 19208 22584
rect 18880 19916 18932 19922
rect 18880 19858 18932 19864
rect 18788 19168 18840 19174
rect 18788 19110 18840 19116
rect 18512 18828 18564 18834
rect 18512 18770 18564 18776
rect 18696 18352 18748 18358
rect 18696 18294 18748 18300
rect 18604 18216 18656 18222
rect 18604 18158 18656 18164
rect 18616 17746 18644 18158
rect 18604 17740 18656 17746
rect 18604 17682 18656 17688
rect 18708 17338 18736 18294
rect 18696 17332 18748 17338
rect 18696 17274 18748 17280
rect 18696 17196 18748 17202
rect 18696 17138 18748 17144
rect 18708 16794 18736 17138
rect 18696 16788 18748 16794
rect 18696 16730 18748 16736
rect 18800 16674 18828 19110
rect 18616 16646 18828 16674
rect 18420 16448 18472 16454
rect 18420 16390 18472 16396
rect 18616 14929 18644 16646
rect 18696 16584 18748 16590
rect 18696 16526 18748 16532
rect 18708 16182 18736 16526
rect 18696 16176 18748 16182
rect 18748 16136 18828 16164
rect 18696 16118 18748 16124
rect 18800 16046 18828 16136
rect 18696 16040 18748 16046
rect 18696 15982 18748 15988
rect 18788 16040 18840 16046
rect 18788 15982 18840 15988
rect 18708 15858 18736 15982
rect 18892 15858 18920 19858
rect 18708 15830 18920 15858
rect 18696 15496 18748 15502
rect 18696 15438 18748 15444
rect 18708 15366 18736 15438
rect 18696 15360 18748 15366
rect 18696 15302 18748 15308
rect 18694 15192 18750 15201
rect 18694 15127 18696 15136
rect 18748 15127 18750 15136
rect 18696 15098 18748 15104
rect 18602 14920 18658 14929
rect 18602 14855 18658 14864
rect 18512 14816 18564 14822
rect 18512 14758 18564 14764
rect 18524 14006 18552 14758
rect 18512 14000 18564 14006
rect 18512 13942 18564 13948
rect 18340 12406 18460 12434
rect 18144 11892 18196 11898
rect 18144 11834 18196 11840
rect 17776 11824 17828 11830
rect 17776 11766 17828 11772
rect 17696 11478 17816 11506
rect 17788 11218 17816 11478
rect 17776 11212 17828 11218
rect 17776 11154 17828 11160
rect 17408 10736 17460 10742
rect 17408 10678 17460 10684
rect 17316 10192 17368 10198
rect 17316 10134 17368 10140
rect 18144 9580 18196 9586
rect 18144 9522 18196 9528
rect 17960 9512 18012 9518
rect 17960 9454 18012 9460
rect 16580 8968 16632 8974
rect 16580 8910 16632 8916
rect 16856 8900 16908 8906
rect 16856 8842 16908 8848
rect 16868 8634 16896 8842
rect 17868 8832 17920 8838
rect 17972 8820 18000 9454
rect 18156 9110 18184 9522
rect 18144 9104 18196 9110
rect 18144 9046 18196 9052
rect 18236 8968 18288 8974
rect 18236 8910 18288 8916
rect 17920 8792 18000 8820
rect 17868 8774 17920 8780
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 15844 8560 15896 8566
rect 15844 8502 15896 8508
rect 17972 8430 18000 8792
rect 18248 8566 18276 8910
rect 18236 8560 18288 8566
rect 18236 8502 18288 8508
rect 17868 8424 17920 8430
rect 17868 8366 17920 8372
rect 17960 8424 18012 8430
rect 17960 8366 18012 8372
rect 16120 8356 16172 8362
rect 16120 8298 16172 8304
rect 15568 7336 15620 7342
rect 15396 7296 15568 7324
rect 15568 7278 15620 7284
rect 15292 6248 15344 6254
rect 15292 6190 15344 6196
rect 14280 3936 14332 3942
rect 14280 3878 14332 3884
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 14188 3596 14240 3602
rect 14188 3538 14240 3544
rect 14200 3369 14228 3538
rect 14186 3360 14242 3369
rect 14186 3295 14242 3304
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 14292 3126 14320 3878
rect 14370 3632 14426 3641
rect 14370 3567 14426 3576
rect 14384 3534 14412 3567
rect 14372 3528 14424 3534
rect 14660 3505 14688 3878
rect 14752 3670 14780 3878
rect 14740 3664 14792 3670
rect 14740 3606 14792 3612
rect 15304 3602 15332 6190
rect 16028 5908 16080 5914
rect 16028 5850 16080 5856
rect 15752 5024 15804 5030
rect 15752 4966 15804 4972
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 15396 3602 15424 3674
rect 15292 3596 15344 3602
rect 15292 3538 15344 3544
rect 15384 3596 15436 3602
rect 15384 3538 15436 3544
rect 15016 3528 15068 3534
rect 14372 3470 14424 3476
rect 14646 3496 14702 3505
rect 14464 3460 14516 3466
rect 15016 3470 15068 3476
rect 14646 3431 14702 3440
rect 14464 3402 14516 3408
rect 14372 3392 14424 3398
rect 14372 3334 14424 3340
rect 14384 3126 14412 3334
rect 11520 3120 11572 3126
rect 11520 3062 11572 3068
rect 12072 3120 12124 3126
rect 12072 3062 12124 3068
rect 14280 3120 14332 3126
rect 14280 3062 14332 3068
rect 14372 3120 14424 3126
rect 14372 3062 14424 3068
rect 12084 2774 12112 3062
rect 14476 2990 14504 3402
rect 14464 2984 14516 2990
rect 14464 2926 14516 2932
rect 11992 2746 12112 2774
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 7760 1970 7788 2382
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 10324 2304 10376 2310
rect 10324 2246 10376 2252
rect 7748 1964 7800 1970
rect 7748 1906 7800 1912
rect 9048 800 9076 2246
rect 10336 800 10364 2246
rect 11624 800 11652 2382
rect 11704 2304 11756 2310
rect 11704 2246 11756 2252
rect 11716 2038 11744 2246
rect 11992 2106 12020 2746
rect 15028 2650 15056 3470
rect 15764 3398 15792 4966
rect 16040 4758 16068 5850
rect 16028 4752 16080 4758
rect 16028 4694 16080 4700
rect 15752 3392 15804 3398
rect 15752 3334 15804 3340
rect 15764 2922 15792 3334
rect 16132 2990 16160 8298
rect 17880 7857 17908 8366
rect 17972 7954 18000 8366
rect 17960 7948 18012 7954
rect 17960 7890 18012 7896
rect 17866 7848 17922 7857
rect 17866 7783 17922 7792
rect 17972 7342 18000 7890
rect 18052 7880 18104 7886
rect 18052 7822 18104 7828
rect 16304 7336 16356 7342
rect 16304 7278 16356 7284
rect 17960 7336 18012 7342
rect 17960 7278 18012 7284
rect 16316 7041 16344 7278
rect 16302 7032 16358 7041
rect 16302 6967 16358 6976
rect 16316 5574 16344 6967
rect 16580 6928 16632 6934
rect 16580 6870 16632 6876
rect 16592 6458 16620 6870
rect 17224 6860 17276 6866
rect 17224 6802 17276 6808
rect 17236 6662 17264 6802
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 16580 6452 16632 6458
rect 16580 6394 16632 6400
rect 16672 6452 16724 6458
rect 16672 6394 16724 6400
rect 16684 6186 16712 6394
rect 16672 6180 16724 6186
rect 16672 6122 16724 6128
rect 16304 5568 16356 5574
rect 16304 5510 16356 5516
rect 17224 5568 17276 5574
rect 17224 5510 17276 5516
rect 17132 5228 17184 5234
rect 17132 5170 17184 5176
rect 17040 5160 17092 5166
rect 17040 5102 17092 5108
rect 17052 4826 17080 5102
rect 17040 4820 17092 4826
rect 17040 4762 17092 4768
rect 16856 4752 16908 4758
rect 16856 4694 16908 4700
rect 16868 4282 16896 4694
rect 17040 4616 17092 4622
rect 17040 4558 17092 4564
rect 16856 4276 16908 4282
rect 16856 4218 16908 4224
rect 17052 3534 17080 4558
rect 17144 4282 17172 5170
rect 17236 5166 17264 5510
rect 17224 5160 17276 5166
rect 17224 5102 17276 5108
rect 17682 4584 17738 4593
rect 17682 4519 17738 4528
rect 17696 4486 17724 4519
rect 17224 4480 17276 4486
rect 17224 4422 17276 4428
rect 17592 4480 17644 4486
rect 17592 4422 17644 4428
rect 17684 4480 17736 4486
rect 17684 4422 17736 4428
rect 17236 4282 17264 4422
rect 17132 4276 17184 4282
rect 17132 4218 17184 4224
rect 17224 4276 17276 4282
rect 17224 4218 17276 4224
rect 17604 4214 17632 4422
rect 17592 4208 17644 4214
rect 17592 4150 17644 4156
rect 17684 4140 17736 4146
rect 17684 4082 17736 4088
rect 17696 4049 17724 4082
rect 17682 4040 17738 4049
rect 17682 3975 17738 3984
rect 17788 3942 17816 6598
rect 17972 5166 18000 7278
rect 17960 5160 18012 5166
rect 17960 5102 18012 5108
rect 17972 4214 18000 5102
rect 18064 4622 18092 7822
rect 18236 7812 18288 7818
rect 18236 7754 18288 7760
rect 18248 7342 18276 7754
rect 18328 7744 18380 7750
rect 18326 7712 18328 7721
rect 18380 7712 18382 7721
rect 18326 7647 18382 7656
rect 18328 7540 18380 7546
rect 18328 7482 18380 7488
rect 18340 7342 18368 7482
rect 18236 7336 18288 7342
rect 18236 7278 18288 7284
rect 18328 7336 18380 7342
rect 18328 7278 18380 7284
rect 18248 6798 18276 7278
rect 18236 6792 18288 6798
rect 18432 6769 18460 12406
rect 18616 9042 18644 14855
rect 19064 13728 19116 13734
rect 19064 13670 19116 13676
rect 18696 13320 18748 13326
rect 18696 13262 18748 13268
rect 18708 12714 18736 13262
rect 18696 12708 18748 12714
rect 18696 12650 18748 12656
rect 18972 11212 19024 11218
rect 18972 11154 19024 11160
rect 18604 9036 18656 9042
rect 18604 8978 18656 8984
rect 18984 8634 19012 11154
rect 18972 8628 19024 8634
rect 18972 8570 19024 8576
rect 18696 8084 18748 8090
rect 18696 8026 18748 8032
rect 18708 7886 18736 8026
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 18512 7744 18564 7750
rect 18512 7686 18564 7692
rect 18236 6734 18288 6740
rect 18418 6760 18474 6769
rect 18418 6695 18474 6704
rect 18432 5896 18460 6695
rect 18248 5868 18460 5896
rect 18142 5672 18198 5681
rect 18142 5607 18144 5616
rect 18196 5607 18198 5616
rect 18144 5578 18196 5584
rect 18248 4758 18276 5868
rect 18326 5400 18382 5409
rect 18326 5335 18382 5344
rect 18340 5166 18368 5335
rect 18524 5302 18552 7686
rect 19076 6798 19104 13670
rect 19168 12986 19196 22578
rect 19352 21962 19380 22986
rect 19432 22976 19484 22982
rect 19432 22918 19484 22924
rect 19340 21956 19392 21962
rect 19340 21898 19392 21904
rect 19444 20942 19472 22918
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19996 22778 20024 23054
rect 20076 22976 20128 22982
rect 20076 22918 20128 22924
rect 19984 22772 20036 22778
rect 19984 22714 20036 22720
rect 19984 21956 20036 21962
rect 19984 21898 20036 21904
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19800 21480 19852 21486
rect 19800 21422 19852 21428
rect 19812 21350 19840 21422
rect 19800 21344 19852 21350
rect 19800 21286 19852 21292
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19444 20602 19472 20878
rect 19812 20806 19840 21286
rect 19800 20800 19852 20806
rect 19800 20742 19852 20748
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19432 20596 19484 20602
rect 19432 20538 19484 20544
rect 19340 19848 19392 19854
rect 19340 19790 19392 19796
rect 19248 19304 19300 19310
rect 19248 19246 19300 19252
rect 19260 18698 19288 19246
rect 19248 18692 19300 18698
rect 19248 18634 19300 18640
rect 19248 17536 19300 17542
rect 19248 17478 19300 17484
rect 19260 17338 19288 17478
rect 19248 17332 19300 17338
rect 19248 17274 19300 17280
rect 19248 15904 19300 15910
rect 19248 15846 19300 15852
rect 19260 13274 19288 15846
rect 19352 15434 19380 19790
rect 19432 19712 19484 19718
rect 19432 19654 19484 19660
rect 19444 19378 19472 19654
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 19432 18624 19484 18630
rect 19432 18566 19484 18572
rect 19340 15428 19392 15434
rect 19340 15370 19392 15376
rect 19444 14958 19472 18566
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19996 18068 20024 21898
rect 20088 21622 20116 22918
rect 20076 21616 20128 21622
rect 20076 21558 20128 21564
rect 20076 20052 20128 20058
rect 20076 19994 20128 20000
rect 20088 18170 20116 19994
rect 20180 19990 20208 27882
rect 20352 26376 20404 26382
rect 20352 26318 20404 26324
rect 20364 26042 20392 26318
rect 20352 26036 20404 26042
rect 20352 25978 20404 25984
rect 20352 25900 20404 25906
rect 20352 25842 20404 25848
rect 20260 21888 20312 21894
rect 20260 21830 20312 21836
rect 20272 20942 20300 21830
rect 20364 21350 20392 25842
rect 20536 22024 20588 22030
rect 20536 21966 20588 21972
rect 20548 21468 20576 21966
rect 20640 21622 20668 27882
rect 20812 26852 20864 26858
rect 20812 26794 20864 26800
rect 20824 24274 20852 26794
rect 20916 24410 20944 28086
rect 20996 26784 21048 26790
rect 20996 26726 21048 26732
rect 21008 26314 21036 26726
rect 20996 26308 21048 26314
rect 20996 26250 21048 26256
rect 20904 24404 20956 24410
rect 20904 24346 20956 24352
rect 20812 24268 20864 24274
rect 20812 24210 20864 24216
rect 20720 24200 20772 24206
rect 20720 24142 20772 24148
rect 20732 22642 20760 24142
rect 20812 23180 20864 23186
rect 20812 23122 20864 23128
rect 20720 22636 20772 22642
rect 20720 22578 20772 22584
rect 20628 21616 20680 21622
rect 20628 21558 20680 21564
rect 20548 21440 20668 21468
rect 20352 21344 20404 21350
rect 20352 21286 20404 21292
rect 20536 21344 20588 21350
rect 20536 21286 20588 21292
rect 20260 20936 20312 20942
rect 20260 20878 20312 20884
rect 20260 20800 20312 20806
rect 20260 20742 20312 20748
rect 20352 20800 20404 20806
rect 20352 20742 20404 20748
rect 20168 19984 20220 19990
rect 20168 19926 20220 19932
rect 20168 19304 20220 19310
rect 20168 19246 20220 19252
rect 20180 18970 20208 19246
rect 20168 18964 20220 18970
rect 20168 18906 20220 18912
rect 20180 18290 20208 18906
rect 20168 18284 20220 18290
rect 20168 18226 20220 18232
rect 20088 18142 20208 18170
rect 19996 18040 20116 18068
rect 19984 17604 20036 17610
rect 19984 17546 20036 17552
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19800 16108 19852 16114
rect 19800 16050 19852 16056
rect 19812 15348 19840 16050
rect 19996 15706 20024 17546
rect 20088 16130 20116 18040
rect 20180 16250 20208 18142
rect 20168 16244 20220 16250
rect 20168 16186 20220 16192
rect 20088 16102 20208 16130
rect 19984 15700 20036 15706
rect 19984 15642 20036 15648
rect 19812 15320 20024 15348
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19432 14952 19484 14958
rect 19432 14894 19484 14900
rect 19524 14884 19576 14890
rect 19524 14826 19576 14832
rect 19536 14618 19564 14826
rect 19996 14618 20024 15320
rect 20180 14958 20208 16102
rect 20168 14952 20220 14958
rect 20168 14894 20220 14900
rect 19524 14612 19576 14618
rect 19524 14554 19576 14560
rect 19984 14612 20036 14618
rect 19984 14554 20036 14560
rect 20180 14278 20208 14894
rect 20168 14272 20220 14278
rect 20168 14214 20220 14220
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19260 13246 19380 13274
rect 19352 13190 19380 13246
rect 19248 13184 19300 13190
rect 19248 13126 19300 13132
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 19260 12986 19288 13126
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19156 12980 19208 12986
rect 19156 12922 19208 12928
rect 19248 12980 19300 12986
rect 19248 12922 19300 12928
rect 19168 10606 19196 12922
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19984 11212 20036 11218
rect 19984 11154 20036 11160
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19156 10600 19208 10606
rect 19156 10542 19208 10548
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19996 9654 20024 11154
rect 20168 11076 20220 11082
rect 20168 11018 20220 11024
rect 20076 9988 20128 9994
rect 20076 9930 20128 9936
rect 19984 9648 20036 9654
rect 19984 9590 20036 9596
rect 19156 9512 19208 9518
rect 19154 9480 19156 9489
rect 19248 9512 19300 9518
rect 19208 9480 19210 9489
rect 19248 9454 19300 9460
rect 19430 9480 19486 9489
rect 19154 9415 19210 9424
rect 19064 6792 19116 6798
rect 19064 6734 19116 6740
rect 18604 6112 18656 6118
rect 18604 6054 18656 6060
rect 18696 6112 18748 6118
rect 18696 6054 18748 6060
rect 18616 5846 18644 6054
rect 18604 5840 18656 5846
rect 18604 5782 18656 5788
rect 18512 5296 18564 5302
rect 18512 5238 18564 5244
rect 18602 5264 18658 5273
rect 18602 5199 18658 5208
rect 18616 5166 18644 5199
rect 18328 5160 18380 5166
rect 18328 5102 18380 5108
rect 18604 5160 18656 5166
rect 18604 5102 18656 5108
rect 18144 4752 18196 4758
rect 18144 4694 18196 4700
rect 18236 4752 18288 4758
rect 18236 4694 18288 4700
rect 18420 4752 18472 4758
rect 18420 4694 18472 4700
rect 18052 4616 18104 4622
rect 18052 4558 18104 4564
rect 18156 4570 18184 4694
rect 18432 4570 18460 4694
rect 18156 4542 18460 4570
rect 17960 4208 18012 4214
rect 17960 4150 18012 4156
rect 18328 4208 18380 4214
rect 18328 4150 18380 4156
rect 18512 4208 18564 4214
rect 18512 4150 18564 4156
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 17316 3664 17368 3670
rect 17314 3632 17316 3641
rect 17368 3632 17370 3641
rect 17314 3567 17370 3576
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 18052 3528 18104 3534
rect 18052 3470 18104 3476
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 17236 3194 17264 3334
rect 17224 3188 17276 3194
rect 17224 3130 17276 3136
rect 17868 3120 17920 3126
rect 17868 3062 17920 3068
rect 16120 2984 16172 2990
rect 16120 2926 16172 2932
rect 15752 2916 15804 2922
rect 15752 2858 15804 2864
rect 17880 2802 17908 3062
rect 18064 3058 18092 3470
rect 18144 3392 18196 3398
rect 18144 3334 18196 3340
rect 18052 3052 18104 3058
rect 18052 2994 18104 3000
rect 17880 2774 18092 2802
rect 18064 2650 18092 2774
rect 15016 2644 15068 2650
rect 15016 2586 15068 2592
rect 17960 2644 18012 2650
rect 17960 2586 18012 2592
rect 18052 2644 18104 2650
rect 18052 2586 18104 2592
rect 16672 2576 16724 2582
rect 16672 2518 16724 2524
rect 13544 2440 13596 2446
rect 13544 2382 13596 2388
rect 14832 2440 14884 2446
rect 14832 2382 14884 2388
rect 11980 2100 12032 2106
rect 11980 2042 12032 2048
rect 11704 2032 11756 2038
rect 11704 1974 11756 1980
rect 13556 800 13584 2382
rect 14844 800 14872 2382
rect 16684 2310 16712 2518
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 16672 2304 16724 2310
rect 16672 2246 16724 2252
rect 16776 800 16804 2382
rect 17972 2106 18000 2586
rect 18156 2446 18184 3334
rect 18340 3058 18368 4150
rect 18524 3738 18552 4150
rect 18512 3732 18564 3738
rect 18512 3674 18564 3680
rect 18604 3732 18656 3738
rect 18604 3674 18656 3680
rect 18328 3052 18380 3058
rect 18328 2994 18380 3000
rect 18616 2922 18644 3674
rect 18708 3534 18736 6054
rect 19076 4078 19104 6734
rect 19260 6322 19288 9454
rect 19430 9415 19486 9424
rect 19340 8968 19392 8974
rect 19340 8910 19392 8916
rect 19352 8090 19380 8910
rect 19340 8084 19392 8090
rect 19340 8026 19392 8032
rect 19340 7812 19392 7818
rect 19340 7754 19392 7760
rect 19352 6458 19380 7754
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19248 6316 19300 6322
rect 19248 6258 19300 6264
rect 19444 5114 19472 9415
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19708 8628 19760 8634
rect 19708 8570 19760 8576
rect 19616 8560 19668 8566
rect 19720 8537 19748 8570
rect 19996 8548 20024 9590
rect 20088 9586 20116 9930
rect 20180 9654 20208 11018
rect 20168 9648 20220 9654
rect 20168 9590 20220 9596
rect 20076 9580 20128 9586
rect 20076 9522 20128 9528
rect 20168 8968 20220 8974
rect 20168 8910 20220 8916
rect 20076 8832 20128 8838
rect 20076 8774 20128 8780
rect 19616 8502 19668 8508
rect 19706 8528 19762 8537
rect 19628 8401 19656 8502
rect 19904 8520 20024 8548
rect 19706 8463 19762 8472
rect 19800 8492 19852 8498
rect 19800 8434 19852 8440
rect 19614 8392 19670 8401
rect 19614 8327 19670 8336
rect 19812 8294 19840 8434
rect 19800 8288 19852 8294
rect 19628 8248 19800 8276
rect 19628 7818 19656 8248
rect 19800 8230 19852 8236
rect 19616 7812 19668 7818
rect 19616 7754 19668 7760
rect 19800 7812 19852 7818
rect 19904 7800 19932 8520
rect 19982 8392 20038 8401
rect 19982 8327 20038 8336
rect 19852 7772 19932 7800
rect 19800 7754 19852 7760
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19892 7336 19944 7342
rect 19892 7278 19944 7284
rect 19904 7002 19932 7278
rect 19892 6996 19944 7002
rect 19892 6938 19944 6944
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19996 6458 20024 8327
rect 20088 8090 20116 8774
rect 20180 8362 20208 8910
rect 20168 8356 20220 8362
rect 20168 8298 20220 8304
rect 20076 8084 20128 8090
rect 20076 8026 20128 8032
rect 20074 7848 20130 7857
rect 20074 7783 20130 7792
rect 19984 6452 20036 6458
rect 19984 6394 20036 6400
rect 20088 6338 20116 7783
rect 20272 6458 20300 20742
rect 20364 19310 20392 20742
rect 20444 20528 20496 20534
rect 20444 20470 20496 20476
rect 20352 19304 20404 19310
rect 20352 19246 20404 19252
rect 20352 17332 20404 17338
rect 20352 17274 20404 17280
rect 20364 16794 20392 17274
rect 20456 17218 20484 20470
rect 20548 19378 20576 21286
rect 20640 21010 20668 21440
rect 20628 21004 20680 21010
rect 20628 20946 20680 20952
rect 20640 19854 20668 20946
rect 20824 20534 20852 23122
rect 20996 22636 21048 22642
rect 20996 22578 21048 22584
rect 21008 22030 21036 22578
rect 21100 22098 21128 29582
rect 22020 29306 22048 37198
rect 27724 37126 27752 39200
rect 27804 37256 27856 37262
rect 27804 37198 27856 37204
rect 28632 37256 28684 37262
rect 28632 37198 28684 37204
rect 22744 37120 22796 37126
rect 22744 37062 22796 37068
rect 23112 37120 23164 37126
rect 23112 37062 23164 37068
rect 25136 37120 25188 37126
rect 25136 37062 25188 37068
rect 27712 37120 27764 37126
rect 27712 37062 27764 37068
rect 22560 30728 22612 30734
rect 22560 30670 22612 30676
rect 22572 30394 22600 30670
rect 22560 30388 22612 30394
rect 22560 30330 22612 30336
rect 22008 29300 22060 29306
rect 22008 29242 22060 29248
rect 22100 28756 22152 28762
rect 22100 28698 22152 28704
rect 21916 28144 21968 28150
rect 21916 28086 21968 28092
rect 21180 26988 21232 26994
rect 21180 26930 21232 26936
rect 21192 26042 21220 26930
rect 21180 26036 21232 26042
rect 21180 25978 21232 25984
rect 21272 25968 21324 25974
rect 21272 25910 21324 25916
rect 21180 24200 21232 24206
rect 21180 24142 21232 24148
rect 21192 23322 21220 24142
rect 21284 23730 21312 25910
rect 21928 24954 21956 28086
rect 22112 27946 22140 28698
rect 22756 28082 22784 37062
rect 23124 30258 23152 37062
rect 24032 30660 24084 30666
rect 24032 30602 24084 30608
rect 23112 30252 23164 30258
rect 23112 30194 23164 30200
rect 23204 30048 23256 30054
rect 23204 29990 23256 29996
rect 22744 28076 22796 28082
rect 22744 28018 22796 28024
rect 23216 28014 23244 29990
rect 24044 29238 24072 30602
rect 24952 30388 25004 30394
rect 24952 30330 25004 30336
rect 24768 30252 24820 30258
rect 24768 30194 24820 30200
rect 24032 29232 24084 29238
rect 24032 29174 24084 29180
rect 23204 28008 23256 28014
rect 23204 27950 23256 27956
rect 22100 27940 22152 27946
rect 22100 27882 22152 27888
rect 23848 27396 23900 27402
rect 23848 27338 23900 27344
rect 23020 26240 23072 26246
rect 23020 26182 23072 26188
rect 23032 25974 23060 26182
rect 23020 25968 23072 25974
rect 23020 25910 23072 25916
rect 22836 25900 22888 25906
rect 22836 25842 22888 25848
rect 21916 24948 21968 24954
rect 21916 24890 21968 24896
rect 21928 24682 21956 24890
rect 22192 24880 22244 24886
rect 22192 24822 22244 24828
rect 21916 24676 21968 24682
rect 21916 24618 21968 24624
rect 22204 23866 22232 24822
rect 22652 24676 22704 24682
rect 22652 24618 22704 24624
rect 22560 24336 22612 24342
rect 22560 24278 22612 24284
rect 22192 23860 22244 23866
rect 22192 23802 22244 23808
rect 21272 23724 21324 23730
rect 21272 23666 21324 23672
rect 21180 23316 21232 23322
rect 21180 23258 21232 23264
rect 22008 23248 22060 23254
rect 22008 23190 22060 23196
rect 21272 23112 21324 23118
rect 21272 23054 21324 23060
rect 21284 22778 21312 23054
rect 21272 22772 21324 22778
rect 21272 22714 21324 22720
rect 22020 22574 22048 23190
rect 22100 22976 22152 22982
rect 22100 22918 22152 22924
rect 22008 22568 22060 22574
rect 22008 22510 22060 22516
rect 21088 22092 21140 22098
rect 21088 22034 21140 22040
rect 21824 22092 21876 22098
rect 21824 22034 21876 22040
rect 20996 22024 21048 22030
rect 20996 21966 21048 21972
rect 20812 20528 20864 20534
rect 20812 20470 20864 20476
rect 20628 19848 20680 19854
rect 20628 19790 20680 19796
rect 20720 19508 20772 19514
rect 20720 19450 20772 19456
rect 20536 19372 20588 19378
rect 20536 19314 20588 19320
rect 20548 17490 20576 19314
rect 20548 17462 20668 17490
rect 20456 17190 20576 17218
rect 20352 16788 20404 16794
rect 20352 16730 20404 16736
rect 20364 13938 20392 16730
rect 20444 16108 20496 16114
rect 20444 16050 20496 16056
rect 20456 15706 20484 16050
rect 20444 15700 20496 15706
rect 20444 15642 20496 15648
rect 20444 15360 20496 15366
rect 20444 15302 20496 15308
rect 20456 15094 20484 15302
rect 20444 15088 20496 15094
rect 20444 15030 20496 15036
rect 20444 14408 20496 14414
rect 20444 14350 20496 14356
rect 20456 13938 20484 14350
rect 20352 13932 20404 13938
rect 20352 13874 20404 13880
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20444 11892 20496 11898
rect 20444 11834 20496 11840
rect 20352 11756 20404 11762
rect 20352 11698 20404 11704
rect 20364 8498 20392 11698
rect 20456 9722 20484 11834
rect 20444 9716 20496 9722
rect 20444 9658 20496 9664
rect 20444 9580 20496 9586
rect 20444 9522 20496 9528
rect 20456 9194 20484 9522
rect 20548 9382 20576 17190
rect 20640 16590 20668 17462
rect 20732 17270 20760 19450
rect 20812 18760 20864 18766
rect 20812 18702 20864 18708
rect 20824 18426 20852 18702
rect 20812 18420 20864 18426
rect 20812 18362 20864 18368
rect 20720 17264 20772 17270
rect 20720 17206 20772 17212
rect 20720 16720 20772 16726
rect 20720 16662 20772 16668
rect 20628 16584 20680 16590
rect 20628 16526 20680 16532
rect 20732 16114 20760 16662
rect 20720 16108 20772 16114
rect 20720 16050 20772 16056
rect 20628 15904 20680 15910
rect 20628 15846 20680 15852
rect 20640 15162 20668 15846
rect 20824 15722 20852 18362
rect 20904 16448 20956 16454
rect 20904 16390 20956 16396
rect 20732 15694 20852 15722
rect 20732 15502 20760 15694
rect 20812 15632 20864 15638
rect 20812 15574 20864 15580
rect 20720 15496 20772 15502
rect 20720 15438 20772 15444
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20628 14272 20680 14278
rect 20628 14214 20680 14220
rect 20640 14006 20668 14214
rect 20732 14074 20760 15098
rect 20824 14074 20852 15574
rect 20720 14068 20772 14074
rect 20720 14010 20772 14016
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20628 14000 20680 14006
rect 20916 13954 20944 16390
rect 21008 16266 21036 21966
rect 21836 21418 21864 22034
rect 22112 21962 22140 22918
rect 22376 22704 22428 22710
rect 22376 22646 22428 22652
rect 22008 21956 22060 21962
rect 22008 21898 22060 21904
rect 22100 21956 22152 21962
rect 22100 21898 22152 21904
rect 22020 21690 22048 21898
rect 22192 21888 22244 21894
rect 22192 21830 22244 21836
rect 22008 21684 22060 21690
rect 22008 21626 22060 21632
rect 22204 21622 22232 21830
rect 22192 21616 22244 21622
rect 22192 21558 22244 21564
rect 22100 21480 22152 21486
rect 22100 21422 22152 21428
rect 21824 21412 21876 21418
rect 21824 21354 21876 21360
rect 21272 20596 21324 20602
rect 21272 20538 21324 20544
rect 21180 20256 21232 20262
rect 21180 20198 21232 20204
rect 21192 19514 21220 20198
rect 21180 19508 21232 19514
rect 21180 19450 21232 19456
rect 21008 16238 21128 16266
rect 21100 14362 21128 16238
rect 21180 16108 21232 16114
rect 21180 16050 21232 16056
rect 20628 13942 20680 13948
rect 20732 13926 20944 13954
rect 21008 14334 21128 14362
rect 20732 11762 20760 13926
rect 21008 13802 21036 14334
rect 20996 13796 21048 13802
rect 20996 13738 21048 13744
rect 21192 13682 21220 16050
rect 20824 13654 21220 13682
rect 20824 11762 20852 13654
rect 21284 13546 21312 20538
rect 21364 20392 21416 20398
rect 21364 20334 21416 20340
rect 21376 20058 21404 20334
rect 22112 20262 22140 21422
rect 22100 20256 22152 20262
rect 22100 20198 22152 20204
rect 21364 20052 21416 20058
rect 21364 19994 21416 20000
rect 22100 19372 22152 19378
rect 22100 19314 22152 19320
rect 22112 19174 22140 19314
rect 22100 19168 22152 19174
rect 22100 19110 22152 19116
rect 22388 18970 22416 22646
rect 22572 22574 22600 24278
rect 22664 24274 22692 24618
rect 22652 24268 22704 24274
rect 22652 24210 22704 24216
rect 22652 24064 22704 24070
rect 22652 24006 22704 24012
rect 22664 23798 22692 24006
rect 22652 23792 22704 23798
rect 22652 23734 22704 23740
rect 22560 22568 22612 22574
rect 22560 22510 22612 22516
rect 22376 18964 22428 18970
rect 22376 18906 22428 18912
rect 21548 18760 21600 18766
rect 21548 18702 21600 18708
rect 22284 18760 22336 18766
rect 22284 18702 22336 18708
rect 21364 18624 21416 18630
rect 21364 18566 21416 18572
rect 21376 18290 21404 18566
rect 21364 18284 21416 18290
rect 21364 18226 21416 18232
rect 21560 17882 21588 18702
rect 22008 18692 22060 18698
rect 22008 18634 22060 18640
rect 22020 18290 22048 18634
rect 22008 18284 22060 18290
rect 22008 18226 22060 18232
rect 22192 18216 22244 18222
rect 22192 18158 22244 18164
rect 22204 17882 22232 18158
rect 21548 17876 21600 17882
rect 21548 17818 21600 17824
rect 22192 17876 22244 17882
rect 22192 17818 22244 17824
rect 21456 17332 21508 17338
rect 21456 17274 21508 17280
rect 21364 17264 21416 17270
rect 21364 17206 21416 17212
rect 21376 16998 21404 17206
rect 21468 16998 21496 17274
rect 21364 16992 21416 16998
rect 21364 16934 21416 16940
rect 21456 16992 21508 16998
rect 21456 16934 21508 16940
rect 21364 16516 21416 16522
rect 21364 16458 21416 16464
rect 21376 13870 21404 16458
rect 22296 16182 22324 18702
rect 22468 17672 22520 17678
rect 22468 17614 22520 17620
rect 22480 16794 22508 17614
rect 22468 16788 22520 16794
rect 22468 16730 22520 16736
rect 22284 16176 22336 16182
rect 22284 16118 22336 16124
rect 22572 16130 22600 22510
rect 22848 22094 22876 25842
rect 23480 25832 23532 25838
rect 23480 25774 23532 25780
rect 23492 25430 23520 25774
rect 23480 25424 23532 25430
rect 23480 25366 23532 25372
rect 23664 22704 23716 22710
rect 23664 22646 23716 22652
rect 23676 22098 23704 22646
rect 22848 22066 22968 22094
rect 22940 22030 22968 22066
rect 23664 22092 23716 22098
rect 23664 22034 23716 22040
rect 22928 22024 22980 22030
rect 22928 21966 22980 21972
rect 22744 20324 22796 20330
rect 22744 20266 22796 20272
rect 22756 19922 22784 20266
rect 22744 19916 22796 19922
rect 22744 19858 22796 19864
rect 22652 19780 22704 19786
rect 22652 19722 22704 19728
rect 22664 19514 22692 19722
rect 22652 19508 22704 19514
rect 22652 19450 22704 19456
rect 22836 16992 22888 16998
rect 22836 16934 22888 16940
rect 22008 15428 22060 15434
rect 22008 15370 22060 15376
rect 21916 15360 21968 15366
rect 21916 15302 21968 15308
rect 21824 15020 21876 15026
rect 21824 14962 21876 14968
rect 21836 14414 21864 14962
rect 21824 14408 21876 14414
rect 21824 14350 21876 14356
rect 21732 13932 21784 13938
rect 21732 13874 21784 13880
rect 21364 13864 21416 13870
rect 21364 13806 21416 13812
rect 21364 13728 21416 13734
rect 21364 13670 21416 13676
rect 21456 13728 21508 13734
rect 21456 13670 21508 13676
rect 20996 13524 21048 13530
rect 20996 13466 21048 13472
rect 21192 13518 21312 13546
rect 20904 12096 20956 12102
rect 20904 12038 20956 12044
rect 20720 11756 20772 11762
rect 20720 11698 20772 11704
rect 20812 11756 20864 11762
rect 20812 11698 20864 11704
rect 20720 11348 20772 11354
rect 20720 11290 20772 11296
rect 20732 10810 20760 11290
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 20812 10668 20864 10674
rect 20812 10610 20864 10616
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 20732 9602 20760 9998
rect 20640 9574 20760 9602
rect 20824 9586 20852 10610
rect 20916 10606 20944 12038
rect 21008 11898 21036 13466
rect 21088 12844 21140 12850
rect 21088 12786 21140 12792
rect 21100 12102 21128 12786
rect 21088 12096 21140 12102
rect 21088 12038 21140 12044
rect 20996 11892 21048 11898
rect 20996 11834 21048 11840
rect 21192 11778 21220 13518
rect 21376 13326 21404 13670
rect 21468 13394 21496 13670
rect 21456 13388 21508 13394
rect 21456 13330 21508 13336
rect 21548 13388 21600 13394
rect 21548 13330 21600 13336
rect 21364 13320 21416 13326
rect 21364 13262 21416 13268
rect 21376 12442 21404 13262
rect 21560 13258 21588 13330
rect 21548 13252 21600 13258
rect 21548 13194 21600 13200
rect 21640 13184 21692 13190
rect 21640 13126 21692 13132
rect 21364 12436 21416 12442
rect 21364 12378 21416 12384
rect 21456 12164 21508 12170
rect 21456 12106 21508 12112
rect 21548 12164 21600 12170
rect 21548 12106 21600 12112
rect 21468 11898 21496 12106
rect 21456 11892 21508 11898
rect 21456 11834 21508 11840
rect 21008 11750 21220 11778
rect 21560 11762 21588 12106
rect 21548 11756 21600 11762
rect 20904 10600 20956 10606
rect 20904 10542 20956 10548
rect 20812 9580 20864 9586
rect 20536 9376 20588 9382
rect 20536 9318 20588 9324
rect 20456 9166 20576 9194
rect 20444 8628 20496 8634
rect 20444 8570 20496 8576
rect 20352 8492 20404 8498
rect 20352 8434 20404 8440
rect 20456 7857 20484 8570
rect 20442 7848 20498 7857
rect 20442 7783 20498 7792
rect 20260 6452 20312 6458
rect 20260 6394 20312 6400
rect 19904 6322 20116 6338
rect 19892 6316 20116 6322
rect 19944 6310 20116 6316
rect 19892 6258 19944 6264
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19340 5092 19392 5098
rect 19444 5086 19564 5114
rect 19340 5034 19392 5040
rect 19352 4690 19380 5034
rect 19536 5030 19564 5086
rect 20088 5030 20116 6310
rect 20168 5568 20220 5574
rect 20168 5510 20220 5516
rect 19432 5024 19484 5030
rect 19432 4966 19484 4972
rect 19524 5024 19576 5030
rect 19524 4966 19576 4972
rect 20076 5024 20128 5030
rect 20076 4966 20128 4972
rect 19340 4684 19392 4690
rect 19340 4626 19392 4632
rect 19248 4616 19300 4622
rect 19248 4558 19300 4564
rect 19064 4072 19116 4078
rect 19064 4014 19116 4020
rect 18696 3528 18748 3534
rect 18880 3528 18932 3534
rect 18696 3470 18748 3476
rect 18800 3488 18880 3516
rect 18800 2990 18828 3488
rect 18880 3470 18932 3476
rect 18972 3460 19024 3466
rect 18972 3402 19024 3408
rect 18984 3369 19012 3402
rect 18970 3360 19026 3369
rect 18970 3295 19026 3304
rect 18788 2984 18840 2990
rect 19076 2972 19104 4014
rect 19156 2984 19208 2990
rect 19076 2944 19156 2972
rect 18788 2926 18840 2932
rect 19156 2926 19208 2932
rect 18604 2916 18656 2922
rect 18604 2858 18656 2864
rect 18144 2440 18196 2446
rect 18144 2382 18196 2388
rect 18052 2304 18104 2310
rect 18052 2246 18104 2252
rect 17960 2100 18012 2106
rect 17960 2042 18012 2048
rect 18064 800 18092 2246
rect 19260 1902 19288 4558
rect 19444 2530 19472 4966
rect 19984 4752 20036 4758
rect 19984 4694 20036 4700
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19996 4282 20024 4694
rect 20088 4622 20116 4966
rect 20076 4616 20128 4622
rect 20076 4558 20128 4564
rect 19984 4276 20036 4282
rect 19984 4218 20036 4224
rect 20088 4146 20116 4558
rect 20180 4146 20208 5510
rect 20076 4140 20128 4146
rect 20076 4082 20128 4088
rect 20168 4140 20220 4146
rect 20168 4082 20220 4088
rect 19984 3392 20036 3398
rect 19984 3334 20036 3340
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19352 2502 19472 2530
rect 19996 2514 20024 3334
rect 20088 2666 20116 4082
rect 20442 3632 20498 3641
rect 20352 3596 20404 3602
rect 20442 3567 20498 3576
rect 20352 3538 20404 3544
rect 20168 3392 20220 3398
rect 20364 3369 20392 3538
rect 20456 3534 20484 3567
rect 20444 3528 20496 3534
rect 20444 3470 20496 3476
rect 20168 3334 20220 3340
rect 20350 3360 20406 3369
rect 20180 2854 20208 3334
rect 20350 3295 20406 3304
rect 20548 2854 20576 9166
rect 20640 8974 20668 9574
rect 20812 9522 20864 9528
rect 20628 8968 20680 8974
rect 20628 8910 20680 8916
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 20720 8832 20772 8838
rect 20720 8774 20772 8780
rect 20640 6934 20668 8774
rect 20732 7954 20760 8774
rect 20824 8498 20852 9522
rect 20916 8634 20944 10542
rect 20904 8628 20956 8634
rect 20904 8570 20956 8576
rect 20812 8492 20864 8498
rect 20812 8434 20864 8440
rect 21008 8022 21036 11750
rect 21548 11698 21600 11704
rect 21180 11688 21232 11694
rect 21180 11630 21232 11636
rect 21192 11150 21220 11630
rect 21560 11150 21588 11698
rect 21180 11144 21232 11150
rect 21180 11086 21232 11092
rect 21548 11144 21600 11150
rect 21548 11086 21600 11092
rect 21088 9648 21140 9654
rect 21088 9590 21140 9596
rect 21100 9382 21128 9590
rect 21088 9376 21140 9382
rect 21088 9318 21140 9324
rect 21192 9178 21220 11086
rect 21456 11008 21508 11014
rect 21456 10950 21508 10956
rect 21272 10532 21324 10538
rect 21272 10474 21324 10480
rect 21088 9172 21140 9178
rect 21088 9114 21140 9120
rect 21180 9172 21232 9178
rect 21180 9114 21232 9120
rect 21100 8634 21128 9114
rect 21284 9058 21312 10474
rect 21468 10470 21496 10950
rect 21560 10674 21588 11086
rect 21652 11082 21680 13126
rect 21744 12850 21772 13874
rect 21836 12850 21864 14350
rect 21928 14346 21956 15302
rect 21916 14340 21968 14346
rect 21916 14282 21968 14288
rect 22020 13326 22048 15370
rect 22008 13320 22060 13326
rect 21928 13268 22008 13274
rect 21928 13262 22060 13268
rect 21928 13246 22048 13262
rect 21928 13190 21956 13246
rect 21916 13184 21968 13190
rect 21916 13126 21968 13132
rect 22008 13184 22060 13190
rect 22008 13126 22060 13132
rect 21732 12844 21784 12850
rect 21732 12786 21784 12792
rect 21824 12844 21876 12850
rect 21824 12786 21876 12792
rect 21836 12238 21864 12786
rect 21824 12232 21876 12238
rect 21824 12174 21876 12180
rect 21732 11688 21784 11694
rect 21732 11630 21784 11636
rect 21640 11076 21692 11082
rect 21640 11018 21692 11024
rect 21548 10668 21600 10674
rect 21548 10610 21600 10616
rect 21364 10464 21416 10470
rect 21364 10406 21416 10412
rect 21456 10464 21508 10470
rect 21456 10406 21508 10412
rect 21376 9722 21404 10406
rect 21548 9988 21600 9994
rect 21548 9930 21600 9936
rect 21364 9716 21416 9722
rect 21364 9658 21416 9664
rect 21192 9030 21312 9058
rect 21088 8628 21140 8634
rect 21088 8570 21140 8576
rect 20812 8016 20864 8022
rect 20812 7958 20864 7964
rect 20996 8016 21048 8022
rect 20996 7958 21048 7964
rect 20720 7948 20772 7954
rect 20720 7890 20772 7896
rect 20628 6928 20680 6934
rect 20628 6870 20680 6876
rect 20824 6662 20852 7958
rect 21088 7404 21140 7410
rect 21088 7346 21140 7352
rect 20812 6656 20864 6662
rect 20812 6598 20864 6604
rect 20904 6248 20956 6254
rect 20904 6190 20956 6196
rect 20916 5642 20944 6190
rect 20994 5808 21050 5817
rect 20994 5743 20996 5752
rect 21048 5743 21050 5752
rect 20996 5714 21048 5720
rect 20904 5636 20956 5642
rect 20904 5578 20956 5584
rect 20628 5568 20680 5574
rect 20628 5510 20680 5516
rect 20640 5302 20668 5510
rect 20628 5296 20680 5302
rect 20628 5238 20680 5244
rect 20628 5160 20680 5166
rect 20628 5102 20680 5108
rect 20640 4758 20668 5102
rect 20718 4856 20774 4865
rect 20718 4791 20774 4800
rect 20628 4752 20680 4758
rect 20628 4694 20680 4700
rect 20732 3942 20760 4791
rect 20810 4176 20866 4185
rect 20810 4111 20866 4120
rect 20720 3936 20772 3942
rect 20720 3878 20772 3884
rect 20824 3126 20852 4111
rect 21100 3534 21128 7346
rect 21192 6118 21220 9030
rect 21272 8288 21324 8294
rect 21272 8230 21324 8236
rect 21180 6112 21232 6118
rect 21180 6054 21232 6060
rect 21284 5370 21312 8230
rect 21456 7472 21508 7478
rect 21376 7420 21456 7426
rect 21376 7414 21508 7420
rect 21376 7398 21496 7414
rect 21376 5642 21404 7398
rect 21560 6934 21588 9930
rect 21652 9382 21680 11018
rect 21640 9376 21692 9382
rect 21640 9318 21692 9324
rect 21652 8974 21680 9318
rect 21640 8968 21692 8974
rect 21640 8910 21692 8916
rect 21744 7410 21772 11630
rect 21836 8838 21864 12174
rect 21916 12096 21968 12102
rect 21916 12038 21968 12044
rect 21928 10742 21956 12038
rect 22020 11830 22048 13126
rect 22192 12708 22244 12714
rect 22192 12650 22244 12656
rect 22204 12594 22232 12650
rect 22112 12566 22232 12594
rect 22008 11824 22060 11830
rect 22008 11766 22060 11772
rect 21916 10736 21968 10742
rect 21916 10678 21968 10684
rect 22112 10130 22140 12566
rect 22100 10124 22152 10130
rect 22100 10066 22152 10072
rect 22100 9920 22152 9926
rect 22100 9862 22152 9868
rect 22112 9625 22140 9862
rect 21914 9616 21970 9625
rect 22098 9616 22154 9625
rect 21914 9551 21970 9560
rect 22008 9580 22060 9586
rect 21928 9450 21956 9551
rect 22098 9551 22154 9560
rect 22008 9522 22060 9528
rect 21916 9444 21968 9450
rect 21916 9386 21968 9392
rect 22020 9382 22048 9522
rect 22296 9489 22324 16118
rect 22572 16102 22784 16130
rect 22560 15904 22612 15910
rect 22560 15846 22612 15852
rect 22468 15496 22520 15502
rect 22468 15438 22520 15444
rect 22480 15026 22508 15438
rect 22468 15020 22520 15026
rect 22468 14962 22520 14968
rect 22480 14482 22508 14962
rect 22468 14476 22520 14482
rect 22468 14418 22520 14424
rect 22480 12434 22508 14418
rect 22572 12782 22600 15846
rect 22756 15706 22784 16102
rect 22744 15700 22796 15706
rect 22744 15642 22796 15648
rect 22848 14482 22876 16934
rect 22836 14476 22888 14482
rect 22836 14418 22888 14424
rect 22744 13932 22796 13938
rect 22744 13874 22796 13880
rect 22756 13258 22784 13874
rect 22744 13252 22796 13258
rect 22744 13194 22796 13200
rect 22560 12776 22612 12782
rect 22560 12718 22612 12724
rect 22388 12406 22508 12434
rect 22388 10742 22416 12406
rect 22756 12170 22784 13194
rect 22744 12164 22796 12170
rect 22744 12106 22796 12112
rect 22468 10804 22520 10810
rect 22468 10746 22520 10752
rect 22376 10736 22428 10742
rect 22376 10678 22428 10684
rect 22388 10062 22416 10678
rect 22376 10056 22428 10062
rect 22376 9998 22428 10004
rect 22282 9480 22338 9489
rect 22282 9415 22338 9424
rect 22008 9376 22060 9382
rect 22008 9318 22060 9324
rect 21916 8968 21968 8974
rect 21916 8910 21968 8916
rect 21824 8832 21876 8838
rect 21824 8774 21876 8780
rect 21928 7886 21956 8910
rect 22020 8242 22048 9318
rect 22388 9058 22416 9998
rect 22296 9030 22416 9058
rect 22192 8560 22244 8566
rect 22192 8502 22244 8508
rect 22020 8214 22140 8242
rect 22112 8090 22140 8214
rect 22100 8084 22152 8090
rect 22100 8026 22152 8032
rect 22098 7984 22154 7993
rect 22098 7919 22154 7928
rect 21916 7880 21968 7886
rect 21916 7822 21968 7828
rect 22008 7880 22060 7886
rect 22008 7822 22060 7828
rect 21732 7404 21784 7410
rect 21732 7346 21784 7352
rect 21640 7336 21692 7342
rect 21640 7278 21692 7284
rect 21652 7002 21680 7278
rect 21744 7177 21772 7346
rect 21730 7168 21786 7177
rect 21730 7103 21786 7112
rect 21730 7032 21786 7041
rect 21640 6996 21692 7002
rect 21730 6967 21732 6976
rect 21640 6938 21692 6944
rect 21784 6967 21786 6976
rect 21732 6938 21784 6944
rect 21548 6928 21600 6934
rect 21548 6870 21600 6876
rect 21928 6798 21956 7822
rect 22020 7410 22048 7822
rect 22008 7404 22060 7410
rect 22008 7346 22060 7352
rect 21916 6792 21968 6798
rect 21916 6734 21968 6740
rect 21456 6316 21508 6322
rect 21456 6258 21508 6264
rect 21468 6186 21496 6258
rect 21456 6180 21508 6186
rect 21456 6122 21508 6128
rect 21548 6112 21600 6118
rect 21548 6054 21600 6060
rect 21456 5840 21508 5846
rect 21456 5782 21508 5788
rect 21364 5636 21416 5642
rect 21364 5578 21416 5584
rect 21272 5364 21324 5370
rect 21272 5306 21324 5312
rect 21468 4729 21496 5782
rect 21560 5642 21588 6054
rect 21638 5808 21694 5817
rect 21638 5743 21640 5752
rect 21692 5743 21694 5752
rect 21640 5714 21692 5720
rect 21732 5704 21784 5710
rect 21732 5646 21784 5652
rect 21548 5636 21600 5642
rect 21548 5578 21600 5584
rect 21454 4720 21510 4729
rect 21454 4655 21510 4664
rect 21272 4140 21324 4146
rect 21272 4082 21324 4088
rect 21088 3528 21140 3534
rect 21088 3470 21140 3476
rect 21284 3194 21312 4082
rect 21560 4049 21588 5578
rect 21744 5030 21772 5646
rect 21732 5024 21784 5030
rect 21732 4966 21784 4972
rect 21928 4146 21956 6734
rect 22020 6322 22048 7346
rect 22008 6316 22060 6322
rect 22008 6258 22060 6264
rect 22112 5914 22140 7919
rect 22204 6662 22232 8502
rect 22296 7886 22324 9030
rect 22480 8090 22508 10746
rect 22756 9994 22784 12106
rect 22940 11626 22968 21966
rect 23480 21140 23532 21146
rect 23480 21082 23532 21088
rect 23492 20398 23520 21082
rect 23480 20392 23532 20398
rect 23480 20334 23532 20340
rect 23492 17542 23520 20334
rect 23572 18896 23624 18902
rect 23572 18838 23624 18844
rect 23480 17536 23532 17542
rect 23480 17478 23532 17484
rect 23584 17338 23612 18838
rect 23572 17332 23624 17338
rect 23572 17274 23624 17280
rect 23664 17264 23716 17270
rect 23664 17206 23716 17212
rect 23676 16794 23704 17206
rect 23860 17066 23888 27338
rect 23940 26784 23992 26790
rect 23940 26726 23992 26732
rect 23952 25974 23980 26726
rect 23940 25968 23992 25974
rect 23940 25910 23992 25916
rect 24044 20330 24072 29174
rect 24308 26852 24360 26858
rect 24308 26794 24360 26800
rect 24216 26444 24268 26450
rect 24216 26386 24268 26392
rect 24228 22710 24256 26386
rect 24320 25974 24348 26794
rect 24492 26512 24544 26518
rect 24492 26454 24544 26460
rect 24308 25968 24360 25974
rect 24308 25910 24360 25916
rect 24504 25838 24532 26454
rect 24780 26450 24808 30194
rect 24768 26444 24820 26450
rect 24768 26386 24820 26392
rect 24492 25832 24544 25838
rect 24492 25774 24544 25780
rect 24860 24200 24912 24206
rect 24860 24142 24912 24148
rect 24676 24064 24728 24070
rect 24676 24006 24728 24012
rect 24216 22704 24268 22710
rect 24216 22646 24268 22652
rect 24688 22098 24716 24006
rect 24872 23118 24900 24142
rect 24860 23112 24912 23118
rect 24860 23054 24912 23060
rect 24676 22092 24728 22098
rect 24964 22094 24992 30330
rect 25148 26994 25176 37062
rect 27528 31884 27580 31890
rect 27528 31826 27580 31832
rect 26792 31680 26844 31686
rect 26792 31622 26844 31628
rect 26148 31340 26200 31346
rect 26148 31282 26200 31288
rect 26160 29850 26188 31282
rect 26148 29844 26200 29850
rect 26148 29786 26200 29792
rect 26240 29640 26292 29646
rect 26240 29582 26292 29588
rect 25136 26988 25188 26994
rect 25136 26930 25188 26936
rect 25320 26988 25372 26994
rect 25320 26930 25372 26936
rect 25044 26784 25096 26790
rect 25044 26726 25096 26732
rect 25056 25362 25084 26726
rect 25332 26382 25360 26930
rect 25964 26920 26016 26926
rect 25964 26862 26016 26868
rect 25976 26450 26004 26862
rect 25964 26444 26016 26450
rect 25964 26386 26016 26392
rect 25320 26376 25372 26382
rect 25320 26318 25372 26324
rect 25044 25356 25096 25362
rect 25044 25298 25096 25304
rect 25136 25220 25188 25226
rect 25136 25162 25188 25168
rect 25148 24410 25176 25162
rect 25136 24404 25188 24410
rect 25136 24346 25188 24352
rect 24964 22066 25176 22094
rect 24676 22034 24728 22040
rect 24768 20868 24820 20874
rect 24768 20810 24820 20816
rect 24032 20324 24084 20330
rect 24032 20266 24084 20272
rect 24780 19990 24808 20810
rect 25148 20466 25176 22066
rect 25136 20460 25188 20466
rect 25136 20402 25188 20408
rect 24768 19984 24820 19990
rect 24768 19926 24820 19932
rect 25148 19378 25176 20402
rect 25136 19372 25188 19378
rect 25136 19314 25188 19320
rect 24768 18760 24820 18766
rect 24768 18702 24820 18708
rect 24584 18624 24636 18630
rect 24584 18566 24636 18572
rect 24596 18358 24624 18566
rect 24780 18426 24808 18702
rect 24768 18420 24820 18426
rect 24768 18362 24820 18368
rect 24584 18352 24636 18358
rect 24584 18294 24636 18300
rect 24860 18216 24912 18222
rect 24860 18158 24912 18164
rect 24400 18148 24452 18154
rect 24400 18090 24452 18096
rect 24124 17808 24176 17814
rect 24124 17750 24176 17756
rect 23848 17060 23900 17066
rect 23848 17002 23900 17008
rect 23664 16788 23716 16794
rect 23664 16730 23716 16736
rect 23296 16584 23348 16590
rect 23296 16526 23348 16532
rect 23308 16250 23336 16526
rect 23296 16244 23348 16250
rect 23296 16186 23348 16192
rect 23572 16108 23624 16114
rect 23572 16050 23624 16056
rect 23480 15428 23532 15434
rect 23480 15370 23532 15376
rect 23492 15162 23520 15370
rect 23480 15156 23532 15162
rect 23480 15098 23532 15104
rect 23480 15020 23532 15026
rect 23584 15008 23612 16050
rect 23664 15632 23716 15638
rect 23664 15574 23716 15580
rect 23532 14980 23612 15008
rect 23480 14962 23532 14968
rect 23204 14408 23256 14414
rect 23204 14350 23256 14356
rect 22928 11620 22980 11626
rect 22928 11562 22980 11568
rect 22836 10600 22888 10606
rect 22836 10542 22888 10548
rect 22744 9988 22796 9994
rect 22744 9930 22796 9936
rect 22560 9580 22612 9586
rect 22560 9522 22612 9528
rect 22572 8974 22600 9522
rect 22560 8968 22612 8974
rect 22560 8910 22612 8916
rect 22652 8900 22704 8906
rect 22652 8842 22704 8848
rect 22664 8566 22692 8842
rect 22652 8560 22704 8566
rect 22652 8502 22704 8508
rect 22468 8084 22520 8090
rect 22468 8026 22520 8032
rect 22560 8016 22612 8022
rect 22560 7958 22612 7964
rect 22284 7880 22336 7886
rect 22468 7880 22520 7886
rect 22284 7822 22336 7828
rect 22388 7840 22468 7868
rect 22388 7750 22416 7840
rect 22468 7822 22520 7828
rect 22376 7744 22428 7750
rect 22376 7686 22428 7692
rect 22572 6882 22600 7958
rect 22480 6854 22600 6882
rect 22192 6656 22244 6662
rect 22192 6598 22244 6604
rect 22100 5908 22152 5914
rect 22100 5850 22152 5856
rect 22376 5704 22428 5710
rect 22376 5646 22428 5652
rect 22388 5302 22416 5646
rect 22376 5296 22428 5302
rect 22376 5238 22428 5244
rect 22388 4622 22416 5238
rect 22480 5234 22508 6854
rect 22652 5704 22704 5710
rect 22756 5692 22784 9930
rect 22848 9722 22876 10542
rect 22836 9716 22888 9722
rect 22836 9658 22888 9664
rect 23216 6798 23244 14350
rect 23296 12368 23348 12374
rect 23296 12310 23348 12316
rect 23308 11150 23336 12310
rect 23492 11558 23520 14962
rect 23676 14482 23704 15574
rect 23860 15570 23888 17002
rect 23940 16040 23992 16046
rect 23940 15982 23992 15988
rect 23848 15564 23900 15570
rect 23848 15506 23900 15512
rect 23756 15360 23808 15366
rect 23756 15302 23808 15308
rect 23768 14618 23796 15302
rect 23756 14612 23808 14618
rect 23756 14554 23808 14560
rect 23664 14476 23716 14482
rect 23664 14418 23716 14424
rect 23768 14074 23796 14554
rect 23756 14068 23808 14074
rect 23756 14010 23808 14016
rect 23480 11552 23532 11558
rect 23480 11494 23532 11500
rect 23296 11144 23348 11150
rect 23296 11086 23348 11092
rect 23664 10736 23716 10742
rect 23664 10678 23716 10684
rect 23676 9722 23704 10678
rect 23952 10470 23980 15982
rect 24032 14272 24084 14278
rect 24032 14214 24084 14220
rect 24044 13938 24072 14214
rect 24032 13932 24084 13938
rect 24032 13874 24084 13880
rect 23940 10464 23992 10470
rect 23940 10406 23992 10412
rect 24032 10464 24084 10470
rect 24032 10406 24084 10412
rect 23952 10062 23980 10406
rect 24044 10198 24072 10406
rect 24032 10192 24084 10198
rect 24032 10134 24084 10140
rect 23940 10056 23992 10062
rect 23940 9998 23992 10004
rect 23664 9716 23716 9722
rect 23664 9658 23716 9664
rect 23480 9376 23532 9382
rect 23480 9318 23532 9324
rect 23386 9072 23442 9081
rect 23386 9007 23442 9016
rect 23400 8634 23428 9007
rect 23388 8628 23440 8634
rect 23388 8570 23440 8576
rect 23492 7274 23520 9318
rect 23572 8968 23624 8974
rect 23572 8910 23624 8916
rect 23584 8498 23612 8910
rect 23756 8900 23808 8906
rect 23756 8842 23808 8848
rect 23572 8492 23624 8498
rect 23572 8434 23624 8440
rect 23584 8362 23612 8434
rect 23572 8356 23624 8362
rect 23572 8298 23624 8304
rect 23664 8288 23716 8294
rect 23664 8230 23716 8236
rect 23676 7818 23704 8230
rect 23664 7812 23716 7818
rect 23664 7754 23716 7760
rect 23572 7744 23624 7750
rect 23572 7686 23624 7692
rect 23584 7478 23612 7686
rect 23572 7472 23624 7478
rect 23572 7414 23624 7420
rect 23664 7404 23716 7410
rect 23664 7346 23716 7352
rect 23480 7268 23532 7274
rect 23480 7210 23532 7216
rect 23386 7168 23442 7177
rect 23676 7154 23704 7346
rect 23386 7103 23442 7112
rect 23492 7126 23704 7154
rect 23296 6928 23348 6934
rect 23296 6870 23348 6876
rect 23204 6792 23256 6798
rect 23204 6734 23256 6740
rect 23020 6452 23072 6458
rect 23020 6394 23072 6400
rect 22928 6248 22980 6254
rect 22928 6190 22980 6196
rect 22704 5664 22784 5692
rect 22652 5646 22704 5652
rect 22940 5370 22968 6190
rect 23032 6118 23060 6394
rect 23204 6384 23256 6390
rect 23204 6326 23256 6332
rect 23020 6112 23072 6118
rect 23020 6054 23072 6060
rect 23216 5914 23244 6326
rect 23204 5908 23256 5914
rect 23204 5850 23256 5856
rect 23308 5846 23336 6870
rect 23400 6798 23428 7103
rect 23388 6792 23440 6798
rect 23388 6734 23440 6740
rect 23296 5840 23348 5846
rect 23296 5782 23348 5788
rect 23492 5710 23520 7126
rect 23572 6384 23624 6390
rect 23572 6326 23624 6332
rect 23480 5704 23532 5710
rect 23480 5646 23532 5652
rect 23492 5370 23520 5646
rect 22928 5364 22980 5370
rect 22928 5306 22980 5312
rect 23480 5364 23532 5370
rect 23480 5306 23532 5312
rect 22652 5296 22704 5302
rect 22652 5238 22704 5244
rect 22468 5228 22520 5234
rect 22468 5170 22520 5176
rect 22480 4690 22508 5170
rect 22468 4684 22520 4690
rect 22468 4626 22520 4632
rect 22376 4616 22428 4622
rect 22376 4558 22428 4564
rect 21916 4140 21968 4146
rect 21916 4082 21968 4088
rect 21546 4040 21602 4049
rect 21546 3975 21602 3984
rect 21362 3496 21418 3505
rect 21362 3431 21418 3440
rect 21376 3398 21404 3431
rect 21364 3392 21416 3398
rect 21364 3334 21416 3340
rect 21272 3188 21324 3194
rect 21272 3130 21324 3136
rect 20812 3120 20864 3126
rect 20812 3062 20864 3068
rect 21928 3058 21956 4082
rect 22192 3936 22244 3942
rect 22192 3878 22244 3884
rect 22204 3126 22232 3878
rect 22480 3534 22508 4626
rect 22664 4146 22692 5238
rect 23388 5160 23440 5166
rect 23388 5102 23440 5108
rect 23400 4690 23428 5102
rect 23388 4684 23440 4690
rect 23388 4626 23440 4632
rect 23492 4146 23520 5306
rect 22652 4140 22704 4146
rect 22652 4082 22704 4088
rect 23204 4140 23256 4146
rect 23204 4082 23256 4088
rect 23480 4140 23532 4146
rect 23480 4082 23532 4088
rect 22836 3936 22888 3942
rect 22836 3878 22888 3884
rect 22468 3528 22520 3534
rect 22468 3470 22520 3476
rect 22192 3120 22244 3126
rect 22192 3062 22244 3068
rect 21916 3052 21968 3058
rect 21916 2994 21968 3000
rect 22100 2984 22152 2990
rect 22100 2926 22152 2932
rect 20720 2916 20772 2922
rect 20720 2858 20772 2864
rect 20168 2848 20220 2854
rect 20168 2790 20220 2796
rect 20536 2848 20588 2854
rect 20536 2790 20588 2796
rect 20088 2638 20208 2666
rect 19984 2508 20036 2514
rect 19352 2446 19380 2502
rect 19984 2450 20036 2456
rect 20180 2446 20208 2638
rect 20732 2582 20760 2858
rect 22112 2650 22140 2926
rect 22100 2644 22152 2650
rect 22100 2586 22152 2592
rect 20720 2576 20772 2582
rect 20720 2518 20772 2524
rect 19340 2440 19392 2446
rect 19340 2382 19392 2388
rect 20168 2440 20220 2446
rect 20168 2382 20220 2388
rect 21272 2440 21324 2446
rect 21272 2382 21324 2388
rect 19340 2304 19392 2310
rect 19340 2246 19392 2252
rect 21180 2304 21232 2310
rect 21180 2246 21232 2252
rect 19248 1896 19300 1902
rect 19248 1838 19300 1844
rect 19352 800 19380 2246
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 21192 1902 21220 2246
rect 21180 1896 21232 1902
rect 21180 1838 21232 1844
rect 21284 800 21312 2382
rect 22560 2372 22612 2378
rect 22560 2314 22612 2320
rect 22572 800 22600 2314
rect 22848 2106 22876 3878
rect 23216 3534 23244 4082
rect 23480 4004 23532 4010
rect 23480 3946 23532 3952
rect 23204 3528 23256 3534
rect 23204 3470 23256 3476
rect 23492 3466 23520 3946
rect 23388 3460 23440 3466
rect 23388 3402 23440 3408
rect 23480 3460 23532 3466
rect 23480 3402 23532 3408
rect 23400 3194 23428 3402
rect 23388 3188 23440 3194
rect 23388 3130 23440 3136
rect 23584 3126 23612 6326
rect 23572 3120 23624 3126
rect 23572 3062 23624 3068
rect 23768 2650 23796 8842
rect 23848 8628 23900 8634
rect 23848 8570 23900 8576
rect 23860 7886 23888 8570
rect 24032 8492 24084 8498
rect 24032 8434 24084 8440
rect 23848 7880 23900 7886
rect 23848 7822 23900 7828
rect 24044 7410 24072 8434
rect 24032 7404 24084 7410
rect 24032 7346 24084 7352
rect 24136 6390 24164 17750
rect 24216 17604 24268 17610
rect 24216 17546 24268 17552
rect 24228 10198 24256 17546
rect 24216 10192 24268 10198
rect 24216 10134 24268 10140
rect 24216 8832 24268 8838
rect 24216 8774 24268 8780
rect 24124 6384 24176 6390
rect 24124 6326 24176 6332
rect 24228 6322 24256 8774
rect 24412 7478 24440 18090
rect 24872 17746 24900 18158
rect 24860 17740 24912 17746
rect 24860 17682 24912 17688
rect 24872 15026 24900 17682
rect 25136 17332 25188 17338
rect 25136 17274 25188 17280
rect 25044 15496 25096 15502
rect 25044 15438 25096 15444
rect 24860 15020 24912 15026
rect 24860 14962 24912 14968
rect 24872 12238 24900 14962
rect 25056 14414 25084 15438
rect 25044 14408 25096 14414
rect 25044 14350 25096 14356
rect 25044 13864 25096 13870
rect 25044 13806 25096 13812
rect 25056 13394 25084 13806
rect 25044 13388 25096 13394
rect 25044 13330 25096 13336
rect 24952 12776 25004 12782
rect 24952 12718 25004 12724
rect 24964 12442 24992 12718
rect 24952 12436 25004 12442
rect 24952 12378 25004 12384
rect 24860 12232 24912 12238
rect 24860 12174 24912 12180
rect 24676 11144 24728 11150
rect 24676 11086 24728 11092
rect 24688 8430 24716 11086
rect 24768 11008 24820 11014
rect 24768 10950 24820 10956
rect 24780 9994 24808 10950
rect 24768 9988 24820 9994
rect 24768 9930 24820 9936
rect 24768 9580 24820 9586
rect 24768 9522 24820 9528
rect 24676 8424 24728 8430
rect 24676 8366 24728 8372
rect 24400 7472 24452 7478
rect 24400 7414 24452 7420
rect 24216 6316 24268 6322
rect 24216 6258 24268 6264
rect 23848 5704 23900 5710
rect 23848 5646 23900 5652
rect 23860 3942 23888 5646
rect 24032 5228 24084 5234
rect 24032 5170 24084 5176
rect 23940 5024 23992 5030
rect 23940 4966 23992 4972
rect 23848 3936 23900 3942
rect 23848 3878 23900 3884
rect 23860 3398 23888 3878
rect 23848 3392 23900 3398
rect 23848 3334 23900 3340
rect 23756 2644 23808 2650
rect 23756 2586 23808 2592
rect 23848 2304 23900 2310
rect 23848 2246 23900 2252
rect 22836 2100 22888 2106
rect 22836 2042 22888 2048
rect 23860 800 23888 2246
rect 23952 1970 23980 4966
rect 24044 4758 24072 5170
rect 24032 4752 24084 4758
rect 24032 4694 24084 4700
rect 24228 3641 24256 6258
rect 24688 6186 24716 8366
rect 24780 7886 24808 9522
rect 24872 8566 24900 12174
rect 25044 11144 25096 11150
rect 25044 11086 25096 11092
rect 25056 10810 25084 11086
rect 25044 10804 25096 10810
rect 25044 10746 25096 10752
rect 24952 10192 25004 10198
rect 24952 10134 25004 10140
rect 24860 8560 24912 8566
rect 24860 8502 24912 8508
rect 24860 8424 24912 8430
rect 24860 8366 24912 8372
rect 24872 8090 24900 8366
rect 24860 8084 24912 8090
rect 24860 8026 24912 8032
rect 24768 7880 24820 7886
rect 24768 7822 24820 7828
rect 24780 7206 24808 7822
rect 24768 7200 24820 7206
rect 24768 7142 24820 7148
rect 24964 6254 24992 10134
rect 25044 10124 25096 10130
rect 25044 10066 25096 10072
rect 25056 8362 25084 10066
rect 25148 9926 25176 17274
rect 25332 14890 25360 26318
rect 26252 24274 26280 29582
rect 26424 28552 26476 28558
rect 26424 28494 26476 28500
rect 26332 26512 26384 26518
rect 26332 26454 26384 26460
rect 26344 25906 26372 26454
rect 26436 25974 26464 28494
rect 26804 27606 26832 31622
rect 27540 30802 27568 31826
rect 27816 31482 27844 37198
rect 28540 34536 28592 34542
rect 28540 34478 28592 34484
rect 27804 31476 27856 31482
rect 27804 31418 27856 31424
rect 27528 30796 27580 30802
rect 27528 30738 27580 30744
rect 28552 28218 28580 34478
rect 28644 32570 28672 37198
rect 28908 37188 28960 37194
rect 28908 37130 28960 37136
rect 28632 32564 28684 32570
rect 28632 32506 28684 32512
rect 28816 32428 28868 32434
rect 28816 32370 28868 32376
rect 28828 29850 28856 32370
rect 28816 29844 28868 29850
rect 28816 29786 28868 29792
rect 28540 28212 28592 28218
rect 28540 28154 28592 28160
rect 27804 28144 27856 28150
rect 27804 28086 27856 28092
rect 27160 27872 27212 27878
rect 27160 27814 27212 27820
rect 27252 27872 27304 27878
rect 27252 27814 27304 27820
rect 26792 27600 26844 27606
rect 26792 27542 26844 27548
rect 26608 27464 26660 27470
rect 26608 27406 26660 27412
rect 26620 27130 26648 27406
rect 26608 27124 26660 27130
rect 26608 27066 26660 27072
rect 27172 26450 27200 27814
rect 27264 27538 27292 27814
rect 27252 27532 27304 27538
rect 27252 27474 27304 27480
rect 27816 27334 27844 28086
rect 27988 28076 28040 28082
rect 27988 28018 28040 28024
rect 28000 27538 28028 28018
rect 27988 27532 28040 27538
rect 27988 27474 28040 27480
rect 27804 27328 27856 27334
rect 27804 27270 27856 27276
rect 27816 26586 27844 27270
rect 27804 26580 27856 26586
rect 27804 26522 27856 26528
rect 27160 26444 27212 26450
rect 27160 26386 27212 26392
rect 27528 26376 27580 26382
rect 27528 26318 27580 26324
rect 27540 26042 27568 26318
rect 27804 26308 27856 26314
rect 27804 26250 27856 26256
rect 27896 26308 27948 26314
rect 27896 26250 27948 26256
rect 27816 26042 27844 26250
rect 27528 26036 27580 26042
rect 27528 25978 27580 25984
rect 27804 26036 27856 26042
rect 27804 25978 27856 25984
rect 26424 25968 26476 25974
rect 27908 25922 27936 26250
rect 26424 25910 26476 25916
rect 27816 25906 27936 25922
rect 26332 25900 26384 25906
rect 26332 25842 26384 25848
rect 27804 25900 27936 25906
rect 27856 25894 27936 25900
rect 27804 25842 27856 25848
rect 27344 25832 27396 25838
rect 27344 25774 27396 25780
rect 27356 24954 27384 25774
rect 27712 25764 27764 25770
rect 27712 25706 27764 25712
rect 27620 25220 27672 25226
rect 27620 25162 27672 25168
rect 27344 24948 27396 24954
rect 27344 24890 27396 24896
rect 26240 24268 26292 24274
rect 26240 24210 26292 24216
rect 25964 24064 26016 24070
rect 25964 24006 26016 24012
rect 25872 22976 25924 22982
rect 25872 22918 25924 22924
rect 25884 22710 25912 22918
rect 25872 22704 25924 22710
rect 25872 22646 25924 22652
rect 25504 22568 25556 22574
rect 25504 22510 25556 22516
rect 25780 22568 25832 22574
rect 25780 22510 25832 22516
rect 25412 20800 25464 20806
rect 25412 20742 25464 20748
rect 25424 20534 25452 20742
rect 25412 20528 25464 20534
rect 25412 20470 25464 20476
rect 25516 16130 25544 22510
rect 25792 22098 25820 22510
rect 25780 22092 25832 22098
rect 25780 22034 25832 22040
rect 25688 22024 25740 22030
rect 25688 21966 25740 21972
rect 25700 21350 25728 21966
rect 25688 21344 25740 21350
rect 25688 21286 25740 21292
rect 25596 20936 25648 20942
rect 25596 20878 25648 20884
rect 25608 20602 25636 20878
rect 25596 20596 25648 20602
rect 25596 20538 25648 20544
rect 25700 20466 25728 21286
rect 25688 20460 25740 20466
rect 25688 20402 25740 20408
rect 25872 20256 25924 20262
rect 25872 20198 25924 20204
rect 25884 19786 25912 20198
rect 25688 19780 25740 19786
rect 25688 19722 25740 19728
rect 25872 19780 25924 19786
rect 25872 19722 25924 19728
rect 25700 19446 25728 19722
rect 25688 19440 25740 19446
rect 25688 19382 25740 19388
rect 25688 18284 25740 18290
rect 25688 18226 25740 18232
rect 25700 16522 25728 18226
rect 25976 18222 26004 24006
rect 26252 22094 26280 24210
rect 27252 23520 27304 23526
rect 27252 23462 27304 23468
rect 27160 23112 27212 23118
rect 27160 23054 27212 23060
rect 26424 23044 26476 23050
rect 26424 22986 26476 22992
rect 26252 22066 26372 22094
rect 26344 19922 26372 22066
rect 26436 22030 26464 22986
rect 27172 22234 27200 23054
rect 27160 22228 27212 22234
rect 27160 22170 27212 22176
rect 26424 22024 26476 22030
rect 26424 21966 26476 21972
rect 26332 19916 26384 19922
rect 26332 19858 26384 19864
rect 25964 18216 26016 18222
rect 25964 18158 26016 18164
rect 25872 17536 25924 17542
rect 25872 17478 25924 17484
rect 25688 16516 25740 16522
rect 25688 16458 25740 16464
rect 25424 16102 25544 16130
rect 25320 14884 25372 14890
rect 25320 14826 25372 14832
rect 25228 14816 25280 14822
rect 25228 14758 25280 14764
rect 25240 13938 25268 14758
rect 25228 13932 25280 13938
rect 25228 13874 25280 13880
rect 25424 12918 25452 16102
rect 25504 16040 25556 16046
rect 25504 15982 25556 15988
rect 25516 14074 25544 15982
rect 25780 15972 25832 15978
rect 25780 15914 25832 15920
rect 25792 15434 25820 15914
rect 25780 15428 25832 15434
rect 25780 15370 25832 15376
rect 25596 14408 25648 14414
rect 25596 14350 25648 14356
rect 25504 14068 25556 14074
rect 25504 14010 25556 14016
rect 25516 12986 25544 14010
rect 25504 12980 25556 12986
rect 25504 12922 25556 12928
rect 25412 12912 25464 12918
rect 25412 12854 25464 12860
rect 25320 11756 25372 11762
rect 25320 11698 25372 11704
rect 25332 11121 25360 11698
rect 25424 11354 25452 12854
rect 25504 12232 25556 12238
rect 25504 12174 25556 12180
rect 25412 11348 25464 11354
rect 25412 11290 25464 11296
rect 25318 11112 25374 11121
rect 25318 11047 25374 11056
rect 25228 10668 25280 10674
rect 25228 10610 25280 10616
rect 25240 10266 25268 10610
rect 25228 10260 25280 10266
rect 25228 10202 25280 10208
rect 25136 9920 25188 9926
rect 25136 9862 25188 9868
rect 25228 9512 25280 9518
rect 25228 9454 25280 9460
rect 25240 9110 25268 9454
rect 25228 9104 25280 9110
rect 25228 9046 25280 9052
rect 25044 8356 25096 8362
rect 25044 8298 25096 8304
rect 25516 6633 25544 12174
rect 25608 7002 25636 14350
rect 25596 6996 25648 7002
rect 25596 6938 25648 6944
rect 25688 6656 25740 6662
rect 25502 6624 25558 6633
rect 25688 6598 25740 6604
rect 25502 6559 25558 6568
rect 25320 6384 25372 6390
rect 25320 6326 25372 6332
rect 24952 6248 25004 6254
rect 24952 6190 25004 6196
rect 24676 6180 24728 6186
rect 24676 6122 24728 6128
rect 24584 5364 24636 5370
rect 24584 5306 24636 5312
rect 24596 5234 24624 5306
rect 24688 5234 24716 6122
rect 24584 5228 24636 5234
rect 24584 5170 24636 5176
rect 24676 5228 24728 5234
rect 24676 5170 24728 5176
rect 24676 5024 24728 5030
rect 24676 4966 24728 4972
rect 24768 5024 24820 5030
rect 24768 4966 24820 4972
rect 24688 4826 24716 4966
rect 24676 4820 24728 4826
rect 24676 4762 24728 4768
rect 24676 4684 24728 4690
rect 24676 4626 24728 4632
rect 24688 4146 24716 4626
rect 24780 4622 24808 4966
rect 25226 4720 25282 4729
rect 25226 4655 25282 4664
rect 25240 4622 25268 4655
rect 24768 4616 24820 4622
rect 24768 4558 24820 4564
rect 25228 4616 25280 4622
rect 25228 4558 25280 4564
rect 24780 4282 24808 4558
rect 25332 4554 25360 6326
rect 25412 5704 25464 5710
rect 25412 5646 25464 5652
rect 25424 5370 25452 5646
rect 25412 5364 25464 5370
rect 25412 5306 25464 5312
rect 25320 4548 25372 4554
rect 25320 4490 25372 4496
rect 24768 4276 24820 4282
rect 24768 4218 24820 4224
rect 24492 4140 24544 4146
rect 24492 4082 24544 4088
rect 24676 4140 24728 4146
rect 24676 4082 24728 4088
rect 24400 4072 24452 4078
rect 24400 4014 24452 4020
rect 24214 3632 24270 3641
rect 24214 3567 24270 3576
rect 24412 3466 24440 4014
rect 24504 3738 24532 4082
rect 25412 4004 25464 4010
rect 25412 3946 25464 3952
rect 24492 3732 24544 3738
rect 24492 3674 24544 3680
rect 24584 3528 24636 3534
rect 24584 3470 24636 3476
rect 24032 3460 24084 3466
rect 24032 3402 24084 3408
rect 24400 3460 24452 3466
rect 24400 3402 24452 3408
rect 24044 2990 24072 3402
rect 24124 3392 24176 3398
rect 24596 3369 24624 3470
rect 24124 3334 24176 3340
rect 24582 3360 24638 3369
rect 24136 3058 24164 3334
rect 24582 3295 24638 3304
rect 24124 3052 24176 3058
rect 24124 2994 24176 3000
rect 24032 2984 24084 2990
rect 24032 2926 24084 2932
rect 25424 2446 25452 3946
rect 25700 3738 25728 6598
rect 25884 5914 25912 17478
rect 25976 16046 26004 18158
rect 25964 16040 26016 16046
rect 25964 15982 26016 15988
rect 26436 14550 26464 21966
rect 27160 19780 27212 19786
rect 27160 19722 27212 19728
rect 27172 19514 27200 19722
rect 27160 19508 27212 19514
rect 27160 19450 27212 19456
rect 27264 17270 27292 23462
rect 27436 23316 27488 23322
rect 27436 23258 27488 23264
rect 27448 22642 27476 23258
rect 27632 22710 27660 25162
rect 27620 22704 27672 22710
rect 27620 22646 27672 22652
rect 27436 22636 27488 22642
rect 27436 22578 27488 22584
rect 27344 20256 27396 20262
rect 27344 20198 27396 20204
rect 27356 19378 27384 20198
rect 27344 19372 27396 19378
rect 27344 19314 27396 19320
rect 27252 17264 27304 17270
rect 27252 17206 27304 17212
rect 27448 17082 27476 22578
rect 27724 19922 27752 25706
rect 27816 23866 27844 25842
rect 28000 24886 28028 27474
rect 28920 27470 28948 37130
rect 29012 37126 29040 39200
rect 30300 37244 30328 39200
rect 32232 37262 32260 39200
rect 33520 37262 33548 39200
rect 30380 37256 30432 37262
rect 30300 37216 30380 37244
rect 30380 37198 30432 37204
rect 32220 37256 32272 37262
rect 32220 37198 32272 37204
rect 33508 37256 33560 37262
rect 33508 37198 33560 37204
rect 33876 37256 33928 37262
rect 33876 37198 33928 37204
rect 32128 37188 32180 37194
rect 32128 37130 32180 37136
rect 29000 37120 29052 37126
rect 29000 37062 29052 37068
rect 32140 34746 32168 37130
rect 32404 37120 32456 37126
rect 32404 37062 32456 37068
rect 33324 37120 33376 37126
rect 33324 37062 33376 37068
rect 32128 34740 32180 34746
rect 32128 34682 32180 34688
rect 31668 34604 31720 34610
rect 31668 34546 31720 34552
rect 31680 33114 31708 34546
rect 31668 33108 31720 33114
rect 31668 33050 31720 33056
rect 31116 32904 31168 32910
rect 31116 32846 31168 32852
rect 30472 31136 30524 31142
rect 30472 31078 30524 31084
rect 30484 29714 30512 31078
rect 30472 29708 30524 29714
rect 30472 29650 30524 29656
rect 29460 28416 29512 28422
rect 29460 28358 29512 28364
rect 29472 28082 29500 28358
rect 29460 28076 29512 28082
rect 29460 28018 29512 28024
rect 29644 28008 29696 28014
rect 29644 27950 29696 27956
rect 29656 27674 29684 27950
rect 29644 27668 29696 27674
rect 29644 27610 29696 27616
rect 28908 27464 28960 27470
rect 28908 27406 28960 27412
rect 28264 27328 28316 27334
rect 28264 27270 28316 27276
rect 27988 24880 28040 24886
rect 27988 24822 28040 24828
rect 28276 24750 28304 27270
rect 28448 25764 28500 25770
rect 28448 25706 28500 25712
rect 28460 25430 28488 25706
rect 28448 25424 28500 25430
rect 28448 25366 28500 25372
rect 28264 24744 28316 24750
rect 28264 24686 28316 24692
rect 27804 23860 27856 23866
rect 27804 23802 27856 23808
rect 28276 23186 28304 24686
rect 28448 24064 28500 24070
rect 28448 24006 28500 24012
rect 28264 23180 28316 23186
rect 28264 23122 28316 23128
rect 28356 23112 28408 23118
rect 28356 23054 28408 23060
rect 28264 22976 28316 22982
rect 28264 22918 28316 22924
rect 27896 22704 27948 22710
rect 27896 22646 27948 22652
rect 27908 22094 27936 22646
rect 28276 22094 28304 22918
rect 28368 22778 28396 23054
rect 28356 22772 28408 22778
rect 28356 22714 28408 22720
rect 28460 22642 28488 24006
rect 28540 23860 28592 23866
rect 28540 23802 28592 23808
rect 28448 22636 28500 22642
rect 28448 22578 28500 22584
rect 28552 22094 28580 23802
rect 29184 23724 29236 23730
rect 29184 23666 29236 23672
rect 29196 23322 29224 23666
rect 29276 23520 29328 23526
rect 29276 23462 29328 23468
rect 29184 23316 29236 23322
rect 29184 23258 29236 23264
rect 29288 23186 29316 23462
rect 29736 23248 29788 23254
rect 29736 23190 29788 23196
rect 29276 23180 29328 23186
rect 29276 23122 29328 23128
rect 28632 22568 28684 22574
rect 28632 22510 28684 22516
rect 28644 22234 28672 22510
rect 29000 22432 29052 22438
rect 29000 22374 29052 22380
rect 28632 22228 28684 22234
rect 28632 22170 28684 22176
rect 27908 22066 28028 22094
rect 28276 22066 28396 22094
rect 28552 22066 28672 22094
rect 27804 22024 27856 22030
rect 27804 21966 27856 21972
rect 27816 20942 27844 21966
rect 27804 20936 27856 20942
rect 27804 20878 27856 20884
rect 27712 19916 27764 19922
rect 27712 19858 27764 19864
rect 27724 18290 27752 19858
rect 27712 18284 27764 18290
rect 27712 18226 27764 18232
rect 27528 18216 27580 18222
rect 27528 18158 27580 18164
rect 27620 18216 27672 18222
rect 27620 18158 27672 18164
rect 27540 17882 27568 18158
rect 27528 17876 27580 17882
rect 27528 17818 27580 17824
rect 27632 17678 27660 18158
rect 27620 17672 27672 17678
rect 27620 17614 27672 17620
rect 27264 17054 27476 17082
rect 26516 15428 26568 15434
rect 26516 15370 26568 15376
rect 26424 14544 26476 14550
rect 26424 14486 26476 14492
rect 26240 13456 26292 13462
rect 26240 13398 26292 13404
rect 26252 12434 26280 13398
rect 26252 12406 26372 12434
rect 26344 12374 26372 12406
rect 26332 12368 26384 12374
rect 26332 12310 26384 12316
rect 25976 8622 26280 8650
rect 25976 8566 26004 8622
rect 26252 8566 26280 8622
rect 25964 8560 26016 8566
rect 25964 8502 26016 8508
rect 26148 8560 26200 8566
rect 26148 8502 26200 8508
rect 26240 8560 26292 8566
rect 26240 8502 26292 8508
rect 26160 8090 26188 8502
rect 26344 8430 26372 12310
rect 26528 11150 26556 15370
rect 27068 13864 27120 13870
rect 27068 13806 27120 13812
rect 26608 12844 26660 12850
rect 26608 12786 26660 12792
rect 26516 11144 26568 11150
rect 26516 11086 26568 11092
rect 26332 8424 26384 8430
rect 26332 8366 26384 8372
rect 26516 8356 26568 8362
rect 26516 8298 26568 8304
rect 26148 8084 26200 8090
rect 26148 8026 26200 8032
rect 26528 7342 26556 8298
rect 26516 7336 26568 7342
rect 26516 7278 26568 7284
rect 25964 6656 26016 6662
rect 25964 6598 26016 6604
rect 25976 6390 26004 6598
rect 25964 6384 26016 6390
rect 25964 6326 26016 6332
rect 25872 5908 25924 5914
rect 25872 5850 25924 5856
rect 26528 5302 26556 7278
rect 26516 5296 26568 5302
rect 26516 5238 26568 5244
rect 25872 5228 25924 5234
rect 25872 5170 25924 5176
rect 25884 4486 25912 5170
rect 26516 5092 26568 5098
rect 26516 5034 26568 5040
rect 26528 4622 26556 5034
rect 26516 4616 26568 4622
rect 26516 4558 26568 4564
rect 25780 4480 25832 4486
rect 25780 4422 25832 4428
rect 25872 4480 25924 4486
rect 25872 4422 25924 4428
rect 25792 4282 25820 4422
rect 25780 4276 25832 4282
rect 25780 4218 25832 4224
rect 26148 4140 26200 4146
rect 26148 4082 26200 4088
rect 25596 3732 25648 3738
rect 25596 3674 25648 3680
rect 25688 3732 25740 3738
rect 25688 3674 25740 3680
rect 25608 3466 25636 3674
rect 25596 3460 25648 3466
rect 25596 3402 25648 3408
rect 25700 2922 25728 3674
rect 25780 3528 25832 3534
rect 25780 3470 25832 3476
rect 25688 2916 25740 2922
rect 25688 2858 25740 2864
rect 25792 2774 25820 3470
rect 26160 3126 26188 4082
rect 26620 3738 26648 12786
rect 27080 12374 27108 13806
rect 27068 12368 27120 12374
rect 27068 12310 27120 12316
rect 26700 12232 26752 12238
rect 26700 12174 26752 12180
rect 26712 11354 26740 12174
rect 26700 11348 26752 11354
rect 26700 11290 26752 11296
rect 27160 8832 27212 8838
rect 27160 8774 27212 8780
rect 27172 8498 27200 8774
rect 27160 8492 27212 8498
rect 27160 8434 27212 8440
rect 27264 7274 27292 17054
rect 27344 16448 27396 16454
rect 27344 16390 27396 16396
rect 27356 16114 27384 16390
rect 27344 16108 27396 16114
rect 27344 16050 27396 16056
rect 27528 15496 27580 15502
rect 27528 15438 27580 15444
rect 27344 15360 27396 15366
rect 27344 15302 27396 15308
rect 27436 15360 27488 15366
rect 27436 15302 27488 15308
rect 27356 13938 27384 15302
rect 27344 13932 27396 13938
rect 27344 13874 27396 13880
rect 27448 13326 27476 15302
rect 27540 14618 27568 15438
rect 27528 14612 27580 14618
rect 27528 14554 27580 14560
rect 27436 13320 27488 13326
rect 27436 13262 27488 13268
rect 27344 7744 27396 7750
rect 27344 7686 27396 7692
rect 27356 7410 27384 7686
rect 27344 7404 27396 7410
rect 27344 7346 27396 7352
rect 27252 7268 27304 7274
rect 27252 7210 27304 7216
rect 27632 6905 27660 17614
rect 27896 17128 27948 17134
rect 27896 17070 27948 17076
rect 27804 14408 27856 14414
rect 27804 14350 27856 14356
rect 27712 14000 27764 14006
rect 27712 13942 27764 13948
rect 27724 12170 27752 13942
rect 27816 12850 27844 14350
rect 27908 12850 27936 17070
rect 28000 15094 28028 22066
rect 28080 21888 28132 21894
rect 28080 21830 28132 21836
rect 28092 21554 28120 21830
rect 28080 21548 28132 21554
rect 28080 21490 28132 21496
rect 28264 21480 28316 21486
rect 28264 21422 28316 21428
rect 28276 21146 28304 21422
rect 28264 21140 28316 21146
rect 28264 21082 28316 21088
rect 28172 20460 28224 20466
rect 28172 20402 28224 20408
rect 28184 19854 28212 20402
rect 28172 19848 28224 19854
rect 28172 19790 28224 19796
rect 28080 18624 28132 18630
rect 28080 18566 28132 18572
rect 28092 17746 28120 18566
rect 28264 18080 28316 18086
rect 28264 18022 28316 18028
rect 28276 17814 28304 18022
rect 28264 17808 28316 17814
rect 28264 17750 28316 17756
rect 28080 17740 28132 17746
rect 28080 17682 28132 17688
rect 27988 15088 28040 15094
rect 27988 15030 28040 15036
rect 27804 12844 27856 12850
rect 27804 12786 27856 12792
rect 27896 12844 27948 12850
rect 27896 12786 27948 12792
rect 27712 12164 27764 12170
rect 27712 12106 27764 12112
rect 27618 6896 27674 6905
rect 27618 6831 27674 6840
rect 27620 6384 27672 6390
rect 27620 6326 27672 6332
rect 27632 5914 27660 6326
rect 27620 5908 27672 5914
rect 27620 5850 27672 5856
rect 27436 5704 27488 5710
rect 27436 5646 27488 5652
rect 27068 3936 27120 3942
rect 27068 3878 27120 3884
rect 26608 3732 26660 3738
rect 26608 3674 26660 3680
rect 26424 3528 26476 3534
rect 26424 3470 26476 3476
rect 26148 3120 26200 3126
rect 26148 3062 26200 3068
rect 25516 2746 25820 2774
rect 25516 2650 25544 2746
rect 25504 2644 25556 2650
rect 25504 2586 25556 2592
rect 25412 2440 25464 2446
rect 25412 2382 25464 2388
rect 26148 2304 26200 2310
rect 26148 2246 26200 2252
rect 23940 1964 23992 1970
rect 23940 1906 23992 1912
rect 25792 870 25912 898
rect 25792 800 25820 870
rect 18 200 74 800
rect 1306 200 1362 800
rect 2594 200 2650 800
rect 4526 200 4582 800
rect 5814 200 5870 800
rect 7102 200 7158 800
rect 9034 200 9090 800
rect 10322 200 10378 800
rect 11610 200 11666 800
rect 13542 200 13598 800
rect 14830 200 14886 800
rect 16762 200 16818 800
rect 18050 200 18106 800
rect 19338 200 19394 800
rect 21270 200 21326 800
rect 22558 200 22614 800
rect 23846 200 23902 800
rect 25778 200 25834 800
rect 25884 762 25912 870
rect 26160 762 26188 2246
rect 26436 2038 26464 3470
rect 27080 3398 27108 3878
rect 27068 3392 27120 3398
rect 27068 3334 27120 3340
rect 27344 3392 27396 3398
rect 27344 3334 27396 3340
rect 27356 2961 27384 3334
rect 27342 2952 27398 2961
rect 27252 2916 27304 2922
rect 27342 2887 27398 2896
rect 27252 2858 27304 2864
rect 27068 2848 27120 2854
rect 27068 2790 27120 2796
rect 27080 2378 27108 2790
rect 27264 2774 27292 2858
rect 27172 2746 27292 2774
rect 27068 2372 27120 2378
rect 27068 2314 27120 2320
rect 26424 2032 26476 2038
rect 26424 1974 26476 1980
rect 27172 1442 27200 2746
rect 27448 2310 27476 5646
rect 27724 4758 27752 12106
rect 27816 10470 27844 12786
rect 28080 12164 28132 12170
rect 28080 12106 28132 12112
rect 28092 11354 28120 12106
rect 28080 11348 28132 11354
rect 28080 11290 28132 11296
rect 27804 10464 27856 10470
rect 27804 10406 27856 10412
rect 27988 8968 28040 8974
rect 27988 8910 28040 8916
rect 27804 6180 27856 6186
rect 27804 6122 27856 6128
rect 27712 4752 27764 4758
rect 27712 4694 27764 4700
rect 27816 3534 27844 6122
rect 28000 5778 28028 8910
rect 28276 8022 28304 17750
rect 28368 13870 28396 22066
rect 28448 18760 28500 18766
rect 28448 18702 28500 18708
rect 28460 18426 28488 18702
rect 28448 18420 28500 18426
rect 28448 18362 28500 18368
rect 28540 16176 28592 16182
rect 28540 16118 28592 16124
rect 28448 14000 28500 14006
rect 28448 13942 28500 13948
rect 28356 13864 28408 13870
rect 28356 13806 28408 13812
rect 28460 12986 28488 13942
rect 28552 13530 28580 16118
rect 28644 16046 28672 22066
rect 29012 21690 29040 22374
rect 29748 22098 29776 23190
rect 30380 22432 30432 22438
rect 30380 22374 30432 22380
rect 30392 22234 30420 22374
rect 30380 22228 30432 22234
rect 30380 22170 30432 22176
rect 29736 22092 29788 22098
rect 29736 22034 29788 22040
rect 29276 22024 29328 22030
rect 29276 21966 29328 21972
rect 29288 21690 29316 21966
rect 29736 21956 29788 21962
rect 29736 21898 29788 21904
rect 29000 21684 29052 21690
rect 29000 21626 29052 21632
rect 29276 21684 29328 21690
rect 29276 21626 29328 21632
rect 29184 21548 29236 21554
rect 29184 21490 29236 21496
rect 29000 20800 29052 20806
rect 29000 20742 29052 20748
rect 29012 20466 29040 20742
rect 29000 20460 29052 20466
rect 29000 20402 29052 20408
rect 29092 18216 29144 18222
rect 29092 18158 29144 18164
rect 29104 17678 29132 18158
rect 29092 17672 29144 17678
rect 29092 17614 29144 17620
rect 28632 16040 28684 16046
rect 28632 15982 28684 15988
rect 29000 14952 29052 14958
rect 29000 14894 29052 14900
rect 29012 13870 29040 14894
rect 29000 13864 29052 13870
rect 29000 13806 29052 13812
rect 28540 13524 28592 13530
rect 28540 13466 28592 13472
rect 29196 13462 29224 21490
rect 29748 20942 29776 21898
rect 30392 20942 30420 22170
rect 29736 20936 29788 20942
rect 29736 20878 29788 20884
rect 30380 20936 30432 20942
rect 30380 20878 30432 20884
rect 29368 20528 29420 20534
rect 29368 20470 29420 20476
rect 29380 20058 29408 20470
rect 29368 20052 29420 20058
rect 29368 19994 29420 20000
rect 29748 19854 29776 20878
rect 30484 20602 30512 29650
rect 30564 22976 30616 22982
rect 30564 22918 30616 22924
rect 30472 20596 30524 20602
rect 30472 20538 30524 20544
rect 29828 20324 29880 20330
rect 29828 20266 29880 20272
rect 29840 19990 29868 20266
rect 30104 20256 30156 20262
rect 30104 20198 30156 20204
rect 29828 19984 29880 19990
rect 29828 19926 29880 19932
rect 29736 19848 29788 19854
rect 29736 19790 29788 19796
rect 30116 19378 30144 20198
rect 30472 19916 30524 19922
rect 30472 19858 30524 19864
rect 30104 19372 30156 19378
rect 30104 19314 30156 19320
rect 29828 19304 29880 19310
rect 29828 19246 29880 19252
rect 29840 18834 29868 19246
rect 29828 18828 29880 18834
rect 29828 18770 29880 18776
rect 29276 16040 29328 16046
rect 29276 15982 29328 15988
rect 29184 13456 29236 13462
rect 29184 13398 29236 13404
rect 28448 12980 28500 12986
rect 28448 12922 28500 12928
rect 29288 12434 29316 15982
rect 30012 15904 30064 15910
rect 30012 15846 30064 15852
rect 30024 15434 30052 15846
rect 30012 15428 30064 15434
rect 30012 15370 30064 15376
rect 29460 15020 29512 15026
rect 29460 14962 29512 14968
rect 29472 14618 29500 14962
rect 29460 14612 29512 14618
rect 29460 14554 29512 14560
rect 29644 13320 29696 13326
rect 29644 13262 29696 13268
rect 29920 13320 29972 13326
rect 29920 13262 29972 13268
rect 29288 12406 29500 12434
rect 28724 12164 28776 12170
rect 28724 12106 28776 12112
rect 28736 11898 28764 12106
rect 29184 12096 29236 12102
rect 29184 12038 29236 12044
rect 28724 11892 28776 11898
rect 28724 11834 28776 11840
rect 28736 10674 28764 11834
rect 29196 11830 29224 12038
rect 29184 11824 29236 11830
rect 29184 11766 29236 11772
rect 29276 11688 29328 11694
rect 29276 11630 29328 11636
rect 29092 11552 29144 11558
rect 29092 11494 29144 11500
rect 29104 11150 29132 11494
rect 29092 11144 29144 11150
rect 29092 11086 29144 11092
rect 28724 10668 28776 10674
rect 28724 10610 28776 10616
rect 28724 9512 28776 9518
rect 28724 9454 28776 9460
rect 28736 9178 28764 9454
rect 28724 9172 28776 9178
rect 28724 9114 28776 9120
rect 28632 8968 28684 8974
rect 28632 8910 28684 8916
rect 28448 8832 28500 8838
rect 28448 8774 28500 8780
rect 28460 8498 28488 8774
rect 28644 8537 28672 8910
rect 28630 8528 28686 8537
rect 28448 8492 28500 8498
rect 28630 8463 28686 8472
rect 28448 8434 28500 8440
rect 28448 8288 28500 8294
rect 28448 8230 28500 8236
rect 28264 8016 28316 8022
rect 28264 7958 28316 7964
rect 28460 7818 28488 8230
rect 28632 7948 28684 7954
rect 28632 7890 28684 7896
rect 28448 7812 28500 7818
rect 28448 7754 28500 7760
rect 28172 6248 28224 6254
rect 28172 6190 28224 6196
rect 28184 5778 28212 6190
rect 28644 6186 28672 7890
rect 28724 7812 28776 7818
rect 28724 7754 28776 7760
rect 28736 6798 28764 7754
rect 29184 7472 29236 7478
rect 29184 7414 29236 7420
rect 29092 7336 29144 7342
rect 29092 7278 29144 7284
rect 28724 6792 28776 6798
rect 28724 6734 28776 6740
rect 28632 6180 28684 6186
rect 28632 6122 28684 6128
rect 27988 5772 28040 5778
rect 27988 5714 28040 5720
rect 28172 5772 28224 5778
rect 28172 5714 28224 5720
rect 27988 5228 28040 5234
rect 27988 5170 28040 5176
rect 28000 4826 28028 5170
rect 28080 5024 28132 5030
rect 28080 4966 28132 4972
rect 27988 4820 28040 4826
rect 27988 4762 28040 4768
rect 28092 4690 28120 4966
rect 28080 4684 28132 4690
rect 28080 4626 28132 4632
rect 27896 4616 27948 4622
rect 27896 4558 27948 4564
rect 27908 4282 27936 4558
rect 27896 4276 27948 4282
rect 27896 4218 27948 4224
rect 28172 4140 28224 4146
rect 28172 4082 28224 4088
rect 28184 3670 28212 4082
rect 28736 3942 28764 6734
rect 28908 6656 28960 6662
rect 28908 6598 28960 6604
rect 28920 6390 28948 6598
rect 28816 6384 28868 6390
rect 28816 6326 28868 6332
rect 28908 6384 28960 6390
rect 28908 6326 28960 6332
rect 28828 5914 28856 6326
rect 28816 5908 28868 5914
rect 28816 5850 28868 5856
rect 29000 5704 29052 5710
rect 29000 5646 29052 5652
rect 29012 5370 29040 5646
rect 29104 5370 29132 7278
rect 29196 6866 29224 7414
rect 29184 6860 29236 6866
rect 29184 6802 29236 6808
rect 29000 5364 29052 5370
rect 29000 5306 29052 5312
rect 29092 5364 29144 5370
rect 29092 5306 29144 5312
rect 29288 4146 29316 11630
rect 29368 10668 29420 10674
rect 29368 10610 29420 10616
rect 29380 8974 29408 10610
rect 29368 8968 29420 8974
rect 29368 8910 29420 8916
rect 29472 8820 29500 12406
rect 29380 8792 29500 8820
rect 29380 8566 29408 8792
rect 29368 8560 29420 8566
rect 29368 8502 29420 8508
rect 29380 7342 29408 8502
rect 29656 8090 29684 13262
rect 29932 12714 29960 13262
rect 29920 12708 29972 12714
rect 29920 12650 29972 12656
rect 30116 10674 30144 19314
rect 30380 17536 30432 17542
rect 30380 17478 30432 17484
rect 30196 17128 30248 17134
rect 30196 17070 30248 17076
rect 30208 16658 30236 17070
rect 30392 16658 30420 17478
rect 30196 16652 30248 16658
rect 30196 16594 30248 16600
rect 30380 16652 30432 16658
rect 30380 16594 30432 16600
rect 30380 16040 30432 16046
rect 30380 15982 30432 15988
rect 30392 15706 30420 15982
rect 30380 15700 30432 15706
rect 30380 15642 30432 15648
rect 30196 13864 30248 13870
rect 30196 13806 30248 13812
rect 30104 10668 30156 10674
rect 30104 10610 30156 10616
rect 29920 10600 29972 10606
rect 29920 10542 29972 10548
rect 29932 10266 29960 10542
rect 30012 10464 30064 10470
rect 30012 10406 30064 10412
rect 29920 10260 29972 10266
rect 29920 10202 29972 10208
rect 30024 10062 30052 10406
rect 30012 10056 30064 10062
rect 30012 9998 30064 10004
rect 29644 8084 29696 8090
rect 29644 8026 29696 8032
rect 30208 7410 30236 13806
rect 30484 13462 30512 19858
rect 30576 18902 30604 22918
rect 30656 22568 30708 22574
rect 30656 22510 30708 22516
rect 30668 22234 30696 22510
rect 31128 22506 31156 32846
rect 31760 30592 31812 30598
rect 31760 30534 31812 30540
rect 31772 25362 31800 30534
rect 32416 26994 32444 37062
rect 32956 32904 33008 32910
rect 32956 32846 33008 32852
rect 32968 30326 32996 32846
rect 33336 30734 33364 37062
rect 33416 35080 33468 35086
rect 33416 35022 33468 35028
rect 33324 30728 33376 30734
rect 33324 30670 33376 30676
rect 32956 30320 33008 30326
rect 32956 30262 33008 30268
rect 33324 30184 33376 30190
rect 33324 30126 33376 30132
rect 33140 28076 33192 28082
rect 33140 28018 33192 28024
rect 33152 27606 33180 28018
rect 33140 27600 33192 27606
rect 33140 27542 33192 27548
rect 32404 26988 32456 26994
rect 32404 26930 32456 26936
rect 31852 26784 31904 26790
rect 31852 26726 31904 26732
rect 31760 25356 31812 25362
rect 31760 25298 31812 25304
rect 31392 24200 31444 24206
rect 31392 24142 31444 24148
rect 31404 23118 31432 24142
rect 31392 23112 31444 23118
rect 31392 23054 31444 23060
rect 31864 23050 31892 26726
rect 32128 25424 32180 25430
rect 32128 25366 32180 25372
rect 31944 25288 31996 25294
rect 31944 25230 31996 25236
rect 31956 24410 31984 25230
rect 31944 24404 31996 24410
rect 31944 24346 31996 24352
rect 32140 23866 32168 25366
rect 33336 23866 33364 30126
rect 33428 30122 33456 35022
rect 33888 34746 33916 37198
rect 34808 37126 34836 39200
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 36740 37126 36768 39200
rect 37462 38176 37518 38185
rect 37462 38111 37518 38120
rect 37476 37330 37504 38111
rect 37464 37324 37516 37330
rect 37464 37266 37516 37272
rect 37740 37256 37792 37262
rect 37740 37198 37792 37204
rect 34796 37120 34848 37126
rect 34796 37062 34848 37068
rect 36728 37120 36780 37126
rect 36728 37062 36780 37068
rect 36910 36816 36966 36825
rect 36910 36751 36912 36760
rect 36964 36751 36966 36760
rect 37004 36780 37056 36786
rect 36912 36722 36964 36728
rect 37004 36722 37056 36728
rect 36728 36576 36780 36582
rect 36728 36518 36780 36524
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 33876 34740 33928 34746
rect 33876 34682 33928 34688
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 35440 32428 35492 32434
rect 35440 32370 35492 32376
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 33600 30252 33652 30258
rect 33600 30194 33652 30200
rect 33416 30116 33468 30122
rect 33416 30058 33468 30064
rect 33612 28762 33640 30194
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34520 29028 34572 29034
rect 34520 28970 34572 28976
rect 33600 28756 33652 28762
rect 33600 28698 33652 28704
rect 34532 28558 34560 28970
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34520 28552 34572 28558
rect 34520 28494 34572 28500
rect 35452 28218 35480 32370
rect 36740 31822 36768 36518
rect 37016 33114 37044 36722
rect 37280 36032 37332 36038
rect 37280 35974 37332 35980
rect 37004 33108 37056 33114
rect 37004 33050 37056 33056
rect 36728 31816 36780 31822
rect 36728 31758 36780 31764
rect 37292 31346 37320 35974
rect 37280 31340 37332 31346
rect 37280 31282 37332 31288
rect 35440 28212 35492 28218
rect 35440 28154 35492 28160
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 37752 26382 37780 37198
rect 38028 36174 38056 39200
rect 39316 36922 39344 39200
rect 39304 36916 39356 36922
rect 39304 36858 39356 36864
rect 38016 36168 38068 36174
rect 38016 36110 38068 36116
rect 38200 34944 38252 34950
rect 38200 34886 38252 34892
rect 38212 34785 38240 34886
rect 38198 34776 38254 34785
rect 38198 34711 38254 34720
rect 38292 33516 38344 33522
rect 38292 33458 38344 33464
rect 38304 33425 38332 33458
rect 38290 33416 38346 33425
rect 38290 33351 38346 33360
rect 38108 33312 38160 33318
rect 38108 33254 38160 33260
rect 37740 26376 37792 26382
rect 37740 26318 37792 26324
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 38120 25498 38148 33254
rect 38200 32224 38252 32230
rect 38200 32166 38252 32172
rect 38212 32065 38240 32166
rect 38198 32056 38254 32065
rect 38198 31991 38254 32000
rect 38200 30048 38252 30054
rect 38198 30016 38200 30025
rect 38252 30016 38254 30025
rect 38198 29951 38254 29960
rect 38292 29164 38344 29170
rect 38292 29106 38344 29112
rect 38304 28665 38332 29106
rect 38290 28656 38346 28665
rect 38290 28591 38346 28600
rect 38200 27328 38252 27334
rect 38198 27296 38200 27305
rect 38252 27296 38254 27305
rect 38198 27231 38254 27240
rect 38108 25492 38160 25498
rect 38108 25434 38160 25440
rect 38292 25288 38344 25294
rect 38290 25256 38292 25265
rect 38344 25256 38346 25265
rect 38290 25191 38346 25200
rect 38108 25152 38160 25158
rect 38108 25094 38160 25100
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 38120 24274 38148 25094
rect 38108 24268 38160 24274
rect 38108 24210 38160 24216
rect 38292 24200 38344 24206
rect 38292 24142 38344 24148
rect 33508 24064 33560 24070
rect 33508 24006 33560 24012
rect 37004 24064 37056 24070
rect 37004 24006 37056 24012
rect 32128 23860 32180 23866
rect 32128 23802 32180 23808
rect 33324 23860 33376 23866
rect 33324 23802 33376 23808
rect 31852 23044 31904 23050
rect 31852 22986 31904 22992
rect 31116 22500 31168 22506
rect 31116 22442 31168 22448
rect 30656 22228 30708 22234
rect 30656 22170 30708 22176
rect 31024 22024 31076 22030
rect 31024 21966 31076 21972
rect 31036 21690 31064 21966
rect 31024 21684 31076 21690
rect 31024 21626 31076 21632
rect 31484 20800 31536 20806
rect 31484 20742 31536 20748
rect 30748 20392 30800 20398
rect 30748 20334 30800 20340
rect 30760 20058 30788 20334
rect 30748 20052 30800 20058
rect 30748 19994 30800 20000
rect 31300 19712 31352 19718
rect 31300 19654 31352 19660
rect 31312 19310 31340 19654
rect 31300 19304 31352 19310
rect 31300 19246 31352 19252
rect 30564 18896 30616 18902
rect 30564 18838 30616 18844
rect 31208 18284 31260 18290
rect 31208 18226 31260 18232
rect 31024 18080 31076 18086
rect 31024 18022 31076 18028
rect 31036 17678 31064 18022
rect 31024 17672 31076 17678
rect 31024 17614 31076 17620
rect 31220 17610 31248 18226
rect 31208 17604 31260 17610
rect 31208 17546 31260 17552
rect 31116 17060 31168 17066
rect 31116 17002 31168 17008
rect 30564 16992 30616 16998
rect 30564 16934 30616 16940
rect 30576 16794 30604 16934
rect 30564 16788 30616 16794
rect 30564 16730 30616 16736
rect 30576 16250 30604 16730
rect 30564 16244 30616 16250
rect 30564 16186 30616 16192
rect 31024 15564 31076 15570
rect 31024 15506 31076 15512
rect 31036 14074 31064 15506
rect 31024 14068 31076 14074
rect 31024 14010 31076 14016
rect 30472 13456 30524 13462
rect 30472 13398 30524 13404
rect 30656 13252 30708 13258
rect 30656 13194 30708 13200
rect 30668 12442 30696 13194
rect 30932 13184 30984 13190
rect 30932 13126 30984 13132
rect 30944 12918 30972 13126
rect 30932 12912 30984 12918
rect 30932 12854 30984 12860
rect 31128 12782 31156 17002
rect 31220 15502 31248 17546
rect 31496 16114 31524 20742
rect 31484 16108 31536 16114
rect 31484 16050 31536 16056
rect 31208 15496 31260 15502
rect 31208 15438 31260 15444
rect 31760 14340 31812 14346
rect 31760 14282 31812 14288
rect 31772 13530 31800 14282
rect 31760 13524 31812 13530
rect 31760 13466 31812 13472
rect 31208 13456 31260 13462
rect 31208 13398 31260 13404
rect 30840 12776 30892 12782
rect 30840 12718 30892 12724
rect 31116 12776 31168 12782
rect 31116 12718 31168 12724
rect 30656 12436 30708 12442
rect 30656 12378 30708 12384
rect 30852 12306 30880 12718
rect 30840 12300 30892 12306
rect 30840 12242 30892 12248
rect 30380 10532 30432 10538
rect 30380 10474 30432 10480
rect 30392 7886 30420 10474
rect 30564 10464 30616 10470
rect 30564 10406 30616 10412
rect 30576 9586 30604 10406
rect 30564 9580 30616 9586
rect 30564 9522 30616 9528
rect 30576 8974 30604 9522
rect 30564 8968 30616 8974
rect 30564 8910 30616 8916
rect 31220 8566 31248 13398
rect 31864 13394 31892 22986
rect 32140 22642 32168 23802
rect 33520 23730 33548 24006
rect 32496 23724 32548 23730
rect 32496 23666 32548 23672
rect 33508 23724 33560 23730
rect 33508 23666 33560 23672
rect 32508 23322 32536 23666
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 32496 23316 32548 23322
rect 32496 23258 32548 23264
rect 37016 23118 37044 24006
rect 38304 23905 38332 24142
rect 38290 23896 38346 23905
rect 38290 23831 38346 23840
rect 37004 23112 37056 23118
rect 37004 23054 37056 23060
rect 32128 22636 32180 22642
rect 32128 22578 32180 22584
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 37464 22024 37516 22030
rect 37464 21966 37516 21972
rect 37740 22024 37792 22030
rect 37740 21966 37792 21972
rect 37476 21865 37504 21966
rect 37462 21856 37518 21865
rect 37462 21791 37518 21800
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34520 20800 34572 20806
rect 34520 20742 34572 20748
rect 34532 19922 34560 20742
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34520 19916 34572 19922
rect 34520 19858 34572 19864
rect 32588 19440 32640 19446
rect 32588 19382 32640 19388
rect 32404 17536 32456 17542
rect 32404 17478 32456 17484
rect 32416 17270 32444 17478
rect 32404 17264 32456 17270
rect 32404 17206 32456 17212
rect 32496 17264 32548 17270
rect 32496 17206 32548 17212
rect 32220 17128 32272 17134
rect 32220 17070 32272 17076
rect 31944 14340 31996 14346
rect 31944 14282 31996 14288
rect 31852 13388 31904 13394
rect 31852 13330 31904 13336
rect 31300 12776 31352 12782
rect 31300 12718 31352 12724
rect 31312 11150 31340 12718
rect 31956 12374 31984 14282
rect 32128 13320 32180 13326
rect 32128 13262 32180 13268
rect 32140 12442 32168 13262
rect 32128 12436 32180 12442
rect 32128 12378 32180 12384
rect 31944 12368 31996 12374
rect 31944 12310 31996 12316
rect 31852 12232 31904 12238
rect 31852 12174 31904 12180
rect 31864 11218 31892 12174
rect 32232 11830 32260 17070
rect 32508 16794 32536 17206
rect 32600 17134 32628 19382
rect 32680 19236 32732 19242
rect 32680 19178 32732 19184
rect 32588 17128 32640 17134
rect 32588 17070 32640 17076
rect 32496 16788 32548 16794
rect 32496 16730 32548 16736
rect 32692 12238 32720 19178
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35900 16992 35952 16998
rect 35900 16934 35952 16940
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 33232 16584 33284 16590
rect 33232 16526 33284 16532
rect 32864 15360 32916 15366
rect 32864 15302 32916 15308
rect 32876 14482 32904 15302
rect 32864 14476 32916 14482
rect 32864 14418 32916 14424
rect 33244 12306 33272 16526
rect 33508 15904 33560 15910
rect 33508 15846 33560 15852
rect 33520 15706 33548 15846
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 33508 15700 33560 15706
rect 33508 15642 33560 15648
rect 35912 15570 35940 16934
rect 35900 15564 35952 15570
rect 35900 15506 35952 15512
rect 34612 15496 34664 15502
rect 34612 15438 34664 15444
rect 34624 14618 34652 15438
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34612 14612 34664 14618
rect 34612 14554 34664 14560
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 36728 12844 36780 12850
rect 36728 12786 36780 12792
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 36740 12442 36768 12786
rect 36728 12436 36780 12442
rect 36728 12378 36780 12384
rect 33232 12300 33284 12306
rect 33232 12242 33284 12248
rect 32680 12232 32732 12238
rect 32680 12174 32732 12180
rect 32404 12096 32456 12102
rect 32404 12038 32456 12044
rect 32416 11830 32444 12038
rect 32220 11824 32272 11830
rect 32220 11766 32272 11772
rect 32404 11824 32456 11830
rect 32404 11766 32456 11772
rect 32496 11824 32548 11830
rect 32496 11766 32548 11772
rect 32508 11354 32536 11766
rect 32692 11694 32720 12174
rect 32680 11688 32732 11694
rect 32680 11630 32732 11636
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 32496 11348 32548 11354
rect 32496 11290 32548 11296
rect 31852 11212 31904 11218
rect 31852 11154 31904 11160
rect 31300 11144 31352 11150
rect 31300 11086 31352 11092
rect 33048 11076 33100 11082
rect 33048 11018 33100 11024
rect 33060 10674 33088 11018
rect 33048 10668 33100 10674
rect 33048 10610 33100 10616
rect 34796 10464 34848 10470
rect 34796 10406 34848 10412
rect 34808 8974 34836 10406
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 37752 9450 37780 21966
rect 38292 20936 38344 20942
rect 38292 20878 38344 20884
rect 38304 20505 38332 20878
rect 38290 20496 38346 20505
rect 38290 20431 38346 20440
rect 38292 17196 38344 17202
rect 38292 17138 38344 17144
rect 38304 17105 38332 17138
rect 38290 17096 38346 17105
rect 38290 17031 38346 17040
rect 38200 15904 38252 15910
rect 38200 15846 38252 15852
rect 38212 15745 38240 15846
rect 38198 15736 38254 15745
rect 38198 15671 38254 15680
rect 38292 14408 38344 14414
rect 38290 14376 38292 14385
rect 38344 14376 38346 14385
rect 38290 14311 38346 14320
rect 38108 13932 38160 13938
rect 38108 13874 38160 13880
rect 38120 11354 38148 13874
rect 38200 12640 38252 12646
rect 38200 12582 38252 12588
rect 38212 12345 38240 12582
rect 38198 12336 38254 12345
rect 38198 12271 38254 12280
rect 38108 11348 38160 11354
rect 38108 11290 38160 11296
rect 38292 11144 38344 11150
rect 38292 11086 38344 11092
rect 38304 10985 38332 11086
rect 38290 10976 38346 10985
rect 38290 10911 38346 10920
rect 37740 9444 37792 9450
rect 37740 9386 37792 9392
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34796 8968 34848 8974
rect 34796 8910 34848 8916
rect 38198 8936 38254 8945
rect 38198 8871 38254 8880
rect 38212 8838 38240 8871
rect 32496 8832 32548 8838
rect 32496 8774 32548 8780
rect 38200 8832 38252 8838
rect 38200 8774 38252 8780
rect 30564 8560 30616 8566
rect 30564 8502 30616 8508
rect 31208 8560 31260 8566
rect 31208 8502 31260 8508
rect 30576 8090 30604 8502
rect 32508 8498 32536 8774
rect 32496 8492 32548 8498
rect 32496 8434 32548 8440
rect 31760 8424 31812 8430
rect 31760 8366 31812 8372
rect 31772 8090 31800 8366
rect 34428 8356 34480 8362
rect 34428 8298 34480 8304
rect 30564 8084 30616 8090
rect 30564 8026 30616 8032
rect 31760 8084 31812 8090
rect 31760 8026 31812 8032
rect 30380 7880 30432 7886
rect 30380 7822 30432 7828
rect 33048 7880 33100 7886
rect 33048 7822 33100 7828
rect 30196 7404 30248 7410
rect 30196 7346 30248 7352
rect 29368 7336 29420 7342
rect 29368 7278 29420 7284
rect 31208 7200 31260 7206
rect 31208 7142 31260 7148
rect 30194 6896 30250 6905
rect 30194 6831 30250 6840
rect 30012 6316 30064 6322
rect 30012 6258 30064 6264
rect 30024 5914 30052 6258
rect 30012 5908 30064 5914
rect 30012 5850 30064 5856
rect 30208 5710 30236 6831
rect 30840 6452 30892 6458
rect 30840 6394 30892 6400
rect 30380 6384 30432 6390
rect 30380 6326 30432 6332
rect 30196 5704 30248 5710
rect 30196 5646 30248 5652
rect 29736 4548 29788 4554
rect 29736 4490 29788 4496
rect 29276 4140 29328 4146
rect 29276 4082 29328 4088
rect 28724 3936 28776 3942
rect 28724 3878 28776 3884
rect 29368 3936 29420 3942
rect 29368 3878 29420 3884
rect 28172 3664 28224 3670
rect 28172 3606 28224 3612
rect 29380 3602 29408 3878
rect 29368 3596 29420 3602
rect 29368 3538 29420 3544
rect 27804 3528 27856 3534
rect 27804 3470 27856 3476
rect 28080 3528 28132 3534
rect 28080 3470 28132 3476
rect 27896 3392 27948 3398
rect 27896 3334 27948 3340
rect 27908 3058 27936 3334
rect 27896 3052 27948 3058
rect 27896 2994 27948 3000
rect 27988 3052 28040 3058
rect 27988 2994 28040 3000
rect 27804 2848 27856 2854
rect 28000 2836 28028 2994
rect 27856 2808 28028 2836
rect 27804 2790 27856 2796
rect 28092 2650 28120 3470
rect 28540 3392 28592 3398
rect 28816 3392 28868 3398
rect 28540 3334 28592 3340
rect 28722 3360 28778 3369
rect 28552 3126 28580 3334
rect 28816 3334 28868 3340
rect 28722 3295 28778 3304
rect 28540 3120 28592 3126
rect 28540 3062 28592 3068
rect 28080 2644 28132 2650
rect 28080 2586 28132 2592
rect 28736 2446 28764 3295
rect 28828 3126 28856 3334
rect 28816 3120 28868 3126
rect 28816 3062 28868 3068
rect 29748 2650 29776 4490
rect 30208 4146 30236 5646
rect 30196 4140 30248 4146
rect 30196 4082 30248 4088
rect 29920 2848 29972 2854
rect 29920 2790 29972 2796
rect 30288 2848 30340 2854
rect 30288 2790 30340 2796
rect 29736 2644 29788 2650
rect 29736 2586 29788 2592
rect 29932 2446 29960 2790
rect 28724 2440 28776 2446
rect 28724 2382 28776 2388
rect 29920 2440 29972 2446
rect 29920 2382 29972 2388
rect 29000 2372 29052 2378
rect 29000 2314 29052 2320
rect 27436 2304 27488 2310
rect 27436 2246 27488 2252
rect 27080 1414 27200 1442
rect 27080 800 27108 1414
rect 29012 800 29040 2314
rect 30300 800 30328 2790
rect 30392 2446 30420 6326
rect 30656 6248 30708 6254
rect 30656 6190 30708 6196
rect 30668 5914 30696 6190
rect 30656 5908 30708 5914
rect 30656 5850 30708 5856
rect 30748 4072 30800 4078
rect 30748 4014 30800 4020
rect 30656 3936 30708 3942
rect 30656 3878 30708 3884
rect 30668 3602 30696 3878
rect 30656 3596 30708 3602
rect 30656 3538 30708 3544
rect 30760 2990 30788 4014
rect 30852 3738 30880 6394
rect 31220 5234 31248 7142
rect 31208 5228 31260 5234
rect 31208 5170 31260 5176
rect 32956 5024 33008 5030
rect 32956 4966 33008 4972
rect 32864 4616 32916 4622
rect 32864 4558 32916 4564
rect 31668 4004 31720 4010
rect 31668 3946 31720 3952
rect 30840 3732 30892 3738
rect 30840 3674 30892 3680
rect 31024 3528 31076 3534
rect 31024 3470 31076 3476
rect 31036 3194 31064 3470
rect 31208 3392 31260 3398
rect 31208 3334 31260 3340
rect 31576 3392 31628 3398
rect 31576 3334 31628 3340
rect 31024 3188 31076 3194
rect 31024 3130 31076 3136
rect 31220 3058 31248 3334
rect 31588 3126 31616 3334
rect 31576 3120 31628 3126
rect 31576 3062 31628 3068
rect 31208 3052 31260 3058
rect 31208 2994 31260 3000
rect 30748 2984 30800 2990
rect 30748 2926 30800 2932
rect 31680 2582 31708 3946
rect 32496 3052 32548 3058
rect 32496 2994 32548 3000
rect 31760 2848 31812 2854
rect 31760 2790 31812 2796
rect 32312 2848 32364 2854
rect 32312 2790 32364 2796
rect 31668 2576 31720 2582
rect 31668 2518 31720 2524
rect 31772 2514 31800 2790
rect 31760 2508 31812 2514
rect 31760 2450 31812 2456
rect 32324 2446 32352 2790
rect 32508 2650 32536 2994
rect 32876 2650 32904 4558
rect 32968 3126 32996 4966
rect 33060 3738 33088 7822
rect 33324 5092 33376 5098
rect 33324 5034 33376 5040
rect 33048 3732 33100 3738
rect 33048 3674 33100 3680
rect 32956 3120 33008 3126
rect 32956 3062 33008 3068
rect 32496 2644 32548 2650
rect 32496 2586 32548 2592
rect 32864 2644 32916 2650
rect 32864 2586 32916 2592
rect 33336 2514 33364 5034
rect 34440 4622 34468 8298
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 38292 7880 38344 7886
rect 38292 7822 38344 7828
rect 37280 7744 37332 7750
rect 37280 7686 37332 7692
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 36728 5296 36780 5302
rect 36728 5238 36780 5244
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34428 4616 34480 4622
rect 34428 4558 34480 4564
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 33692 3528 33744 3534
rect 33692 3470 33744 3476
rect 33704 2650 33732 3470
rect 36740 3194 36768 5238
rect 37292 3670 37320 7686
rect 38304 7585 38332 7822
rect 38290 7576 38346 7585
rect 38290 7511 38346 7520
rect 38292 6316 38344 6322
rect 38292 6258 38344 6264
rect 38304 6225 38332 6258
rect 38290 6216 38346 6225
rect 38290 6151 38346 6160
rect 38108 6112 38160 6118
rect 38108 6054 38160 6060
rect 38120 5710 38148 6054
rect 38108 5704 38160 5710
rect 38108 5646 38160 5652
rect 38200 4480 38252 4486
rect 38200 4422 38252 4428
rect 38212 4185 38240 4422
rect 38198 4176 38254 4185
rect 38198 4111 38254 4120
rect 37280 3664 37332 3670
rect 37280 3606 37332 3612
rect 38292 3528 38344 3534
rect 38292 3470 38344 3476
rect 36728 3188 36780 3194
rect 36728 3130 36780 3136
rect 38200 2848 38252 2854
rect 38304 2825 38332 3470
rect 39304 2984 39356 2990
rect 39304 2926 39356 2932
rect 38200 2790 38252 2796
rect 38290 2816 38346 2825
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 33692 2644 33744 2650
rect 33692 2586 33744 2592
rect 33324 2508 33376 2514
rect 33324 2450 33376 2456
rect 30380 2440 30432 2446
rect 30380 2382 30432 2388
rect 32312 2440 32364 2446
rect 32312 2382 32364 2388
rect 33508 2440 33560 2446
rect 33508 2382 33560 2388
rect 34796 2440 34848 2446
rect 34796 2382 34848 2388
rect 36084 2440 36136 2446
rect 36084 2382 36136 2388
rect 31576 2304 31628 2310
rect 31576 2246 31628 2252
rect 31588 800 31616 2246
rect 33520 800 33548 2382
rect 34808 800 34836 2382
rect 36096 800 36124 2382
rect 38016 2304 38068 2310
rect 38016 2246 38068 2252
rect 38028 800 38056 2246
rect 38212 1465 38240 2790
rect 38290 2751 38346 2760
rect 38198 1456 38254 1465
rect 38198 1391 38254 1400
rect 39316 800 39344 2926
rect 25884 734 26188 762
rect 27066 200 27122 800
rect 28998 200 29054 800
rect 30286 200 30342 800
rect 31574 200 31630 800
rect 33506 200 33562 800
rect 34794 200 34850 800
rect 36082 200 36138 800
rect 38014 200 38070 800
rect 39302 200 39358 800
<< via2 >>
rect 3146 38120 3202 38176
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 2778 36760 2834 36816
rect 1766 33360 1822 33416
rect 1766 32000 1822 32056
rect 1582 30676 1584 30696
rect 1584 30676 1636 30696
rect 1636 30676 1638 30696
rect 1582 30640 1638 30676
rect 1766 28600 1822 28656
rect 1766 27240 1822 27296
rect 1766 25236 1768 25256
rect 1768 25236 1820 25256
rect 1820 25236 1822 25256
rect 1766 25200 1822 25236
rect 1766 23840 1822 23896
rect 1766 22480 1822 22536
rect 1766 20440 1822 20496
rect 1766 19116 1768 19136
rect 1768 19116 1820 19136
rect 1820 19116 1822 19136
rect 1766 19080 1822 19116
rect 1766 17720 1822 17776
rect 1766 15680 1822 15736
rect 1766 14320 1822 14376
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 1766 12280 1822 12336
rect 1766 10920 1822 10976
rect 1766 9560 1822 9616
rect 1766 6160 1822 6216
rect 1766 4800 1822 4856
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 2778 7520 2834 7576
rect 1766 2760 1822 2816
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 5906 9016 5962 9072
rect 5170 5616 5226 5672
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 5354 4800 5410 4856
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 3330 2896 3386 2952
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 2778 1400 2834 1456
rect 10506 16124 10508 16144
rect 10508 16124 10560 16144
rect 10560 16124 10562 16144
rect 10506 16088 10562 16124
rect 10966 16088 11022 16144
rect 11978 18944 12034 19000
rect 11610 12588 11612 12608
rect 11612 12588 11664 12608
rect 11664 12588 11666 12608
rect 11610 12552 11666 12588
rect 11242 7928 11298 7984
rect 11150 4528 11206 4584
rect 12438 14900 12440 14920
rect 12440 14900 12492 14920
rect 12492 14900 12494 14920
rect 12438 14864 12494 14900
rect 12622 12588 12624 12608
rect 12624 12588 12676 12608
rect 12676 12588 12678 12608
rect 12622 12552 12678 12588
rect 14554 16516 14610 16552
rect 14554 16496 14556 16516
rect 14556 16496 14608 16516
rect 14608 16496 14610 16516
rect 15014 15308 15016 15328
rect 15016 15308 15068 15328
rect 15068 15308 15070 15328
rect 15014 15272 15070 15308
rect 14462 6840 14518 6896
rect 13634 5208 13690 5264
rect 13910 4120 13966 4176
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 16670 24112 16726 24168
rect 16026 15272 16082 15328
rect 17590 15136 17646 15192
rect 18234 18944 18290 19000
rect 18050 16516 18106 16552
rect 18050 16496 18052 16516
rect 18052 16496 18104 16516
rect 18104 16496 18106 16516
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 18694 15156 18750 15192
rect 18694 15136 18696 15156
rect 18696 15136 18748 15156
rect 18748 15136 18750 15156
rect 18602 14864 18658 14920
rect 14186 3304 14242 3360
rect 14370 3576 14426 3632
rect 14646 3440 14702 3496
rect 17866 7792 17922 7848
rect 16302 6976 16358 7032
rect 17682 4528 17738 4584
rect 17682 3984 17738 4040
rect 18326 7692 18328 7712
rect 18328 7692 18380 7712
rect 18380 7692 18382 7712
rect 18326 7656 18382 7692
rect 18418 6704 18474 6760
rect 18142 5636 18198 5672
rect 18142 5616 18144 5636
rect 18144 5616 18196 5636
rect 18196 5616 18198 5636
rect 18326 5344 18382 5400
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19154 9460 19156 9480
rect 19156 9460 19208 9480
rect 19208 9460 19210 9480
rect 19154 9424 19210 9460
rect 18602 5208 18658 5264
rect 17314 3612 17316 3632
rect 17316 3612 17368 3632
rect 17368 3612 17370 3632
rect 17314 3576 17370 3612
rect 19430 9424 19486 9480
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19706 8472 19762 8528
rect 19614 8336 19670 8392
rect 19982 8336 20038 8392
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 20074 7792 20130 7848
rect 20442 7792 20498 7848
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 18970 3304 19026 3360
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 20442 3576 20498 3632
rect 20350 3304 20406 3360
rect 20994 5772 21050 5808
rect 20994 5752 20996 5772
rect 20996 5752 21048 5772
rect 21048 5752 21050 5772
rect 20718 4800 20774 4856
rect 20810 4120 20866 4176
rect 21914 9560 21970 9616
rect 22098 9560 22154 9616
rect 22282 9424 22338 9480
rect 22098 7928 22154 7984
rect 21730 7112 21786 7168
rect 21730 6996 21786 7032
rect 21730 6976 21732 6996
rect 21732 6976 21784 6996
rect 21784 6976 21786 6996
rect 21638 5772 21694 5808
rect 21638 5752 21640 5772
rect 21640 5752 21692 5772
rect 21692 5752 21694 5772
rect 21454 4664 21510 4720
rect 23386 9016 23442 9072
rect 23386 7112 23442 7168
rect 21546 3984 21602 4040
rect 21362 3440 21418 3496
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 25318 11056 25374 11112
rect 25502 6568 25558 6624
rect 25226 4664 25282 4720
rect 24214 3576 24270 3632
rect 24582 3304 24638 3360
rect 27618 6840 27674 6896
rect 27342 2896 27398 2952
rect 28630 8472 28686 8528
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 37462 38120 37518 38176
rect 36910 36780 36966 36816
rect 36910 36760 36912 36780
rect 36912 36760 36964 36780
rect 36964 36760 36966 36780
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 38198 34720 38254 34776
rect 38290 33360 38346 33416
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 38198 32000 38254 32056
rect 38198 29996 38200 30016
rect 38200 29996 38252 30016
rect 38252 29996 38254 30016
rect 38198 29960 38254 29996
rect 38290 28600 38346 28656
rect 38198 27276 38200 27296
rect 38200 27276 38252 27296
rect 38252 27276 38254 27296
rect 38198 27240 38254 27276
rect 38290 25236 38292 25256
rect 38292 25236 38344 25256
rect 38344 25236 38346 25256
rect 38290 25200 38346 25236
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 38290 23840 38346 23896
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 37462 21800 37518 21856
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 38290 20440 38346 20496
rect 38290 17040 38346 17096
rect 38198 15680 38254 15736
rect 38290 14356 38292 14376
rect 38292 14356 38344 14376
rect 38344 14356 38346 14376
rect 38290 14320 38346 14356
rect 38198 12280 38254 12336
rect 38290 10920 38346 10976
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 38198 8880 38254 8936
rect 30194 6840 30250 6896
rect 28722 3304 28778 3360
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 38290 7520 38346 7576
rect 38290 6160 38346 6216
rect 38198 4120 38254 4176
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 38290 2760 38346 2816
rect 38198 1400 38254 1456
<< metal3 >>
rect 200 38178 800 38208
rect 3141 38178 3207 38181
rect 200 38176 3207 38178
rect 200 38120 3146 38176
rect 3202 38120 3207 38176
rect 200 38118 3207 38120
rect 200 38088 800 38118
rect 3141 38115 3207 38118
rect 37457 38178 37523 38181
rect 39200 38178 39800 38208
rect 37457 38176 39800 38178
rect 37457 38120 37462 38176
rect 37518 38120 39800 38176
rect 37457 38118 39800 38120
rect 37457 38115 37523 38118
rect 39200 38088 39800 38118
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 200 36818 800 36848
rect 2773 36818 2839 36821
rect 200 36816 2839 36818
rect 200 36760 2778 36816
rect 2834 36760 2839 36816
rect 200 36758 2839 36760
rect 200 36728 800 36758
rect 2773 36755 2839 36758
rect 36905 36818 36971 36821
rect 39200 36818 39800 36848
rect 36905 36816 39800 36818
rect 36905 36760 36910 36816
rect 36966 36760 39800 36816
rect 36905 36758 39800 36760
rect 36905 36755 36971 36758
rect 39200 36728 39800 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 200 35368 800 35488
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 38193 34778 38259 34781
rect 39200 34778 39800 34808
rect 38193 34776 39800 34778
rect 38193 34720 38198 34776
rect 38254 34720 39800 34776
rect 38193 34718 39800 34720
rect 38193 34715 38259 34718
rect 39200 34688 39800 34718
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 200 33418 800 33448
rect 1761 33418 1827 33421
rect 200 33416 1827 33418
rect 200 33360 1766 33416
rect 1822 33360 1827 33416
rect 200 33358 1827 33360
rect 200 33328 800 33358
rect 1761 33355 1827 33358
rect 38285 33418 38351 33421
rect 39200 33418 39800 33448
rect 38285 33416 39800 33418
rect 38285 33360 38290 33416
rect 38346 33360 39800 33416
rect 38285 33358 39800 33360
rect 38285 33355 38351 33358
rect 39200 33328 39800 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 200 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 1761 32058 1827 32061
rect 200 32056 1827 32058
rect 200 32000 1766 32056
rect 1822 32000 1827 32056
rect 200 31998 1827 32000
rect 200 31968 800 31998
rect 1761 31995 1827 31998
rect 38193 32058 38259 32061
rect 39200 32058 39800 32088
rect 38193 32056 39800 32058
rect 38193 32000 38198 32056
rect 38254 32000 39800 32056
rect 38193 31998 39800 32000
rect 38193 31995 38259 31998
rect 39200 31968 39800 31998
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 200 30698 800 30728
rect 1577 30698 1643 30701
rect 200 30696 1643 30698
rect 200 30640 1582 30696
rect 1638 30640 1643 30696
rect 200 30638 1643 30640
rect 200 30608 800 30638
rect 1577 30635 1643 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 38193 30018 38259 30021
rect 39200 30018 39800 30048
rect 38193 30016 39800 30018
rect 38193 29960 38198 30016
rect 38254 29960 39800 30016
rect 38193 29958 39800 29960
rect 38193 29955 38259 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 39200 29928 39800 29958
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 200 28658 800 28688
rect 1761 28658 1827 28661
rect 200 28656 1827 28658
rect 200 28600 1766 28656
rect 1822 28600 1827 28656
rect 200 28598 1827 28600
rect 200 28568 800 28598
rect 1761 28595 1827 28598
rect 38285 28658 38351 28661
rect 39200 28658 39800 28688
rect 38285 28656 39800 28658
rect 38285 28600 38290 28656
rect 38346 28600 39800 28656
rect 38285 28598 39800 28600
rect 38285 28595 38351 28598
rect 39200 28568 39800 28598
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 200 27298 800 27328
rect 1761 27298 1827 27301
rect 200 27296 1827 27298
rect 200 27240 1766 27296
rect 1822 27240 1827 27296
rect 200 27238 1827 27240
rect 200 27208 800 27238
rect 1761 27235 1827 27238
rect 38193 27298 38259 27301
rect 39200 27298 39800 27328
rect 38193 27296 39800 27298
rect 38193 27240 38198 27296
rect 38254 27240 39800 27296
rect 38193 27238 39800 27240
rect 38193 27235 38259 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 39200 27208 39800 27238
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 200 25258 800 25288
rect 1761 25258 1827 25261
rect 200 25256 1827 25258
rect 200 25200 1766 25256
rect 1822 25200 1827 25256
rect 200 25198 1827 25200
rect 200 25168 800 25198
rect 1761 25195 1827 25198
rect 38285 25258 38351 25261
rect 39200 25258 39800 25288
rect 38285 25256 39800 25258
rect 38285 25200 38290 25256
rect 38346 25200 39800 25256
rect 38285 25198 39800 25200
rect 38285 25195 38351 25198
rect 39200 25168 39800 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 16665 24170 16731 24173
rect 18270 24170 18276 24172
rect 16665 24168 18276 24170
rect 16665 24112 16670 24168
rect 16726 24112 18276 24168
rect 16665 24110 18276 24112
rect 16665 24107 16731 24110
rect 18270 24108 18276 24110
rect 18340 24108 18346 24172
rect 19570 23968 19886 23969
rect 200 23898 800 23928
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 1761 23898 1827 23901
rect 200 23896 1827 23898
rect 200 23840 1766 23896
rect 1822 23840 1827 23896
rect 200 23838 1827 23840
rect 200 23808 800 23838
rect 1761 23835 1827 23838
rect 38285 23898 38351 23901
rect 39200 23898 39800 23928
rect 38285 23896 39800 23898
rect 38285 23840 38290 23896
rect 38346 23840 39800 23896
rect 38285 23838 39800 23840
rect 38285 23835 38351 23838
rect 39200 23808 39800 23838
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 200 22538 800 22568
rect 1761 22538 1827 22541
rect 200 22536 1827 22538
rect 200 22480 1766 22536
rect 1822 22480 1827 22536
rect 200 22478 1827 22480
rect 200 22448 800 22478
rect 1761 22475 1827 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 37457 21858 37523 21861
rect 39200 21858 39800 21888
rect 37457 21856 39800 21858
rect 37457 21800 37462 21856
rect 37518 21800 39800 21856
rect 37457 21798 39800 21800
rect 37457 21795 37523 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 39200 21768 39800 21798
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 200 20498 800 20528
rect 1761 20498 1827 20501
rect 200 20496 1827 20498
rect 200 20440 1766 20496
rect 1822 20440 1827 20496
rect 200 20438 1827 20440
rect 200 20408 800 20438
rect 1761 20435 1827 20438
rect 38285 20498 38351 20501
rect 39200 20498 39800 20528
rect 38285 20496 39800 20498
rect 38285 20440 38290 20496
rect 38346 20440 39800 20496
rect 38285 20438 39800 20440
rect 38285 20435 38351 20438
rect 39200 20408 39800 20438
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 200 19138 800 19168
rect 1761 19138 1827 19141
rect 200 19136 1827 19138
rect 200 19080 1766 19136
rect 1822 19080 1827 19136
rect 200 19078 1827 19080
rect 200 19048 800 19078
rect 1761 19075 1827 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 39200 19048 39800 19168
rect 34930 19007 35246 19008
rect 11973 19002 12039 19005
rect 18229 19002 18295 19005
rect 11973 19000 18295 19002
rect 11973 18944 11978 19000
rect 12034 18944 18234 19000
rect 18290 18944 18295 19000
rect 11973 18942 18295 18944
rect 11973 18939 12039 18942
rect 18229 18939 18295 18942
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 200 17778 800 17808
rect 1761 17778 1827 17781
rect 200 17776 1827 17778
rect 200 17720 1766 17776
rect 1822 17720 1827 17776
rect 200 17718 1827 17720
rect 200 17688 800 17718
rect 1761 17715 1827 17718
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 38285 17098 38351 17101
rect 39200 17098 39800 17128
rect 38285 17096 39800 17098
rect 38285 17040 38290 17096
rect 38346 17040 39800 17096
rect 38285 17038 39800 17040
rect 38285 17035 38351 17038
rect 39200 17008 39800 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 14549 16554 14615 16557
rect 18045 16554 18111 16557
rect 14549 16552 18111 16554
rect 14549 16496 14554 16552
rect 14610 16496 18050 16552
rect 18106 16496 18111 16552
rect 14549 16494 18111 16496
rect 14549 16491 14615 16494
rect 18045 16491 18111 16494
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 10501 16146 10567 16149
rect 10961 16146 11027 16149
rect 10501 16144 11027 16146
rect 10501 16088 10506 16144
rect 10562 16088 10966 16144
rect 11022 16088 11027 16144
rect 10501 16086 11027 16088
rect 10501 16083 10567 16086
rect 10961 16083 11027 16086
rect 4210 15808 4526 15809
rect 200 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 1761 15738 1827 15741
rect 200 15736 1827 15738
rect 200 15680 1766 15736
rect 1822 15680 1827 15736
rect 200 15678 1827 15680
rect 200 15648 800 15678
rect 1761 15675 1827 15678
rect 38193 15738 38259 15741
rect 39200 15738 39800 15768
rect 38193 15736 39800 15738
rect 38193 15680 38198 15736
rect 38254 15680 39800 15736
rect 38193 15678 39800 15680
rect 38193 15675 38259 15678
rect 39200 15648 39800 15678
rect 15009 15330 15075 15333
rect 16021 15330 16087 15333
rect 15009 15328 16087 15330
rect 15009 15272 15014 15328
rect 15070 15272 16026 15328
rect 16082 15272 16087 15328
rect 15009 15270 16087 15272
rect 15009 15267 15075 15270
rect 16021 15267 16087 15270
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 17585 15194 17651 15197
rect 18689 15194 18755 15197
rect 17585 15192 18755 15194
rect 17585 15136 17590 15192
rect 17646 15136 18694 15192
rect 18750 15136 18755 15192
rect 17585 15134 18755 15136
rect 17585 15131 17651 15134
rect 18689 15131 18755 15134
rect 12433 14922 12499 14925
rect 18597 14922 18663 14925
rect 12433 14920 18663 14922
rect 12433 14864 12438 14920
rect 12494 14864 18602 14920
rect 18658 14864 18663 14920
rect 12433 14862 18663 14864
rect 12433 14859 12499 14862
rect 18597 14859 18663 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 200 14378 800 14408
rect 1761 14378 1827 14381
rect 200 14376 1827 14378
rect 200 14320 1766 14376
rect 1822 14320 1827 14376
rect 200 14318 1827 14320
rect 200 14288 800 14318
rect 1761 14315 1827 14318
rect 38285 14378 38351 14381
rect 39200 14378 39800 14408
rect 38285 14376 39800 14378
rect 38285 14320 38290 14376
rect 38346 14320 39800 14376
rect 38285 14318 39800 14320
rect 38285 14315 38351 14318
rect 39200 14288 39800 14318
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 11605 12610 11671 12613
rect 12617 12610 12683 12613
rect 11605 12608 12683 12610
rect 11605 12552 11610 12608
rect 11666 12552 12622 12608
rect 12678 12552 12683 12608
rect 11605 12550 12683 12552
rect 11605 12547 11671 12550
rect 12617 12547 12683 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 200 12338 800 12368
rect 1761 12338 1827 12341
rect 200 12336 1827 12338
rect 200 12280 1766 12336
rect 1822 12280 1827 12336
rect 200 12278 1827 12280
rect 200 12248 800 12278
rect 1761 12275 1827 12278
rect 38193 12338 38259 12341
rect 39200 12338 39800 12368
rect 38193 12336 39800 12338
rect 38193 12280 38198 12336
rect 38254 12280 39800 12336
rect 38193 12278 39800 12280
rect 38193 12275 38259 12278
rect 39200 12248 39800 12278
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 18454 11052 18460 11116
rect 18524 11114 18530 11116
rect 25313 11114 25379 11117
rect 18524 11112 25379 11114
rect 18524 11056 25318 11112
rect 25374 11056 25379 11112
rect 18524 11054 25379 11056
rect 18524 11052 18530 11054
rect 25313 11051 25379 11054
rect 200 10978 800 11008
rect 1761 10978 1827 10981
rect 200 10976 1827 10978
rect 200 10920 1766 10976
rect 1822 10920 1827 10976
rect 200 10918 1827 10920
rect 200 10888 800 10918
rect 1761 10915 1827 10918
rect 38285 10978 38351 10981
rect 39200 10978 39800 11008
rect 38285 10976 39800 10978
rect 38285 10920 38290 10976
rect 38346 10920 39800 10976
rect 38285 10918 39800 10920
rect 38285 10915 38351 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 39200 10888 39800 10918
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 200 9618 800 9648
rect 1761 9618 1827 9621
rect 200 9616 1827 9618
rect 200 9560 1766 9616
rect 1822 9560 1827 9616
rect 200 9558 1827 9560
rect 200 9528 800 9558
rect 1761 9555 1827 9558
rect 21909 9618 21975 9621
rect 22093 9618 22159 9621
rect 21909 9616 22159 9618
rect 21909 9560 21914 9616
rect 21970 9560 22098 9616
rect 22154 9560 22159 9616
rect 21909 9558 22159 9560
rect 21909 9555 21975 9558
rect 22093 9555 22159 9558
rect 19149 9482 19215 9485
rect 19425 9482 19491 9485
rect 22277 9482 22343 9485
rect 19149 9480 22343 9482
rect 19149 9424 19154 9480
rect 19210 9424 19430 9480
rect 19486 9424 22282 9480
rect 22338 9424 22343 9480
rect 19149 9422 22343 9424
rect 19149 9419 19215 9422
rect 19425 9419 19491 9422
rect 22277 9419 22343 9422
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 5901 9074 5967 9077
rect 23381 9074 23447 9077
rect 5901 9072 23447 9074
rect 5901 9016 5906 9072
rect 5962 9016 23386 9072
rect 23442 9016 23447 9072
rect 5901 9014 23447 9016
rect 5901 9011 5967 9014
rect 23381 9011 23447 9014
rect 38193 8938 38259 8941
rect 39200 8938 39800 8968
rect 38193 8936 39800 8938
rect 38193 8880 38198 8936
rect 38254 8880 39800 8936
rect 38193 8878 39800 8880
rect 38193 8875 38259 8878
rect 39200 8848 39800 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 19701 8530 19767 8533
rect 28625 8530 28691 8533
rect 19701 8528 28691 8530
rect 19701 8472 19706 8528
rect 19762 8472 28630 8528
rect 28686 8472 28691 8528
rect 19701 8470 28691 8472
rect 19701 8467 19767 8470
rect 28625 8467 28691 8470
rect 19609 8394 19675 8397
rect 19977 8394 20043 8397
rect 19609 8392 20043 8394
rect 19609 8336 19614 8392
rect 19670 8336 19982 8392
rect 20038 8336 20043 8392
rect 19609 8334 20043 8336
rect 19609 8331 19675 8334
rect 19977 8331 20043 8334
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 11237 7986 11303 7989
rect 22093 7986 22159 7989
rect 11237 7984 22159 7986
rect 11237 7928 11242 7984
rect 11298 7928 22098 7984
rect 22154 7928 22159 7984
rect 11237 7926 22159 7928
rect 11237 7923 11303 7926
rect 22093 7923 22159 7926
rect 17861 7850 17927 7853
rect 20069 7850 20135 7853
rect 20437 7850 20503 7853
rect 17861 7848 20503 7850
rect 17861 7792 17866 7848
rect 17922 7792 20074 7848
rect 20130 7792 20442 7848
rect 20498 7792 20503 7848
rect 17861 7790 20503 7792
rect 17861 7787 17927 7790
rect 20069 7787 20135 7790
rect 20437 7787 20503 7790
rect 18321 7714 18387 7717
rect 18454 7714 18460 7716
rect 18321 7712 18460 7714
rect 18321 7656 18326 7712
rect 18382 7656 18460 7712
rect 18321 7654 18460 7656
rect 18321 7651 18387 7654
rect 18454 7652 18460 7654
rect 18524 7652 18530 7716
rect 19570 7648 19886 7649
rect 200 7578 800 7608
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 2773 7578 2839 7581
rect 200 7576 2839 7578
rect 200 7520 2778 7576
rect 2834 7520 2839 7576
rect 200 7518 2839 7520
rect 200 7488 800 7518
rect 2773 7515 2839 7518
rect 38285 7578 38351 7581
rect 39200 7578 39800 7608
rect 38285 7576 39800 7578
rect 38285 7520 38290 7576
rect 38346 7520 39800 7576
rect 38285 7518 39800 7520
rect 38285 7515 38351 7518
rect 39200 7488 39800 7518
rect 21725 7170 21791 7173
rect 23381 7170 23447 7173
rect 21725 7168 23447 7170
rect 21725 7112 21730 7168
rect 21786 7112 23386 7168
rect 23442 7112 23447 7168
rect 21725 7110 23447 7112
rect 21725 7107 21791 7110
rect 23381 7107 23447 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 16297 7034 16363 7037
rect 21725 7034 21791 7037
rect 16297 7032 21791 7034
rect 16297 6976 16302 7032
rect 16358 6976 21730 7032
rect 21786 6976 21791 7032
rect 16297 6974 21791 6976
rect 16297 6971 16363 6974
rect 21725 6971 21791 6974
rect 14457 6898 14523 6901
rect 27613 6898 27679 6901
rect 30189 6898 30255 6901
rect 14457 6896 30255 6898
rect 14457 6840 14462 6896
rect 14518 6840 27618 6896
rect 27674 6840 30194 6896
rect 30250 6840 30255 6896
rect 14457 6838 30255 6840
rect 14457 6835 14523 6838
rect 27613 6835 27679 6838
rect 30189 6835 30255 6838
rect 18413 6762 18479 6765
rect 18413 6760 20730 6762
rect 18413 6704 18418 6760
rect 18474 6704 20730 6760
rect 18413 6702 20730 6704
rect 18413 6699 18479 6702
rect 20670 6626 20730 6702
rect 25497 6626 25563 6629
rect 20670 6624 25563 6626
rect 20670 6568 25502 6624
rect 25558 6568 25563 6624
rect 20670 6566 25563 6568
rect 25497 6563 25563 6566
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 200 6218 800 6248
rect 1761 6218 1827 6221
rect 200 6216 1827 6218
rect 200 6160 1766 6216
rect 1822 6160 1827 6216
rect 200 6158 1827 6160
rect 200 6128 800 6158
rect 1761 6155 1827 6158
rect 38285 6218 38351 6221
rect 39200 6218 39800 6248
rect 38285 6216 39800 6218
rect 38285 6160 38290 6216
rect 38346 6160 39800 6216
rect 38285 6158 39800 6160
rect 38285 6155 38351 6158
rect 39200 6128 39800 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 20989 5810 21055 5813
rect 21633 5810 21699 5813
rect 20989 5808 21699 5810
rect 20989 5752 20994 5808
rect 21050 5752 21638 5808
rect 21694 5752 21699 5808
rect 20989 5750 21699 5752
rect 20989 5747 21055 5750
rect 21633 5747 21699 5750
rect 5165 5674 5231 5677
rect 18137 5674 18203 5677
rect 18270 5674 18276 5676
rect 5165 5672 18276 5674
rect 5165 5616 5170 5672
rect 5226 5616 18142 5672
rect 18198 5616 18276 5672
rect 5165 5614 18276 5616
rect 5165 5611 5231 5614
rect 18137 5611 18203 5614
rect 18270 5612 18276 5614
rect 18340 5612 18346 5676
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 18321 5402 18387 5405
rect 18454 5402 18460 5404
rect 18321 5400 18460 5402
rect 18321 5344 18326 5400
rect 18382 5344 18460 5400
rect 18321 5342 18460 5344
rect 18321 5339 18387 5342
rect 18454 5340 18460 5342
rect 18524 5340 18530 5404
rect 13629 5266 13695 5269
rect 18597 5266 18663 5269
rect 13629 5264 18663 5266
rect 13629 5208 13634 5264
rect 13690 5208 18602 5264
rect 18658 5208 18663 5264
rect 13629 5206 18663 5208
rect 13629 5203 13695 5206
rect 18597 5203 18663 5206
rect 4210 4928 4526 4929
rect 200 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 1761 4858 1827 4861
rect 200 4856 1827 4858
rect 200 4800 1766 4856
rect 1822 4800 1827 4856
rect 200 4798 1827 4800
rect 200 4768 800 4798
rect 1761 4795 1827 4798
rect 5349 4858 5415 4861
rect 20713 4858 20779 4861
rect 5349 4856 20779 4858
rect 5349 4800 5354 4856
rect 5410 4800 20718 4856
rect 20774 4800 20779 4856
rect 5349 4798 20779 4800
rect 5349 4795 5415 4798
rect 20713 4795 20779 4798
rect 21449 4722 21515 4725
rect 25221 4722 25287 4725
rect 21449 4720 25287 4722
rect 21449 4664 21454 4720
rect 21510 4664 25226 4720
rect 25282 4664 25287 4720
rect 21449 4662 25287 4664
rect 21449 4659 21515 4662
rect 25221 4659 25287 4662
rect 11145 4586 11211 4589
rect 17677 4586 17743 4589
rect 11145 4584 17743 4586
rect 11145 4528 11150 4584
rect 11206 4528 17682 4584
rect 17738 4528 17743 4584
rect 11145 4526 17743 4528
rect 11145 4523 11211 4526
rect 17677 4523 17743 4526
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 13905 4178 13971 4181
rect 20805 4178 20871 4181
rect 13905 4176 20871 4178
rect 13905 4120 13910 4176
rect 13966 4120 20810 4176
rect 20866 4120 20871 4176
rect 13905 4118 20871 4120
rect 13905 4115 13971 4118
rect 20805 4115 20871 4118
rect 38193 4178 38259 4181
rect 39200 4178 39800 4208
rect 38193 4176 39800 4178
rect 38193 4120 38198 4176
rect 38254 4120 39800 4176
rect 38193 4118 39800 4120
rect 38193 4115 38259 4118
rect 39200 4088 39800 4118
rect 17677 4042 17743 4045
rect 21541 4042 21607 4045
rect 17677 4040 21607 4042
rect 17677 3984 17682 4040
rect 17738 3984 21546 4040
rect 21602 3984 21607 4040
rect 17677 3982 21607 3984
rect 17677 3979 17743 3982
rect 21541 3979 21607 3982
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 14365 3634 14431 3637
rect 17309 3634 17375 3637
rect 14365 3632 17375 3634
rect 14365 3576 14370 3632
rect 14426 3576 17314 3632
rect 17370 3576 17375 3632
rect 14365 3574 17375 3576
rect 14365 3571 14431 3574
rect 17309 3571 17375 3574
rect 20437 3634 20503 3637
rect 24209 3634 24275 3637
rect 20437 3632 24275 3634
rect 20437 3576 20442 3632
rect 20498 3576 24214 3632
rect 24270 3576 24275 3632
rect 20437 3574 24275 3576
rect 20437 3571 20503 3574
rect 24209 3571 24275 3574
rect 14641 3498 14707 3501
rect 21357 3498 21423 3501
rect 14641 3496 21423 3498
rect 14641 3440 14646 3496
rect 14702 3440 21362 3496
rect 21418 3440 21423 3496
rect 14641 3438 21423 3440
rect 14641 3435 14707 3438
rect 21357 3435 21423 3438
rect 14181 3362 14247 3365
rect 18965 3362 19031 3365
rect 14181 3360 19031 3362
rect 14181 3304 14186 3360
rect 14242 3304 18970 3360
rect 19026 3304 19031 3360
rect 14181 3302 19031 3304
rect 14181 3299 14247 3302
rect 18965 3299 19031 3302
rect 20345 3362 20411 3365
rect 24577 3362 24643 3365
rect 28717 3362 28783 3365
rect 20345 3360 28783 3362
rect 20345 3304 20350 3360
rect 20406 3304 24582 3360
rect 24638 3304 28722 3360
rect 28778 3304 28783 3360
rect 20345 3302 28783 3304
rect 20345 3299 20411 3302
rect 24577 3299 24643 3302
rect 28717 3299 28783 3302
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 3325 2954 3391 2957
rect 27337 2954 27403 2957
rect 3325 2952 27403 2954
rect 3325 2896 3330 2952
rect 3386 2896 27342 2952
rect 27398 2896 27403 2952
rect 3325 2894 27403 2896
rect 3325 2891 3391 2894
rect 27337 2891 27403 2894
rect 200 2818 800 2848
rect 1761 2818 1827 2821
rect 200 2816 1827 2818
rect 200 2760 1766 2816
rect 1822 2760 1827 2816
rect 200 2758 1827 2760
rect 200 2728 800 2758
rect 1761 2755 1827 2758
rect 38285 2818 38351 2821
rect 39200 2818 39800 2848
rect 38285 2816 39800 2818
rect 38285 2760 38290 2816
rect 38346 2760 39800 2816
rect 38285 2758 39800 2760
rect 38285 2755 38351 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 39200 2728 39800 2758
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 200 1458 800 1488
rect 2773 1458 2839 1461
rect 200 1456 2839 1458
rect 200 1400 2778 1456
rect 2834 1400 2839 1456
rect 200 1398 2839 1400
rect 200 1368 800 1398
rect 2773 1395 2839 1398
rect 38193 1458 38259 1461
rect 39200 1458 39800 1488
rect 38193 1456 39800 1458
rect 38193 1400 38198 1456
rect 38254 1400 39800 1456
rect 38193 1398 39800 1400
rect 38193 1395 38259 1398
rect 39200 1368 39800 1398
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 18276 24108 18340 24172
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 18460 11052 18524 11116
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 18460 7652 18524 7716
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 18276 5612 18340 5676
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 18460 5340 18524 5404
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 18275 24172 18341 24173
rect 18275 24108 18276 24172
rect 18340 24108 18341 24172
rect 18275 24107 18341 24108
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 18278 5677 18338 24107
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 18459 11116 18525 11117
rect 18459 11052 18460 11116
rect 18524 11052 18525 11116
rect 18459 11051 18525 11052
rect 18462 7717 18522 11051
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 18459 7716 18525 7717
rect 18459 7652 18460 7716
rect 18524 7652 18525 7716
rect 18459 7651 18525 7652
rect 18275 5676 18341 5677
rect 18275 5612 18276 5676
rect 18340 5612 18341 5676
rect 18275 5611 18341 5612
rect 18462 5405 18522 7651
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 18459 5404 18525 5405
rect 18459 5340 18460 5404
rect 18524 5340 18525 5404
rect 18459 5339 18525 5340
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6348 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1667941163
transform 1 0 11868 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2484 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1667941163
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1667941163
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63
timestamp 1667941163
transform 1 0 6900 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69
timestamp 1667941163
transform 1 0 7452 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 7820 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_91
timestamp 1667941163
transform 1 0 9476 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_99
timestamp 1667941163
transform 1 0 10212 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105
timestamp 1667941163
transform 1 0 10764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1667941163
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 11960 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_130
timestamp 1667941163
transform 1 0 13064 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1667941163
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1667941163
transform 1 0 14536 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1667941163
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1667941163
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_174
timestamp 1667941163
transform 1 0 17112 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_182
timestamp 1667941163
transform 1 0 17848 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_189
timestamp 1667941163
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1667941163
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_203
timestamp 1667941163
transform 1 0 19780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_210
timestamp 1667941163
transform 1 0 20424 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_218
timestamp 1667941163
transform 1 0 21160 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1667941163
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_233
timestamp 1667941163
transform 1 0 22540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_240
timestamp 1667941163
transform 1 0 23184 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_247
timestamp 1667941163
transform 1 0 23828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1667941163
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_259
timestamp 1667941163
transform 1 0 24932 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_267
timestamp 1667941163
transform 1 0 25668 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273
timestamp 1667941163
transform 1 0 26220 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1667941163
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_287
timestamp 1667941163
transform 1 0 27508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_294
timestamp 1667941163
transform 1 0 28152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1667941163
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1667941163
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_314
timestamp 1667941163
transform 1 0 29992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_321
timestamp 1667941163
transform 1 0 30636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_328
timestamp 1667941163
transform 1 0 31280 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_343
timestamp 1667941163
transform 1 0 32660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_350
timestamp 1667941163
transform 1 0 33304 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_357
timestamp 1667941163
transform 1 0 33948 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1667941163
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_370
timestamp 1667941163
transform 1 0 35144 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_378
timestamp 1667941163
transform 1 0 35880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_384
timestamp 1667941163
transform 1 0 36432 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_405
timestamp 1667941163
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1667941163
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_16
timestamp 1667941163
transform 1 0 2576 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_25
timestamp 1667941163
transform 1 0 3404 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1667941163
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_83
timestamp 1667941163
transform 1 0 8740 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1667941163
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_135
timestamp 1667941163
transform 1 0 13524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1667941163
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_181
timestamp 1667941163
transform 1 0 17756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_188
timestamp 1667941163
transform 1 0 18400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_192
timestamp 1667941163
transform 1 0 18768 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_214
timestamp 1667941163
transform 1 0 20792 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_218
timestamp 1667941163
transform 1 0 21160 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1667941163
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_236
timestamp 1667941163
transform 1 0 22816 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_243
timestamp 1667941163
transform 1 0 23460 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_247
timestamp 1667941163
transform 1 0 23828 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_256
timestamp 1667941163
transform 1 0 24656 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_263
timestamp 1667941163
transform 1 0 25300 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1667941163
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1667941163
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_291
timestamp 1667941163
transform 1 0 27876 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_308
timestamp 1667941163
transform 1 0 29440 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_321
timestamp 1667941163
transform 1 0 30636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_328
timestamp 1667941163
transform 1 0 31280 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_342
timestamp 1667941163
transform 1 0 32568 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_354
timestamp 1667941163
transform 1 0 33672 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_366
timestamp 1667941163
transform 1 0 34776 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_378
timestamp 1667941163
transform 1 0 35880 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_386
timestamp 1667941163
transform 1 0 36616 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1667941163
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_8
timestamp 1667941163
transform 1 0 1840 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1667941163
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_41
timestamp 1667941163
transform 1 0 4876 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_63
timestamp 1667941163
transform 1 0 6900 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_75
timestamp 1667941163
transform 1 0 8004 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1667941163
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1667941163
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1667941163
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1667941163
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1667941163
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_149
timestamp 1667941163
transform 1 0 14812 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_154
timestamp 1667941163
transform 1 0 15272 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_166
timestamp 1667941163
transform 1 0 16376 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_177
timestamp 1667941163
transform 1 0 17388 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_184
timestamp 1667941163
transform 1 0 18032 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_188
timestamp 1667941163
transform 1 0 18400 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1667941163
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_203
timestamp 1667941163
transform 1 0 19780 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_207
timestamp 1667941163
transform 1 0 20148 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_214
timestamp 1667941163
transform 1 0 20792 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_221
timestamp 1667941163
transform 1 0 21436 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_229
timestamp 1667941163
transform 1 0 22172 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_237
timestamp 1667941163
transform 1 0 22908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1667941163
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_258
timestamp 1667941163
transform 1 0 24840 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_264
timestamp 1667941163
transform 1 0 25392 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_273
timestamp 1667941163
transform 1 0 26220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_280
timestamp 1667941163
transform 1 0 26864 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_287
timestamp 1667941163
transform 1 0 27508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_294
timestamp 1667941163
transform 1 0 28152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1667941163
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1667941163
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_314
timestamp 1667941163
transform 1 0 29992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_318
timestamp 1667941163
transform 1 0 30360 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_327
timestamp 1667941163
transform 1 0 31188 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_334
timestamp 1667941163
transform 1 0 31832 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_341
timestamp 1667941163
transform 1 0 32476 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_353
timestamp 1667941163
transform 1 0 33580 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_361
timestamp 1667941163
transform 1 0 34316 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1667941163
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1667941163
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_401
timestamp 1667941163
transform 1 0 37996 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_405
timestamp 1667941163
transform 1 0 38364 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_8
timestamp 1667941163
transform 1 0 1840 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_20
timestamp 1667941163
transform 1 0 2944 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_32
timestamp 1667941163
transform 1 0 4048 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_44
timestamp 1667941163
transform 1 0 5152 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_69
timestamp 1667941163
transform 1 0 7452 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_77
timestamp 1667941163
transform 1 0 8188 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1667941163
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1667941163
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1667941163
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1667941163
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_125
timestamp 1667941163
transform 1 0 12604 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_147
timestamp 1667941163
transform 1 0 14628 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_159
timestamp 1667941163
transform 1 0 15732 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1667941163
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_174
timestamp 1667941163
transform 1 0 17112 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_180
timestamp 1667941163
transform 1 0 17664 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_202
timestamp 1667941163
transform 1 0 19688 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_209
timestamp 1667941163
transform 1 0 20332 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_217
timestamp 1667941163
transform 1 0 21068 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1667941163
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_230
timestamp 1667941163
transform 1 0 22264 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_237
timestamp 1667941163
transform 1 0 22908 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_244
timestamp 1667941163
transform 1 0 23552 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_252
timestamp 1667941163
transform 1 0 24288 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_257
timestamp 1667941163
transform 1 0 24748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_264
timestamp 1667941163
transform 1 0 25392 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_271
timestamp 1667941163
transform 1 0 26036 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1667941163
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_286
timestamp 1667941163
transform 1 0 27416 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_296
timestamp 1667941163
transform 1 0 28336 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_303
timestamp 1667941163
transform 1 0 28980 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_310
timestamp 1667941163
transform 1 0 29624 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_314
timestamp 1667941163
transform 1 0 29992 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_318
timestamp 1667941163
transform 1 0 30360 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_325
timestamp 1667941163
transform 1 0 31004 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_333
timestamp 1667941163
transform 1 0 31740 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1667941163
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1667941163
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1667941163
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1667941163
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1667941163
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1667941163
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_54
timestamp 1667941163
transform 1 0 6072 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_66
timestamp 1667941163
transform 1 0 7176 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_78
timestamp 1667941163
transform 1 0 8280 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_97
timestamp 1667941163
transform 1 0 10028 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_101
timestamp 1667941163
transform 1 0 10396 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_122
timestamp 1667941163
transform 1 0 12328 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_134
timestamp 1667941163
transform 1 0 13432 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_163
timestamp 1667941163
transform 1 0 16100 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_174
timestamp 1667941163
transform 1 0 17112 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_181
timestamp 1667941163
transform 1 0 17756 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_188
timestamp 1667941163
transform 1 0 18400 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_209
timestamp 1667941163
transform 1 0 20332 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_213
timestamp 1667941163
transform 1 0 20700 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1667941163
transform 1 0 21252 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_223
timestamp 1667941163
transform 1 0 21620 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_230
timestamp 1667941163
transform 1 0 22264 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1667941163
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_258
timestamp 1667941163
transform 1 0 24840 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_270
timestamp 1667941163
transform 1 0 25944 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_277
timestamp 1667941163
transform 1 0 26588 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_283
timestamp 1667941163
transform 1 0 27140 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_287
timestamp 1667941163
transform 1 0 27508 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_299
timestamp 1667941163
transform 1 0 28612 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_306
timestamp 1667941163
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1667941163
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1667941163
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1667941163
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1667941163
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1667941163
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_405
timestamp 1667941163
transform 1 0 38364 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_9
timestamp 1667941163
transform 1 0 1932 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_16
timestamp 1667941163
transform 1 0 2576 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_49
timestamp 1667941163
transform 1 0 5612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1667941163
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1667941163
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_81
timestamp 1667941163
transform 1 0 8556 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_87
timestamp 1667941163
transform 1 0 9108 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1667941163
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1667941163
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_137
timestamp 1667941163
transform 1 0 13708 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_160
timestamp 1667941163
transform 1 0 15824 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_175
timestamp 1667941163
transform 1 0 17204 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_204
timestamp 1667941163
transform 1 0 19872 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_216
timestamp 1667941163
transform 1 0 20976 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1667941163
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_231
timestamp 1667941163
transform 1 0 22356 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_239
timestamp 1667941163
transform 1 0 23092 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_244
timestamp 1667941163
transform 1 0 23552 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_251
timestamp 1667941163
transform 1 0 24196 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_258
timestamp 1667941163
transform 1 0 24840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_265
timestamp 1667941163
transform 1 0 25484 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_272
timestamp 1667941163
transform 1 0 26128 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_286
timestamp 1667941163
transform 1 0 27416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_293
timestamp 1667941163
transform 1 0 28060 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_300
timestamp 1667941163
transform 1 0 28704 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_308
timestamp 1667941163
transform 1 0 29440 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_314
timestamp 1667941163
transform 1 0 29992 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_321
timestamp 1667941163
transform 1 0 30636 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_328
timestamp 1667941163
transform 1 0 31280 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1667941163
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1667941163
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1667941163
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1667941163
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1667941163
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1667941163
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_8
timestamp 1667941163
transform 1 0 1840 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_20
timestamp 1667941163
transform 1 0 2944 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_52
timestamp 1667941163
transform 1 0 5888 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_64
timestamp 1667941163
transform 1 0 6992 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_76
timestamp 1667941163
transform 1 0 8096 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1667941163
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_109
timestamp 1667941163
transform 1 0 11132 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1667941163
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1667941163
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_153
timestamp 1667941163
transform 1 0 15180 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_161
timestamp 1667941163
transform 1 0 15916 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_186
timestamp 1667941163
transform 1 0 18216 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1667941163
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_209
timestamp 1667941163
transform 1 0 20332 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_213
timestamp 1667941163
transform 1 0 20700 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_223
timestamp 1667941163
transform 1 0 21620 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_230
timestamp 1667941163
transform 1 0 22264 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_237
timestamp 1667941163
transform 1 0 22908 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_244
timestamp 1667941163
transform 1 0 23552 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_258
timestamp 1667941163
transform 1 0 24840 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_265
timestamp 1667941163
transform 1 0 25484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_269
timestamp 1667941163
transform 1 0 25852 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_273
timestamp 1667941163
transform 1 0 26220 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_285
timestamp 1667941163
transform 1 0 27324 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_290
timestamp 1667941163
transform 1 0 27784 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_297
timestamp 1667941163
transform 1 0 28428 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_304
timestamp 1667941163
transform 1 0 29072 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_313
timestamp 1667941163
transform 1 0 29900 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_317
timestamp 1667941163
transform 1 0 30268 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_326
timestamp 1667941163
transform 1 0 31096 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_338
timestamp 1667941163
transform 1 0 32200 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_350
timestamp 1667941163
transform 1 0 33304 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_362
timestamp 1667941163
transform 1 0 34408 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1667941163
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1667941163
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_401
timestamp 1667941163
transform 1 0 37996 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7
timestamp 1667941163
transform 1 0 1748 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_12
timestamp 1667941163
transform 1 0 2208 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_24
timestamp 1667941163
transform 1 0 3312 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_30
timestamp 1667941163
transform 1 0 3864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1667941163
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1667941163
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_81
timestamp 1667941163
transform 1 0 8556 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_103
timestamp 1667941163
transform 1 0 10580 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1667941163
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1667941163
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1667941163
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1667941163
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1667941163
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1667941163
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_181
timestamp 1667941163
transform 1 0 17756 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_191
timestamp 1667941163
transform 1 0 18676 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_198
timestamp 1667941163
transform 1 0 19320 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_207
timestamp 1667941163
transform 1 0 20148 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_215
timestamp 1667941163
transform 1 0 20884 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_219
timestamp 1667941163
transform 1 0 21252 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1667941163
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_230
timestamp 1667941163
transform 1 0 22264 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_247
timestamp 1667941163
transform 1 0 23828 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_254
timestamp 1667941163
transform 1 0 24472 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_260
timestamp 1667941163
transform 1 0 25024 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_270
timestamp 1667941163
transform 1 0 25944 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp 1667941163
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_292
timestamp 1667941163
transform 1 0 27968 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_305
timestamp 1667941163
transform 1 0 29164 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_313
timestamp 1667941163
transform 1 0 29900 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_317
timestamp 1667941163
transform 1 0 30268 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1667941163
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1667941163
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1667941163
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1667941163
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1667941163
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1667941163
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1667941163
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_401
timestamp 1667941163
transform 1 0 37996 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_9
timestamp 1667941163
transform 1 0 1932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_14
timestamp 1667941163
transform 1 0 2392 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_21
timestamp 1667941163
transform 1 0 3036 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1667941163
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1667941163
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_53
timestamp 1667941163
transform 1 0 5980 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_75
timestamp 1667941163
transform 1 0 8004 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1667941163
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_93
timestamp 1667941163
transform 1 0 9660 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_116
timestamp 1667941163
transform 1 0 11776 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_128
timestamp 1667941163
transform 1 0 12880 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1667941163
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1667941163
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1667941163
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1667941163
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1667941163
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_209
timestamp 1667941163
transform 1 0 20332 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1667941163
transform 1 0 20700 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_217
timestamp 1667941163
transform 1 0 21068 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_224
timestamp 1667941163
transform 1 0 21712 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_230
timestamp 1667941163
transform 1 0 22264 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_239
timestamp 1667941163
transform 1 0 23092 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_246
timestamp 1667941163
transform 1 0 23736 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1667941163
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1667941163
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_289
timestamp 1667941163
transform 1 0 27692 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_297
timestamp 1667941163
transform 1 0 28428 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_303
timestamp 1667941163
transform 1 0 28980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1667941163
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1667941163
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1667941163
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1667941163
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1667941163
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1667941163
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1667941163
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_401
timestamp 1667941163
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_12
timestamp 1667941163
transform 1 0 2208 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_24
timestamp 1667941163
transform 1 0 3312 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_36
timestamp 1667941163
transform 1 0 4416 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_48
timestamp 1667941163
transform 1 0 5520 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_69
timestamp 1667941163
transform 1 0 7452 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_90
timestamp 1667941163
transform 1 0 9384 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_102
timestamp 1667941163
transform 1 0 10488 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1667941163
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1667941163
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_137
timestamp 1667941163
transform 1 0 13708 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1667941163
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1667941163
transform 1 0 17756 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_206
timestamp 1667941163
transform 1 0 20056 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_218
timestamp 1667941163
transform 1 0 21160 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1667941163
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_230
timestamp 1667941163
transform 1 0 22264 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_237
timestamp 1667941163
transform 1 0 22908 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_246
timestamp 1667941163
transform 1 0 23736 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_254
timestamp 1667941163
transform 1 0 24472 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_265
timestamp 1667941163
transform 1 0 25484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp 1667941163
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_286
timestamp 1667941163
transform 1 0 27416 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_298
timestamp 1667941163
transform 1 0 28520 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_302
timestamp 1667941163
transform 1 0 28888 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_312
timestamp 1667941163
transform 1 0 29808 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_319
timestamp 1667941163
transform 1 0 30452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_331
timestamp 1667941163
transform 1 0 31556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1667941163
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1667941163
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1667941163
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1667941163
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1667941163
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_12
timestamp 1667941163
transform 1 0 2208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_19
timestamp 1667941163
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1667941163
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_51
timestamp 1667941163
transform 1 0 5796 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1667941163
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1667941163
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_130
timestamp 1667941163
transform 1 0 13064 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1667941163
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_164
timestamp 1667941163
transform 1 0 16192 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_176
timestamp 1667941163
transform 1 0 17296 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_188
timestamp 1667941163
transform 1 0 18400 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1667941163
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_220
timestamp 1667941163
transform 1 0 21344 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_227
timestamp 1667941163
transform 1 0 21988 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_234
timestamp 1667941163
transform 1 0 22632 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_246
timestamp 1667941163
transform 1 0 23736 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1667941163
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_258
timestamp 1667941163
transform 1 0 24840 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_265
timestamp 1667941163
transform 1 0 25484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_272
timestamp 1667941163
transform 1 0 26128 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_281
timestamp 1667941163
transform 1 0 26956 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_293
timestamp 1667941163
transform 1 0 28060 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_304
timestamp 1667941163
transform 1 0 29072 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_314
timestamp 1667941163
transform 1 0 29992 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_321
timestamp 1667941163
transform 1 0 30636 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_329
timestamp 1667941163
transform 1 0 31372 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_335
timestamp 1667941163
transform 1 0 31924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_347
timestamp 1667941163
transform 1 0 33028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_359
timestamp 1667941163
transform 1 0 34132 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1667941163
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1667941163
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_401
timestamp 1667941163
transform 1 0 37996 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_405
timestamp 1667941163
transform 1 0 38364 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_12
timestamp 1667941163
transform 1 0 2208 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_24
timestamp 1667941163
transform 1 0 3312 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1667941163
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1667941163
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_69
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_98
timestamp 1667941163
transform 1 0 10120 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1667941163
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1667941163
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1667941163
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_149
timestamp 1667941163
transform 1 0 14812 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_154
timestamp 1667941163
transform 1 0 15272 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1667941163
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_181
timestamp 1667941163
transform 1 0 17756 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_205
timestamp 1667941163
transform 1 0 19964 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_213
timestamp 1667941163
transform 1 0 20700 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_219
timestamp 1667941163
transform 1 0 21252 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1667941163
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_240
timestamp 1667941163
transform 1 0 23184 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_247
timestamp 1667941163
transform 1 0 23828 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_255
timestamp 1667941163
transform 1 0 24564 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_264
timestamp 1667941163
transform 1 0 25392 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_268
timestamp 1667941163
transform 1 0 25760 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp 1667941163
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_291
timestamp 1667941163
transform 1 0 27876 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_298
timestamp 1667941163
transform 1 0 28520 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_305
timestamp 1667941163
transform 1 0 29164 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_312
timestamp 1667941163
transform 1 0 29808 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_327
timestamp 1667941163
transform 1 0 31188 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1667941163
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_342
timestamp 1667941163
transform 1 0 32568 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_354
timestamp 1667941163
transform 1 0 33672 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_366
timestamp 1667941163
transform 1 0 34776 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_378
timestamp 1667941163
transform 1 0 35880 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_390
timestamp 1667941163
transform 1 0 36984 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_7
timestamp 1667941163
transform 1 0 1748 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_11
timestamp 1667941163
transform 1 0 2116 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_23
timestamp 1667941163
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1667941163
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_41
timestamp 1667941163
transform 1 0 4876 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_49
timestamp 1667941163
transform 1 0 5612 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_61
timestamp 1667941163
transform 1 0 6716 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_73
timestamp 1667941163
transform 1 0 7820 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_81
timestamp 1667941163
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1667941163
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_109
timestamp 1667941163
transform 1 0 11132 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_114
timestamp 1667941163
transform 1 0 11592 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1667941163
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1667941163
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1667941163
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1667941163
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_165
timestamp 1667941163
transform 1 0 16284 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_191
timestamp 1667941163
transform 1 0 18676 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1667941163
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_209
timestamp 1667941163
transform 1 0 20332 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_214
timestamp 1667941163
transform 1 0 20792 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_222
timestamp 1667941163
transform 1 0 21528 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_226
timestamp 1667941163
transform 1 0 21896 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_232
timestamp 1667941163
transform 1 0 22448 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_239
timestamp 1667941163
transform 1 0 23092 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_246
timestamp 1667941163
transform 1 0 23736 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_264
timestamp 1667941163
transform 1 0 25392 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_271
timestamp 1667941163
transform 1 0 26036 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_275
timestamp 1667941163
transform 1 0 26404 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_279
timestamp 1667941163
transform 1 0 26772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_291
timestamp 1667941163
transform 1 0 27876 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_295
timestamp 1667941163
transform 1 0 28244 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_302
timestamp 1667941163
transform 1 0 28888 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_317
timestamp 1667941163
transform 1 0 30268 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_323
timestamp 1667941163
transform 1 0 30820 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_335
timestamp 1667941163
transform 1 0 31924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_347
timestamp 1667941163
transform 1 0 33028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_359
timestamp 1667941163
transform 1 0 34132 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1667941163
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1667941163
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_405
timestamp 1667941163
transform 1 0 38364 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1667941163
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1667941163
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1667941163
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1667941163
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1667941163
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_82
timestamp 1667941163
transform 1 0 8648 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_86
timestamp 1667941163
transform 1 0 9016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1667941163
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1667941163
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_137
timestamp 1667941163
transform 1 0 13708 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1667941163
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1667941163
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_181
timestamp 1667941163
transform 1 0 17756 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_185
timestamp 1667941163
transform 1 0 18124 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_207
timestamp 1667941163
transform 1 0 20148 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_214
timestamp 1667941163
transform 1 0 20792 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_221
timestamp 1667941163
transform 1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_231
timestamp 1667941163
transform 1 0 22356 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_238
timestamp 1667941163
transform 1 0 23000 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_247
timestamp 1667941163
transform 1 0 23828 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_259
timestamp 1667941163
transform 1 0 24932 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_271
timestamp 1667941163
transform 1 0 26036 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1667941163
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_293
timestamp 1667941163
transform 1 0 28060 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_307
timestamp 1667941163
transform 1 0 29348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_319
timestamp 1667941163
transform 1 0 30452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_331
timestamp 1667941163
transform 1 0 31556 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1667941163
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1667941163
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1667941163
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1667941163
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1667941163
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_8
timestamp 1667941163
transform 1 0 1840 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_20
timestamp 1667941163
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_54
timestamp 1667941163
transform 1 0 6072 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_67
timestamp 1667941163
transform 1 0 7268 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_79
timestamp 1667941163
transform 1 0 8372 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1667941163
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1667941163
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1667941163
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1667941163
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1667941163
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1667941163
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1667941163
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1667941163
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1667941163
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1667941163
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1667941163
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_209
timestamp 1667941163
transform 1 0 20332 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_213
timestamp 1667941163
transform 1 0 20700 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1667941163
transform 1 0 21252 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_223
timestamp 1667941163
transform 1 0 21620 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_230
timestamp 1667941163
transform 1 0 22264 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_237
timestamp 1667941163
transform 1 0 22908 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_246
timestamp 1667941163
transform 1 0 23736 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_268
timestamp 1667941163
transform 1 0 25760 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_280
timestamp 1667941163
transform 1 0 26864 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_292
timestamp 1667941163
transform 1 0 27968 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_304
timestamp 1667941163
transform 1 0 29072 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_315
timestamp 1667941163
transform 1 0 30084 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_327
timestamp 1667941163
transform 1 0 31188 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_339
timestamp 1667941163
transform 1 0 32292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_351
timestamp 1667941163
transform 1 0 33396 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1667941163
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1667941163
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_401
timestamp 1667941163
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_7
timestamp 1667941163
transform 1 0 1748 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_11
timestamp 1667941163
transform 1 0 2116 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_23
timestamp 1667941163
transform 1 0 3220 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_35
timestamp 1667941163
transform 1 0 4324 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_43
timestamp 1667941163
transform 1 0 5060 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1667941163
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_73
timestamp 1667941163
transform 1 0 7820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_85
timestamp 1667941163
transform 1 0 8924 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_97
timestamp 1667941163
transform 1 0 10028 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_101
timestamp 1667941163
transform 1 0 10396 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1667941163
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1667941163
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_145
timestamp 1667941163
transform 1 0 14444 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_157
timestamp 1667941163
transform 1 0 15548 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_165
timestamp 1667941163
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_192
timestamp 1667941163
transform 1 0 18768 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_204
timestamp 1667941163
transform 1 0 19872 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_212
timestamp 1667941163
transform 1 0 20608 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_220
timestamp 1667941163
transform 1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_233
timestamp 1667941163
transform 1 0 22540 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_241
timestamp 1667941163
transform 1 0 23276 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_252
timestamp 1667941163
transform 1 0 24288 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_263
timestamp 1667941163
transform 1 0 25300 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_275
timestamp 1667941163
transform 1 0 26404 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1667941163
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_293
timestamp 1667941163
transform 1 0 28060 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_297
timestamp 1667941163
transform 1 0 28428 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_301
timestamp 1667941163
transform 1 0 28796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_308
timestamp 1667941163
transform 1 0 29440 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_320
timestamp 1667941163
transform 1 0 30544 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_332
timestamp 1667941163
transform 1 0 31648 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_358
timestamp 1667941163
transform 1 0 34040 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_370
timestamp 1667941163
transform 1 0 35144 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_382
timestamp 1667941163
transform 1 0 36248 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_390
timestamp 1667941163
transform 1 0 36984 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_8
timestamp 1667941163
transform 1 0 1840 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_20
timestamp 1667941163
transform 1 0 2944 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_55
timestamp 1667941163
transform 1 0 6164 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_59
timestamp 1667941163
transform 1 0 6532 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1667941163
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1667941163
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1667941163
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1667941163
transform 1 0 9476 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_113
timestamp 1667941163
transform 1 0 11500 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_125
timestamp 1667941163
transform 1 0 12604 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_137
timestamp 1667941163
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1667941163
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_165
timestamp 1667941163
transform 1 0 16284 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_173
timestamp 1667941163
transform 1 0 17020 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1667941163
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1667941163
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_221
timestamp 1667941163
transform 1 0 21436 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_228
timestamp 1667941163
transform 1 0 22080 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_236
timestamp 1667941163
transform 1 0 22816 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_242
timestamp 1667941163
transform 1 0 23368 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_249
timestamp 1667941163
transform 1 0 24012 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_263
timestamp 1667941163
transform 1 0 25300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_275
timestamp 1667941163
transform 1 0 26404 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_280
timestamp 1667941163
transform 1 0 26864 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_295
timestamp 1667941163
transform 1 0 28244 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_301
timestamp 1667941163
transform 1 0 28796 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_305
timestamp 1667941163
transform 1 0 29164 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_321
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_332
timestamp 1667941163
transform 1 0 31648 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_344
timestamp 1667941163
transform 1 0 32752 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_356
timestamp 1667941163
transform 1 0 33856 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1667941163
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_401
timestamp 1667941163
transform 1 0 37996 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_405
timestamp 1667941163
transform 1 0 38364 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1667941163
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_27
timestamp 1667941163
transform 1 0 3588 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_33
timestamp 1667941163
transform 1 0 4140 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1667941163
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_65
timestamp 1667941163
transform 1 0 7084 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_89
timestamp 1667941163
transform 1 0 9292 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_101
timestamp 1667941163
transform 1 0 10396 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_109
timestamp 1667941163
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_136
timestamp 1667941163
transform 1 0 13616 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_144
timestamp 1667941163
transform 1 0 14352 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1667941163
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_181
timestamp 1667941163
transform 1 0 17756 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_185
timestamp 1667941163
transform 1 0 18124 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_209
timestamp 1667941163
transform 1 0 20332 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_217
timestamp 1667941163
transform 1 0 21068 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1667941163
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1667941163
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1667941163
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_264
timestamp 1667941163
transform 1 0 25392 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_276
timestamp 1667941163
transform 1 0 26496 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_293
timestamp 1667941163
transform 1 0 28060 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_301
timestamp 1667941163
transform 1 0 28796 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_312
timestamp 1667941163
transform 1 0 29808 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_324
timestamp 1667941163
transform 1 0 30912 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_348
timestamp 1667941163
transform 1 0 33120 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_360
timestamp 1667941163
transform 1 0 34224 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_372
timestamp 1667941163
transform 1 0 35328 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_384
timestamp 1667941163
transform 1 0 36432 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_7
timestamp 1667941163
transform 1 0 1748 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_11
timestamp 1667941163
transform 1 0 2116 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_23
timestamp 1667941163
transform 1 0 3220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1667941163
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_54
timestamp 1667941163
transform 1 0 6072 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_66
timestamp 1667941163
transform 1 0 7176 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_78
timestamp 1667941163
transform 1 0 8280 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1667941163
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_109
timestamp 1667941163
transform 1 0 11132 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_124
timestamp 1667941163
transform 1 0 12512 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1667941163
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_146
timestamp 1667941163
transform 1 0 14536 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_158
timestamp 1667941163
transform 1 0 15640 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_170
timestamp 1667941163
transform 1 0 16744 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_182
timestamp 1667941163
transform 1 0 17848 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1667941163
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1667941163
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_221
timestamp 1667941163
transform 1 0 21436 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_225
timestamp 1667941163
transform 1 0 21804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_229
timestamp 1667941163
transform 1 0 22172 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_239
timestamp 1667941163
transform 1 0 23092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1667941163
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_257
timestamp 1667941163
transform 1 0 24748 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_261
timestamp 1667941163
transform 1 0 25116 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_269
timestamp 1667941163
transform 1 0 25852 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_278
timestamp 1667941163
transform 1 0 26680 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_286
timestamp 1667941163
transform 1 0 27416 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_297
timestamp 1667941163
transform 1 0 28428 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_304
timestamp 1667941163
transform 1 0 29072 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_320
timestamp 1667941163
transform 1 0 30544 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_327
timestamp 1667941163
transform 1 0 31188 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_331
timestamp 1667941163
transform 1 0 31556 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_335
timestamp 1667941163
transform 1 0 31924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_342
timestamp 1667941163
transform 1 0 32568 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_353
timestamp 1667941163
transform 1 0 33580 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_361
timestamp 1667941163
transform 1 0 34316 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_380
timestamp 1667941163
transform 1 0 36064 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_392
timestamp 1667941163
transform 1 0 37168 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_404
timestamp 1667941163
transform 1 0 38272 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_8
timestamp 1667941163
transform 1 0 1840 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_20
timestamp 1667941163
transform 1 0 2944 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_32
timestamp 1667941163
transform 1 0 4048 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_44
timestamp 1667941163
transform 1 0 5152 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1667941163
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_81
timestamp 1667941163
transform 1 0 8556 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1667941163
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1667941163
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_119
timestamp 1667941163
transform 1 0 12052 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_144
timestamp 1667941163
transform 1 0 14352 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_156
timestamp 1667941163
transform 1 0 15456 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_197
timestamp 1667941163
transform 1 0 19228 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_209
timestamp 1667941163
transform 1 0 20332 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_220
timestamp 1667941163
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_230
timestamp 1667941163
transform 1 0 22264 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_242
timestamp 1667941163
transform 1 0 23368 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_251
timestamp 1667941163
transform 1 0 24196 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_263
timestamp 1667941163
transform 1 0 25300 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_275
timestamp 1667941163
transform 1 0 26404 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1667941163
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_289
timestamp 1667941163
transform 1 0 27692 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_293
timestamp 1667941163
transform 1 0 28060 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_300
timestamp 1667941163
transform 1 0 28704 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_312
timestamp 1667941163
transform 1 0 29808 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_320
timestamp 1667941163
transform 1 0 30544 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_331
timestamp 1667941163
transform 1 0 31556 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1667941163
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1667941163
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1667941163
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1667941163
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1667941163
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1667941163
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_7
timestamp 1667941163
transform 1 0 1748 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_11
timestamp 1667941163
transform 1 0 2116 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_23
timestamp 1667941163
transform 1 0 3220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1667941163
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_51
timestamp 1667941163
transform 1 0 5796 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_63
timestamp 1667941163
transform 1 0 6900 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_75
timestamp 1667941163
transform 1 0 8004 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1667941163
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_90
timestamp 1667941163
transform 1 0 9384 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_102
timestamp 1667941163
transform 1 0 10488 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_129
timestamp 1667941163
transform 1 0 12972 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_137
timestamp 1667941163
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_164
timestamp 1667941163
transform 1 0 16192 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_176
timestamp 1667941163
transform 1 0 17296 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_188
timestamp 1667941163
transform 1 0 18400 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_209
timestamp 1667941163
transform 1 0 20332 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_220
timestamp 1667941163
transform 1 0 21344 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_227
timestamp 1667941163
transform 1 0 21988 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_234
timestamp 1667941163
transform 1 0 22632 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_246
timestamp 1667941163
transform 1 0 23736 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_264
timestamp 1667941163
transform 1 0 25392 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_280
timestamp 1667941163
transform 1 0 26864 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_292
timestamp 1667941163
transform 1 0 27968 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_303
timestamp 1667941163
transform 1 0 28980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1667941163
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_314
timestamp 1667941163
transform 1 0 29992 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_318
timestamp 1667941163
transform 1 0 30360 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_328
timestamp 1667941163
transform 1 0 31280 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_334
timestamp 1667941163
transform 1 0 31832 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_338
timestamp 1667941163
transform 1 0 32200 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_350
timestamp 1667941163
transform 1 0 33304 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_362
timestamp 1667941163
transform 1 0 34408 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_401
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_10
timestamp 1667941163
transform 1 0 2024 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_17
timestamp 1667941163
transform 1 0 2668 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_25
timestamp 1667941163
transform 1 0 3404 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_49
timestamp 1667941163
transform 1 0 5612 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1667941163
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_69
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_94
timestamp 1667941163
transform 1 0 9752 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_106
timestamp 1667941163
transform 1 0 10856 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_125
timestamp 1667941163
transform 1 0 12604 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_133
timestamp 1667941163
transform 1 0 13340 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_155
timestamp 1667941163
transform 1 0 15364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1667941163
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_181
timestamp 1667941163
transform 1 0 17756 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_210
timestamp 1667941163
transform 1 0 20424 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_221
timestamp 1667941163
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_230
timestamp 1667941163
transform 1 0 22264 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_237
timestamp 1667941163
transform 1 0 22908 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_245
timestamp 1667941163
transform 1 0 23644 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_255
timestamp 1667941163
transform 1 0 24564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_259
timestamp 1667941163
transform 1 0 24932 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_268
timestamp 1667941163
transform 1 0 25760 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_291
timestamp 1667941163
transform 1 0 27876 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_304
timestamp 1667941163
transform 1 0 29072 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_316
timestamp 1667941163
transform 1 0 30176 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_327
timestamp 1667941163
transform 1 0 31188 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1667941163
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1667941163
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1667941163
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1667941163
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_10
timestamp 1667941163
transform 1 0 2024 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_22
timestamp 1667941163
transform 1 0 3128 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1667941163
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1667941163
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1667941163
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1667941163
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1667941163
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_97
timestamp 1667941163
transform 1 0 10028 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_105
timestamp 1667941163
transform 1 0 10764 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_110
timestamp 1667941163
transform 1 0 11224 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_122
timestamp 1667941163
transform 1 0 12328 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_134
timestamp 1667941163
transform 1 0 13432 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_153
timestamp 1667941163
transform 1 0 15180 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_159
timestamp 1667941163
transform 1 0 15732 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_180
timestamp 1667941163
transform 1 0 17664 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1667941163
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_209
timestamp 1667941163
transform 1 0 20332 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_220
timestamp 1667941163
transform 1 0 21344 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_228
timestamp 1667941163
transform 1 0 22080 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_232
timestamp 1667941163
transform 1 0 22448 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_244
timestamp 1667941163
transform 1 0 23552 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_261
timestamp 1667941163
transform 1 0 25116 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1667941163
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_277
timestamp 1667941163
transform 1 0 26588 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_282
timestamp 1667941163
transform 1 0 27048 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_294
timestamp 1667941163
transform 1 0 28152 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_298
timestamp 1667941163
transform 1 0 28520 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1667941163
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_321
timestamp 1667941163
transform 1 0 30636 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_336
timestamp 1667941163
transform 1 0 32016 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_348
timestamp 1667941163
transform 1 0 33120 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_360
timestamp 1667941163
transform 1 0 34224 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1667941163
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1667941163
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_401
timestamp 1667941163
transform 1 0 37996 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_405
timestamp 1667941163
transform 1 0 38364 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_8
timestamp 1667941163
transform 1 0 1840 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_20
timestamp 1667941163
transform 1 0 2944 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_26
timestamp 1667941163
transform 1 0 3496 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_48
timestamp 1667941163
transform 1 0 5520 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1667941163
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_81
timestamp 1667941163
transform 1 0 8556 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_104
timestamp 1667941163
transform 1 0 10672 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_119
timestamp 1667941163
transform 1 0 12052 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_141
timestamp 1667941163
transform 1 0 14076 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1667941163
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_181
timestamp 1667941163
transform 1 0 17756 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_208
timestamp 1667941163
transform 1 0 20240 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1667941163
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_229
timestamp 1667941163
transform 1 0 22172 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_233
timestamp 1667941163
transform 1 0 22540 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_240
timestamp 1667941163
transform 1 0 23184 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_247
timestamp 1667941163
transform 1 0 23828 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_259
timestamp 1667941163
transform 1 0 24932 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_274
timestamp 1667941163
transform 1 0 26312 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_286
timestamp 1667941163
transform 1 0 27416 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_292
timestamp 1667941163
transform 1 0 27968 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_302
timestamp 1667941163
transform 1 0 28888 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_309
timestamp 1667941163
transform 1 0 29532 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_321
timestamp 1667941163
transform 1 0 30636 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_333
timestamp 1667941163
transform 1 0 31740 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1667941163
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1667941163
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1667941163
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1667941163
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1667941163
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1667941163
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1667941163
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_57
timestamp 1667941163
transform 1 0 6348 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1667941163
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_107
timestamp 1667941163
transform 1 0 10948 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_134
timestamp 1667941163
transform 1 0 13432 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_153
timestamp 1667941163
transform 1 0 15180 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1667941163
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1667941163
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_212
timestamp 1667941163
transform 1 0 20608 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_221
timestamp 1667941163
transform 1 0 21436 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_228
timestamp 1667941163
transform 1 0 22080 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_232
timestamp 1667941163
transform 1 0 22448 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_236
timestamp 1667941163
transform 1 0 22816 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_240
timestamp 1667941163
transform 1 0 23184 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1667941163
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_257
timestamp 1667941163
transform 1 0 24748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_261
timestamp 1667941163
transform 1 0 25116 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_268
timestamp 1667941163
transform 1 0 25760 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_280
timestamp 1667941163
transform 1 0 26864 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_284
timestamp 1667941163
transform 1 0 27232 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_288
timestamp 1667941163
transform 1 0 27600 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_297
timestamp 1667941163
transform 1 0 28428 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_304
timestamp 1667941163
transform 1 0 29072 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_321
timestamp 1667941163
transform 1 0 30636 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_332
timestamp 1667941163
transform 1 0 31648 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_347
timestamp 1667941163
transform 1 0 33028 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_354
timestamp 1667941163
transform 1 0 33672 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_362
timestamp 1667941163
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1667941163
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_401
timestamp 1667941163
transform 1 0 37996 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_9
timestamp 1667941163
transform 1 0 1932 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_17
timestamp 1667941163
transform 1 0 2668 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_21
timestamp 1667941163
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_33
timestamp 1667941163
transform 1 0 4140 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_25_42
timestamp 1667941163
transform 1 0 4968 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1667941163
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1667941163
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1667941163
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1667941163
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_93
timestamp 1667941163
transform 1 0 9660 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1667941163
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1667941163
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1667941163
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1667941163
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1667941163
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1667941163
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_181
timestamp 1667941163
transform 1 0 17756 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_187
timestamp 1667941163
transform 1 0 18308 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_209
timestamp 1667941163
transform 1 0 20332 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_25_218
timestamp 1667941163
transform 1 0 21160 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_231
timestamp 1667941163
transform 1 0 22356 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_235
timestamp 1667941163
transform 1 0 22724 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_244
timestamp 1667941163
transform 1 0 23552 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_251
timestamp 1667941163
transform 1 0 24196 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_263
timestamp 1667941163
transform 1 0 25300 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1667941163
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1667941163
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_286
timestamp 1667941163
transform 1 0 27416 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_294
timestamp 1667941163
transform 1 0 28152 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_305
timestamp 1667941163
transform 1 0 29164 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_312
timestamp 1667941163
transform 1 0 29808 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_324
timestamp 1667941163
transform 1 0 30912 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_331
timestamp 1667941163
transform 1 0 31556 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1667941163
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1667941163
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1667941163
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1667941163
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1667941163
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1667941163
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_11
timestamp 1667941163
transform 1 0 2116 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_16
timestamp 1667941163
transform 1 0 2576 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_22
timestamp 1667941163
transform 1 0 3128 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1667941163
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_35
timestamp 1667941163
transform 1 0 4324 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_42
timestamp 1667941163
transform 1 0 4968 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_49
timestamp 1667941163
transform 1 0 5612 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_57
timestamp 1667941163
transform 1 0 6348 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_62
timestamp 1667941163
transform 1 0 6808 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_69
timestamp 1667941163
transform 1 0 7452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_81
timestamp 1667941163
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_90
timestamp 1667941163
transform 1 0 9384 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_102
timestamp 1667941163
transform 1 0 10488 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_114
timestamp 1667941163
transform 1 0 11592 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_118
timestamp 1667941163
transform 1 0 11960 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_122
timestamp 1667941163
transform 1 0 12328 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_134
timestamp 1667941163
transform 1 0 13432 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1667941163
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1667941163
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_177
timestamp 1667941163
transform 1 0 17388 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_181
timestamp 1667941163
transform 1 0 17756 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_185
timestamp 1667941163
transform 1 0 18124 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1667941163
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1667941163
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1667941163
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1667941163
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_248
timestamp 1667941163
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_265
timestamp 1667941163
transform 1 0 25484 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_271
timestamp 1667941163
transform 1 0 26036 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_283
timestamp 1667941163
transform 1 0 27140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_295
timestamp 1667941163
transform 1 0 28244 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1667941163
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_315
timestamp 1667941163
transform 1 0 30084 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_324
timestamp 1667941163
transform 1 0 30912 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_336
timestamp 1667941163
transform 1 0 32016 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_343
timestamp 1667941163
transform 1 0 32660 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_350
timestamp 1667941163
transform 1 0 33304 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_362
timestamp 1667941163
transform 1 0 34408 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1667941163
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_401
timestamp 1667941163
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_11
timestamp 1667941163
transform 1 0 2116 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_22
timestamp 1667941163
transform 1 0 3128 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_33
timestamp 1667941163
transform 1 0 4140 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_40
timestamp 1667941163
transform 1 0 4784 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_47
timestamp 1667941163
transform 1 0 5428 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1667941163
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_63
timestamp 1667941163
transform 1 0 6900 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_67
timestamp 1667941163
transform 1 0 7268 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_74
timestamp 1667941163
transform 1 0 7912 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_80
timestamp 1667941163
transform 1 0 8464 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_90
timestamp 1667941163
transform 1 0 9384 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_98
timestamp 1667941163
transform 1 0 10120 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_103
timestamp 1667941163
transform 1 0 10580 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1667941163
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_119
timestamp 1667941163
transform 1 0 12052 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_123
timestamp 1667941163
transform 1 0 12420 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_130
timestamp 1667941163
transform 1 0 13064 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_142
timestamp 1667941163
transform 1 0 14168 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_154
timestamp 1667941163
transform 1 0 15272 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_162
timestamp 1667941163
transform 1 0 16008 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1667941163
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_179
timestamp 1667941163
transform 1 0 17572 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_187
timestamp 1667941163
transform 1 0 18308 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_192
timestamp 1667941163
transform 1 0 18768 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_204
timestamp 1667941163
transform 1 0 19872 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_221
timestamp 1667941163
transform 1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_237
timestamp 1667941163
transform 1 0 22908 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1667941163
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_261
timestamp 1667941163
transform 1 0 25116 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_265
timestamp 1667941163
transform 1 0 25484 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_269
timestamp 1667941163
transform 1 0 25852 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_277
timestamp 1667941163
transform 1 0 26588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_292
timestamp 1667941163
transform 1 0 27968 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_304
timestamp 1667941163
transform 1 0 29072 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_319
timestamp 1667941163
transform 1 0 30452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_331
timestamp 1667941163
transform 1 0 31556 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1667941163
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_348
timestamp 1667941163
transform 1 0 33120 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_360
timestamp 1667941163
transform 1 0 34224 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_372
timestamp 1667941163
transform 1 0 35328 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_384
timestamp 1667941163
transform 1 0 36432 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_401
timestamp 1667941163
transform 1 0 37996 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1667941163
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_14
timestamp 1667941163
transform 1 0 2392 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_22
timestamp 1667941163
transform 1 0 3128 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1667941163
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_39
timestamp 1667941163
transform 1 0 4692 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_50
timestamp 1667941163
transform 1 0 5704 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_57
timestamp 1667941163
transform 1 0 6348 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_66
timestamp 1667941163
transform 1 0 7176 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_70
timestamp 1667941163
transform 1 0 7544 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_74
timestamp 1667941163
transform 1 0 7912 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_78
timestamp 1667941163
transform 1 0 8280 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1667941163
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_96
timestamp 1667941163
transform 1 0 9936 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_112
timestamp 1667941163
transform 1 0 11408 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_125
timestamp 1667941163
transform 1 0 12604 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_133
timestamp 1667941163
transform 1 0 13340 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1667941163
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_146
timestamp 1667941163
transform 1 0 14536 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_158
timestamp 1667941163
transform 1 0 15640 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_174
timestamp 1667941163
transform 1 0 17112 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_186
timestamp 1667941163
transform 1 0 18216 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_190
timestamp 1667941163
transform 1 0 18584 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1667941163
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_201
timestamp 1667941163
transform 1 0 19596 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_211
timestamp 1667941163
transform 1 0 20516 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_223
timestamp 1667941163
transform 1 0 21620 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_228
timestamp 1667941163
transform 1 0 22080 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_235
timestamp 1667941163
transform 1 0 22724 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_247
timestamp 1667941163
transform 1 0 23828 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1667941163
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1667941163
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_277
timestamp 1667941163
transform 1 0 26588 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_282
timestamp 1667941163
transform 1 0 27048 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_290
timestamp 1667941163
transform 1 0 27784 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_300
timestamp 1667941163
transform 1 0 28704 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_321
timestamp 1667941163
transform 1 0 30636 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_326
timestamp 1667941163
transform 1 0 31096 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_334
timestamp 1667941163
transform 1 0 31832 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_338
timestamp 1667941163
transform 1 0 32200 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_350
timestamp 1667941163
transform 1 0 33304 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_362
timestamp 1667941163
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1667941163
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1667941163
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_8
timestamp 1667941163
transform 1 0 1840 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_20
timestamp 1667941163
transform 1 0 2944 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_32
timestamp 1667941163
transform 1 0 4048 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_44
timestamp 1667941163
transform 1 0 5152 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_50
timestamp 1667941163
transform 1 0 5704 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_68
timestamp 1667941163
transform 1 0 7360 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_76
timestamp 1667941163
transform 1 0 8096 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_91
timestamp 1667941163
transform 1 0 9476 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_98
timestamp 1667941163
transform 1 0 10120 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1667941163
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_122
timestamp 1667941163
transform 1 0 12328 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_135
timestamp 1667941163
transform 1 0 13524 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_139
timestamp 1667941163
transform 1 0 13892 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1667941163
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1667941163
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1667941163
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_178
timestamp 1667941163
transform 1 0 17480 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_185
timestamp 1667941163
transform 1 0 18124 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_198
timestamp 1667941163
transform 1 0 19320 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_210
timestamp 1667941163
transform 1 0 20424 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_219
timestamp 1667941163
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1667941163
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_235
timestamp 1667941163
transform 1 0 22724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_250
timestamp 1667941163
transform 1 0 24104 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_263
timestamp 1667941163
transform 1 0 25300 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_270
timestamp 1667941163
transform 1 0 25944 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1667941163
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_293
timestamp 1667941163
transform 1 0 28060 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_300
timestamp 1667941163
transform 1 0 28704 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_307
timestamp 1667941163
transform 1 0 29348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_319
timestamp 1667941163
transform 1 0 30452 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_328
timestamp 1667941163
transform 1 0 31280 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1667941163
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1667941163
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1667941163
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1667941163
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1667941163
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1667941163
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1667941163
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_35
timestamp 1667941163
transform 1 0 4324 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_39
timestamp 1667941163
transform 1 0 4692 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_46
timestamp 1667941163
transform 1 0 5336 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_59
timestamp 1667941163
transform 1 0 6532 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_71
timestamp 1667941163
transform 1 0 7636 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_78
timestamp 1667941163
transform 1 0 8280 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_91
timestamp 1667941163
transform 1 0 9476 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_103
timestamp 1667941163
transform 1 0 10580 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_107
timestamp 1667941163
transform 1 0 10948 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_111
timestamp 1667941163
transform 1 0 11316 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_126
timestamp 1667941163
transform 1 0 12696 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1667941163
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_146
timestamp 1667941163
transform 1 0 14536 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_158
timestamp 1667941163
transform 1 0 15640 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_165
timestamp 1667941163
transform 1 0 16284 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_173
timestamp 1667941163
transform 1 0 17020 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_187
timestamp 1667941163
transform 1 0 18308 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1667941163
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_209
timestamp 1667941163
transform 1 0 20332 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1667941163
transform 1 0 20884 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1667941163
transform 1 0 21252 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_223
timestamp 1667941163
transform 1 0 21620 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_229
timestamp 1667941163
transform 1 0 22172 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1667941163
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1667941163
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1667941163
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_263
timestamp 1667941163
transform 1 0 25300 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_275
timestamp 1667941163
transform 1 0 26404 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_287
timestamp 1667941163
transform 1 0 27508 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_296
timestamp 1667941163
transform 1 0 28336 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_316
timestamp 1667941163
transform 1 0 30176 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_328
timestamp 1667941163
transform 1 0 31280 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_340
timestamp 1667941163
transform 1 0 32384 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_352
timestamp 1667941163
transform 1 0 33488 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1667941163
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1667941163
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_401
timestamp 1667941163
transform 1 0 37996 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_9
timestamp 1667941163
transform 1 0 1932 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_21
timestamp 1667941163
transform 1 0 3036 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_33
timestamp 1667941163
transform 1 0 4140 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_42
timestamp 1667941163
transform 1 0 4968 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_49
timestamp 1667941163
transform 1 0 5612 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1667941163
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1667941163
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_96
timestamp 1667941163
transform 1 0 9936 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_104
timestamp 1667941163
transform 1 0 10672 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1667941163
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_119
timestamp 1667941163
transform 1 0 12052 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_131
timestamp 1667941163
transform 1 0 13156 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_139
timestamp 1667941163
transform 1 0 13892 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_149
timestamp 1667941163
transform 1 0 14812 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1667941163
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1667941163
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_173
timestamp 1667941163
transform 1 0 17020 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_177
timestamp 1667941163
transform 1 0 17388 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_190
timestamp 1667941163
transform 1 0 18584 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_196
timestamp 1667941163
transform 1 0 19136 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_200
timestamp 1667941163
transform 1 0 19504 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_206
timestamp 1667941163
transform 1 0 20056 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_215
timestamp 1667941163
transform 1 0 20884 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1667941163
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_230
timestamp 1667941163
transform 1 0 22264 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_242
timestamp 1667941163
transform 1 0 23368 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_254
timestamp 1667941163
transform 1 0 24472 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_266
timestamp 1667941163
transform 1 0 25576 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1667941163
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_286
timestamp 1667941163
transform 1 0 27416 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_298
timestamp 1667941163
transform 1 0 28520 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_310
timestamp 1667941163
transform 1 0 29624 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_320
timestamp 1667941163
transform 1 0 30544 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_332
timestamp 1667941163
transform 1 0 31648 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1667941163
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1667941163
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1667941163
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1667941163
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1667941163
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1667941163
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1667941163
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1667941163
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_41
timestamp 1667941163
transform 1 0 4876 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_51
timestamp 1667941163
transform 1 0 5796 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_58
timestamp 1667941163
transform 1 0 6440 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_70
timestamp 1667941163
transform 1 0 7544 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1667941163
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_93
timestamp 1667941163
transform 1 0 9660 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_97
timestamp 1667941163
transform 1 0 10028 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_110
timestamp 1667941163
transform 1 0 11224 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_118
timestamp 1667941163
transform 1 0 11960 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_122
timestamp 1667941163
transform 1 0 12328 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_129
timestamp 1667941163
transform 1 0 12972 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_137
timestamp 1667941163
transform 1 0 13708 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_146
timestamp 1667941163
transform 1 0 14536 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_153
timestamp 1667941163
transform 1 0 15180 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_157
timestamp 1667941163
transform 1 0 15548 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_161
timestamp 1667941163
transform 1 0 15916 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_168
timestamp 1667941163
transform 1 0 16560 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_172
timestamp 1667941163
transform 1 0 16928 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_182
timestamp 1667941163
transform 1 0 17848 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1667941163
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_209
timestamp 1667941163
transform 1 0 20332 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_217
timestamp 1667941163
transform 1 0 21068 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_222
timestamp 1667941163
transform 1 0 21528 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_230
timestamp 1667941163
transform 1 0 22264 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_241
timestamp 1667941163
transform 1 0 23276 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_249
timestamp 1667941163
transform 1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_265
timestamp 1667941163
transform 1 0 25484 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_275
timestamp 1667941163
transform 1 0 26404 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_288
timestamp 1667941163
transform 1 0 27600 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_296
timestamp 1667941163
transform 1 0 28336 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_300
timestamp 1667941163
transform 1 0 28704 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_313
timestamp 1667941163
transform 1 0 29900 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_317
timestamp 1667941163
transform 1 0 30268 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_324
timestamp 1667941163
transform 1 0 30912 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_331
timestamp 1667941163
transform 1 0 31556 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_343
timestamp 1667941163
transform 1 0 32660 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_355
timestamp 1667941163
transform 1 0 33764 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1667941163
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1667941163
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_401
timestamp 1667941163
transform 1 0 37996 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_15
timestamp 1667941163
transform 1 0 2484 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_26
timestamp 1667941163
transform 1 0 3496 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_38
timestamp 1667941163
transform 1 0 4600 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_50
timestamp 1667941163
transform 1 0 5704 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1667941163
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_62
timestamp 1667941163
transform 1 0 6808 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_74
timestamp 1667941163
transform 1 0 7912 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_84
timestamp 1667941163
transform 1 0 8832 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_96
timestamp 1667941163
transform 1 0 9936 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_104
timestamp 1667941163
transform 1 0 10672 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1667941163
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_120
timestamp 1667941163
transform 1 0 12144 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_132
timestamp 1667941163
transform 1 0 13248 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_144
timestamp 1667941163
transform 1 0 14352 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_148
timestamp 1667941163
transform 1 0 14720 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_156
timestamp 1667941163
transform 1 0 15456 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1667941163
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1667941163
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1667941163
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_205
timestamp 1667941163
transform 1 0 19964 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_213
timestamp 1667941163
transform 1 0 20700 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1667941163
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_237
timestamp 1667941163
transform 1 0 22908 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_241
timestamp 1667941163
transform 1 0 23276 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_251
timestamp 1667941163
transform 1 0 24196 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_262
timestamp 1667941163
transform 1 0 25208 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_266
timestamp 1667941163
transform 1 0 25576 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_270
timestamp 1667941163
transform 1 0 25944 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_277
timestamp 1667941163
transform 1 0 26588 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_286
timestamp 1667941163
transform 1 0 27416 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_292
timestamp 1667941163
transform 1 0 27968 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_301
timestamp 1667941163
transform 1 0 28796 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_314
timestamp 1667941163
transform 1 0 29992 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_326
timestamp 1667941163
transform 1 0 31096 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_334
timestamp 1667941163
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1667941163
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1667941163
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1667941163
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1667941163
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1667941163
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_8
timestamp 1667941163
transform 1 0 1840 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_20
timestamp 1667941163
transform 1 0 2944 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_44
timestamp 1667941163
transform 1 0 5152 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_56
timestamp 1667941163
transform 1 0 6256 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_34_67
timestamp 1667941163
transform 1 0 7268 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1667941163
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_90
timestamp 1667941163
transform 1 0 9384 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_94
timestamp 1667941163
transform 1 0 9752 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_98
timestamp 1667941163
transform 1 0 10120 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_110
timestamp 1667941163
transform 1 0 11224 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_122
timestamp 1667941163
transform 1 0 12328 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_128
timestamp 1667941163
transform 1 0 12880 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_132
timestamp 1667941163
transform 1 0 13248 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_147
timestamp 1667941163
transform 1 0 14628 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_160
timestamp 1667941163
transform 1 0 15824 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_172
timestamp 1667941163
transform 1 0 16928 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_185
timestamp 1667941163
transform 1 0 18124 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_193
timestamp 1667941163
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_202
timestamp 1667941163
transform 1 0 19688 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_210
timestamp 1667941163
transform 1 0 20424 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_215
timestamp 1667941163
transform 1 0 20884 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_227
timestamp 1667941163
transform 1 0 21988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_239
timestamp 1667941163
transform 1 0 23092 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1667941163
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_261
timestamp 1667941163
transform 1 0 25116 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_267
timestamp 1667941163
transform 1 0 25668 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_279
timestamp 1667941163
transform 1 0 26772 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_287
timestamp 1667941163
transform 1 0 27508 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_291
timestamp 1667941163
transform 1 0 27876 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_298
timestamp 1667941163
transform 1 0 28520 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_306
timestamp 1667941163
transform 1 0 29256 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_314
timestamp 1667941163
transform 1 0 29992 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1667941163
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1667941163
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1667941163
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1667941163
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1667941163
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1667941163
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_401
timestamp 1667941163
transform 1 0 37996 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_405
timestamp 1667941163
transform 1 0 38364 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1667941163
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1667941163
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1667941163
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1667941163
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1667941163
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_35_68
timestamp 1667941163
transform 1 0 7360 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_77
timestamp 1667941163
transform 1 0 8188 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_81
timestamp 1667941163
transform 1 0 8556 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_85
timestamp 1667941163
transform 1 0 8924 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_102
timestamp 1667941163
transform 1 0 10488 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_109
timestamp 1667941163
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_122
timestamp 1667941163
transform 1 0 12328 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_130
timestamp 1667941163
transform 1 0 13064 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_140
timestamp 1667941163
transform 1 0 13984 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_152
timestamp 1667941163
transform 1 0 15088 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_164
timestamp 1667941163
transform 1 0 16192 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_190
timestamp 1667941163
transform 1 0 18584 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_211
timestamp 1667941163
transform 1 0 20516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1667941163
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_236
timestamp 1667941163
transform 1 0 22816 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_248
timestamp 1667941163
transform 1 0 23920 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_260
timestamp 1667941163
transform 1 0 25024 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_272
timestamp 1667941163
transform 1 0 26128 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_301
timestamp 1667941163
transform 1 0 28796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_308
timestamp 1667941163
transform 1 0 29440 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_315
timestamp 1667941163
transform 1 0 30084 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_327
timestamp 1667941163
transform 1 0 31188 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1667941163
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1667941163
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1667941163
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1667941163
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1667941163
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1667941163
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1667941163
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1667941163
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_53
timestamp 1667941163
transform 1 0 5980 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_59
timestamp 1667941163
transform 1 0 6532 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_72
timestamp 1667941163
transform 1 0 7728 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_36_81
timestamp 1667941163
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_90
timestamp 1667941163
transform 1 0 9384 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_36_106
timestamp 1667941163
transform 1 0 10856 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_112
timestamp 1667941163
transform 1 0 11408 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_116
timestamp 1667941163
transform 1 0 11776 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_128
timestamp 1667941163
transform 1 0 12880 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1667941163
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1667941163
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_153
timestamp 1667941163
transform 1 0 15180 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_161
timestamp 1667941163
transform 1 0 15916 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_166
timestamp 1667941163
transform 1 0 16376 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_178
timestamp 1667941163
transform 1 0 17480 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_190
timestamp 1667941163
transform 1 0 18584 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_205
timestamp 1667941163
transform 1 0 19964 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_211
timestamp 1667941163
transform 1 0 20516 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_218
timestamp 1667941163
transform 1 0 21160 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_235
timestamp 1667941163
transform 1 0 22724 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_242
timestamp 1667941163
transform 1 0 23368 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1667941163
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_258
timestamp 1667941163
transform 1 0 24840 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_266
timestamp 1667941163
transform 1 0 25576 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_272
timestamp 1667941163
transform 1 0 26128 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_279
timestamp 1667941163
transform 1 0 26772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_291
timestamp 1667941163
transform 1 0 27876 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_296
timestamp 1667941163
transform 1 0 28336 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_303
timestamp 1667941163
transform 1 0 28980 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1667941163
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_319
timestamp 1667941163
transform 1 0 30452 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_326
timestamp 1667941163
transform 1 0 31096 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_338
timestamp 1667941163
transform 1 0 32200 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_350
timestamp 1667941163
transform 1 0 33304 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_362
timestamp 1667941163
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1667941163
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_389
timestamp 1667941163
transform 1 0 36892 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_405
timestamp 1667941163
transform 1 0 38364 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_8
timestamp 1667941163
transform 1 0 1840 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_20
timestamp 1667941163
transform 1 0 2944 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_25
timestamp 1667941163
transform 1 0 3404 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_37
timestamp 1667941163
transform 1 0 4508 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1667941163
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1667941163
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_81
timestamp 1667941163
transform 1 0 8556 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_91
timestamp 1667941163
transform 1 0 9476 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_102
timestamp 1667941163
transform 1 0 10488 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1667941163
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_124
timestamp 1667941163
transform 1 0 12512 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_135
timestamp 1667941163
transform 1 0 13524 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_147
timestamp 1667941163
transform 1 0 14628 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_151
timestamp 1667941163
transform 1 0 14996 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_155
timestamp 1667941163
transform 1 0 15364 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1667941163
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_175
timestamp 1667941163
transform 1 0 17204 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_183
timestamp 1667941163
transform 1 0 17940 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_187
timestamp 1667941163
transform 1 0 18308 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_194
timestamp 1667941163
transform 1 0 18952 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_202
timestamp 1667941163
transform 1 0 19688 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_206
timestamp 1667941163
transform 1 0 20056 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_218
timestamp 1667941163
transform 1 0 21160 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1667941163
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_238
timestamp 1667941163
transform 1 0 23000 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_242
timestamp 1667941163
transform 1 0 23368 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_252
timestamp 1667941163
transform 1 0 24288 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_264
timestamp 1667941163
transform 1 0 25392 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_276
timestamp 1667941163
transform 1 0 26496 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_286
timestamp 1667941163
transform 1 0 27416 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_293
timestamp 1667941163
transform 1 0 28060 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1667941163
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_317
timestamp 1667941163
transform 1 0 30268 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_327
timestamp 1667941163
transform 1 0 31188 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1667941163
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1667941163
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1667941163
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1667941163
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1667941163
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1667941163
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1667941163
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1667941163
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1667941163
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_65
timestamp 1667941163
transform 1 0 7084 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_76
timestamp 1667941163
transform 1 0 8096 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1667941163
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_109
timestamp 1667941163
transform 1 0 11132 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_117
timestamp 1667941163
transform 1 0 11868 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_123
timestamp 1667941163
transform 1 0 12420 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_135
timestamp 1667941163
transform 1 0 13524 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1667941163
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_156
timestamp 1667941163
transform 1 0 15456 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_168
timestamp 1667941163
transform 1 0 16560 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_38_177
timestamp 1667941163
transform 1 0 17388 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_186
timestamp 1667941163
transform 1 0 18216 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1667941163
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_201
timestamp 1667941163
transform 1 0 19596 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_205
timestamp 1667941163
transform 1 0 19964 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_212
timestamp 1667941163
transform 1 0 20608 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_220
timestamp 1667941163
transform 1 0 21344 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_226
timestamp 1667941163
transform 1 0 21896 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_238
timestamp 1667941163
transform 1 0 23000 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1667941163
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_261
timestamp 1667941163
transform 1 0 25116 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_267
timestamp 1667941163
transform 1 0 25668 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_274
timestamp 1667941163
transform 1 0 26312 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_280
timestamp 1667941163
transform 1 0 26864 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_289
timestamp 1667941163
transform 1 0 27692 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_303
timestamp 1667941163
transform 1 0 28980 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1667941163
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_319
timestamp 1667941163
transform 1 0 30452 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_330
timestamp 1667941163
transform 1 0 31464 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_342
timestamp 1667941163
transform 1 0 32568 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_354
timestamp 1667941163
transform 1 0 33672 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_362
timestamp 1667941163
transform 1 0 34408 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_370
timestamp 1667941163
transform 1 0 35144 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_382
timestamp 1667941163
transform 1 0 36248 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_394
timestamp 1667941163
transform 1 0 37352 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_406
timestamp 1667941163
transform 1 0 38456 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1667941163
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1667941163
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1667941163
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1667941163
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1667941163
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_68
timestamp 1667941163
transform 1 0 7360 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_80
timestamp 1667941163
transform 1 0 8464 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_92
timestamp 1667941163
transform 1 0 9568 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_100
timestamp 1667941163
transform 1 0 10304 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1667941163
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_119
timestamp 1667941163
transform 1 0 12052 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_128
timestamp 1667941163
transform 1 0 12880 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_135
timestamp 1667941163
transform 1 0 13524 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_147
timestamp 1667941163
transform 1 0 14628 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_152
timestamp 1667941163
transform 1 0 15088 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 1667941163
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_180
timestamp 1667941163
transform 1 0 17664 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_192
timestamp 1667941163
transform 1 0 18768 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_204
timestamp 1667941163
transform 1 0 19872 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_216
timestamp 1667941163
transform 1 0 20976 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1667941163
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_231
timestamp 1667941163
transform 1 0 22356 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_241
timestamp 1667941163
transform 1 0 23276 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_253
timestamp 1667941163
transform 1 0 24380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_265
timestamp 1667941163
transform 1 0 25484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_277
timestamp 1667941163
transform 1 0 26588 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1667941163
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_308
timestamp 1667941163
transform 1 0 29440 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_316
timestamp 1667941163
transform 1 0 30176 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_322
timestamp 1667941163
transform 1 0 30728 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_334
timestamp 1667941163
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_342
timestamp 1667941163
transform 1 0 32568 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_353
timestamp 1667941163
transform 1 0 33580 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_365
timestamp 1667941163
transform 1 0 34684 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_377
timestamp 1667941163
transform 1 0 35788 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_389
timestamp 1667941163
transform 1 0 36892 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1667941163
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_9
timestamp 1667941163
transform 1 0 1932 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_21
timestamp 1667941163
transform 1 0 3036 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1667941163
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_36
timestamp 1667941163
transform 1 0 4416 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_48
timestamp 1667941163
transform 1 0 5520 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_60
timestamp 1667941163
transform 1 0 6624 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_68
timestamp 1667941163
transform 1 0 7360 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_78
timestamp 1667941163
transform 1 0 8280 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_97
timestamp 1667941163
transform 1 0 10028 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_101
timestamp 1667941163
transform 1 0 10396 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_105
timestamp 1667941163
transform 1 0 10764 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_112
timestamp 1667941163
transform 1 0 11408 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_124
timestamp 1667941163
transform 1 0 12512 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_130
timestamp 1667941163
transform 1 0 13064 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_137
timestamp 1667941163
transform 1 0 13708 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_153
timestamp 1667941163
transform 1 0 15180 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_164
timestamp 1667941163
transform 1 0 16192 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_176
timestamp 1667941163
transform 1 0 17296 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_184
timestamp 1667941163
transform 1 0 18032 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1667941163
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_209
timestamp 1667941163
transform 1 0 20332 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_216
timestamp 1667941163
transform 1 0 20976 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_224
timestamp 1667941163
transform 1 0 21712 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_230
timestamp 1667941163
transform 1 0 22264 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_242
timestamp 1667941163
transform 1 0 23368 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1667941163
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_259
timestamp 1667941163
transform 1 0 24932 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_272
timestamp 1667941163
transform 1 0 26128 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_284
timestamp 1667941163
transform 1 0 27232 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_292
timestamp 1667941163
transform 1 0 27968 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_299
timestamp 1667941163
transform 1 0 28612 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1667941163
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_321
timestamp 1667941163
transform 1 0 30636 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_327
timestamp 1667941163
transform 1 0 31188 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_331
timestamp 1667941163
transform 1 0 31556 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_338
timestamp 1667941163
transform 1 0 32200 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_350
timestamp 1667941163
transform 1 0 33304 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_362
timestamp 1667941163
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1667941163
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1667941163
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_401
timestamp 1667941163
transform 1 0 37996 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_405
timestamp 1667941163
transform 1 0 38364 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1667941163
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1667941163
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_39
timestamp 1667941163
transform 1 0 4692 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_45
timestamp 1667941163
transform 1 0 5244 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_49
timestamp 1667941163
transform 1 0 5612 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1667941163
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_69
timestamp 1667941163
transform 1 0 7452 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_73
timestamp 1667941163
transform 1 0 7820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_85
timestamp 1667941163
transform 1 0 8924 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_97
timestamp 1667941163
transform 1 0 10028 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_105
timestamp 1667941163
transform 1 0 10764 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_109
timestamp 1667941163
transform 1 0 11132 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_121
timestamp 1667941163
transform 1 0 12236 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_125
timestamp 1667941163
transform 1 0 12604 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_137
timestamp 1667941163
transform 1 0 13708 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_145
timestamp 1667941163
transform 1 0 14444 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_157
timestamp 1667941163
transform 1 0 15548 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_165
timestamp 1667941163
transform 1 0 16284 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1667941163
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1667941163
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1667941163
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1667941163
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1667941163
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_236
timestamp 1667941163
transform 1 0 22816 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_248
timestamp 1667941163
transform 1 0 23920 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_260
timestamp 1667941163
transform 1 0 25024 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_272
timestamp 1667941163
transform 1 0 26128 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_286
timestamp 1667941163
transform 1 0 27416 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_298
timestamp 1667941163
transform 1 0 28520 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_310
timestamp 1667941163
transform 1 0 29624 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_322
timestamp 1667941163
transform 1 0 30728 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_334
timestamp 1667941163
transform 1 0 31832 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1667941163
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1667941163
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1667941163
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1667941163
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1667941163
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_8
timestamp 1667941163
transform 1 0 1840 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_20
timestamp 1667941163
transform 1 0 2944 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1667941163
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1667941163
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_80
timestamp 1667941163
transform 1 0 8464 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_93
timestamp 1667941163
transform 1 0 9660 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1667941163
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_109
timestamp 1667941163
transform 1 0 11132 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_116
timestamp 1667941163
transform 1 0 11776 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_124
timestamp 1667941163
transform 1 0 12512 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_134
timestamp 1667941163
transform 1 0 13432 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_153
timestamp 1667941163
transform 1 0 15180 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_159
timestamp 1667941163
transform 1 0 15732 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_166
timestamp 1667941163
transform 1 0 16376 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_173
timestamp 1667941163
transform 1 0 17020 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_185
timestamp 1667941163
transform 1 0 18124 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1667941163
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_208
timestamp 1667941163
transform 1 0 20240 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_220
timestamp 1667941163
transform 1 0 21344 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_232
timestamp 1667941163
transform 1 0 22448 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_244
timestamp 1667941163
transform 1 0 23552 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_268
timestamp 1667941163
transform 1 0 25760 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_280
timestamp 1667941163
transform 1 0 26864 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_292
timestamp 1667941163
transform 1 0 27968 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_299
timestamp 1667941163
transform 1 0 28612 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1667941163
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1667941163
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_341
timestamp 1667941163
transform 1 0 32476 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_353
timestamp 1667941163
transform 1 0 33580 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_361
timestamp 1667941163
transform 1 0 34316 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1667941163
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_401
timestamp 1667941163
transform 1 0 37996 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_405
timestamp 1667941163
transform 1 0 38364 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1667941163
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1667941163
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1667941163
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1667941163
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1667941163
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_65
timestamp 1667941163
transform 1 0 7084 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_75
timestamp 1667941163
transform 1 0 8004 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_83
timestamp 1667941163
transform 1 0 8740 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1667941163
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_105
timestamp 1667941163
transform 1 0 10764 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1667941163
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_123
timestamp 1667941163
transform 1 0 12420 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_130
timestamp 1667941163
transform 1 0 13064 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_137
timestamp 1667941163
transform 1 0 13708 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_143
timestamp 1667941163
transform 1 0 14260 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_147
timestamp 1667941163
transform 1 0 14628 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1667941163
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1667941163
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_196
timestamp 1667941163
transform 1 0 19136 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_204
timestamp 1667941163
transform 1 0 19872 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_210
timestamp 1667941163
transform 1 0 20424 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1667941163
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1667941163
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_246
timestamp 1667941163
transform 1 0 23736 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_259
timestamp 1667941163
transform 1 0 24932 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_271
timestamp 1667941163
transform 1 0 26036 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_275
timestamp 1667941163
transform 1 0 26404 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1667941163
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_291
timestamp 1667941163
transform 1 0 27876 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_303
timestamp 1667941163
transform 1 0 28980 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_315
timestamp 1667941163
transform 1 0 30084 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_327
timestamp 1667941163
transform 1 0 31188 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1667941163
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1667941163
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1667941163
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1667941163
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1667941163
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1667941163
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1667941163
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1667941163
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1667941163
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_65
timestamp 1667941163
transform 1 0 7084 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_70
timestamp 1667941163
transform 1 0 7544 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_82
timestamp 1667941163
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_95
timestamp 1667941163
transform 1 0 9844 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_107
timestamp 1667941163
transform 1 0 10948 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_122
timestamp 1667941163
transform 1 0 12328 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_129
timestamp 1667941163
transform 1 0 12972 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1667941163
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_148
timestamp 1667941163
transform 1 0 14720 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_160
timestamp 1667941163
transform 1 0 15824 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_166
timestamp 1667941163
transform 1 0 16376 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_175
timestamp 1667941163
transform 1 0 17204 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_182
timestamp 1667941163
transform 1 0 17848 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1667941163
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_205
timestamp 1667941163
transform 1 0 19964 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_210
timestamp 1667941163
transform 1 0 20424 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_223
timestamp 1667941163
transform 1 0 21620 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_235
timestamp 1667941163
transform 1 0 22724 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_242
timestamp 1667941163
transform 1 0 23368 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 1667941163
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_44_262
timestamp 1667941163
transform 1 0 25208 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_44_278
timestamp 1667941163
transform 1 0 26680 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_294
timestamp 1667941163
transform 1 0 28152 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_300
timestamp 1667941163
transform 1 0 28704 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_304
timestamp 1667941163
transform 1 0 29072 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1667941163
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1667941163
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1667941163
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1667941163
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1667941163
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1667941163
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1667941163
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_401
timestamp 1667941163
transform 1 0 37996 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1667941163
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1667941163
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1667941163
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1667941163
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1667941163
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_73
timestamp 1667941163
transform 1 0 7820 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_88
timestamp 1667941163
transform 1 0 9200 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_96
timestamp 1667941163
transform 1 0 9936 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_101
timestamp 1667941163
transform 1 0 10396 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_108
timestamp 1667941163
transform 1 0 11040 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_118
timestamp 1667941163
transform 1 0 11960 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_130
timestamp 1667941163
transform 1 0 13064 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_140
timestamp 1667941163
transform 1 0 13984 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_45_156
timestamp 1667941163
transform 1 0 15456 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_162
timestamp 1667941163
transform 1 0 16008 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1667941163
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_178
timestamp 1667941163
transform 1 0 17480 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_182
timestamp 1667941163
transform 1 0 17848 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_187
timestamp 1667941163
transform 1 0 18308 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_195
timestamp 1667941163
transform 1 0 19044 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_199
timestamp 1667941163
transform 1 0 19412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_211
timestamp 1667941163
transform 1 0 20516 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_215
timestamp 1667941163
transform 1 0 20884 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_219
timestamp 1667941163
transform 1 0 21252 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1667941163
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_230
timestamp 1667941163
transform 1 0 22264 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_237
timestamp 1667941163
transform 1 0 22908 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_244
timestamp 1667941163
transform 1 0 23552 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_251
timestamp 1667941163
transform 1 0 24196 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_259
timestamp 1667941163
transform 1 0 24932 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_264
timestamp 1667941163
transform 1 0 25392 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_271
timestamp 1667941163
transform 1 0 26036 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_278
timestamp 1667941163
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1667941163
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1667941163
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1667941163
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1667941163
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1667941163
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_343
timestamp 1667941163
transform 1 0 32660 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_355
timestamp 1667941163
transform 1 0 33764 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_367
timestamp 1667941163
transform 1 0 34868 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_379
timestamp 1667941163
transform 1 0 35972 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1667941163
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1667941163
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_8
timestamp 1667941163
transform 1 0 1840 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_20
timestamp 1667941163
transform 1 0 2944 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_49
timestamp 1667941163
transform 1 0 5612 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_53
timestamp 1667941163
transform 1 0 5980 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_62
timestamp 1667941163
transform 1 0 6808 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_69
timestamp 1667941163
transform 1 0 7452 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_76
timestamp 1667941163
transform 1 0 8096 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_90
timestamp 1667941163
transform 1 0 9384 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_106
timestamp 1667941163
transform 1 0 10856 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_118
timestamp 1667941163
transform 1 0 11960 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_129
timestamp 1667941163
transform 1 0 12972 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_137
timestamp 1667941163
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1667941163
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_165
timestamp 1667941163
transform 1 0 16284 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_169
timestamp 1667941163
transform 1 0 16652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_173
timestamp 1667941163
transform 1 0 17020 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_186
timestamp 1667941163
transform 1 0 18216 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1667941163
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1667941163
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1667941163
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1667941163
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1667941163
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1667941163
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_265
timestamp 1667941163
transform 1 0 25484 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_273
timestamp 1667941163
transform 1 0 26220 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_283
timestamp 1667941163
transform 1 0 27140 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_295
timestamp 1667941163
transform 1 0 28244 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_304
timestamp 1667941163
transform 1 0 29072 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_314
timestamp 1667941163
transform 1 0 29992 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_326
timestamp 1667941163
transform 1 0 31096 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_338
timestamp 1667941163
transform 1 0 32200 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_344
timestamp 1667941163
transform 1 0 32752 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_348
timestamp 1667941163
transform 1 0 33120 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_360
timestamp 1667941163
transform 1 0 34224 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1667941163
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_405
timestamp 1667941163
transform 1 0 38364 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1667941163
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1667941163
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1667941163
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1667941163
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1667941163
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_66
timestamp 1667941163
transform 1 0 7176 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_74
timestamp 1667941163
transform 1 0 7912 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_80
timestamp 1667941163
transform 1 0 8464 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_84
timestamp 1667941163
transform 1 0 8832 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_88
timestamp 1667941163
transform 1 0 9200 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_94
timestamp 1667941163
transform 1 0 9752 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_103
timestamp 1667941163
transform 1 0 10580 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1667941163
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_117
timestamp 1667941163
transform 1 0 11868 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_121
timestamp 1667941163
transform 1 0 12236 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_133
timestamp 1667941163
transform 1 0 13340 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_141
timestamp 1667941163
transform 1 0 14076 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_153
timestamp 1667941163
transform 1 0 15180 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_165
timestamp 1667941163
transform 1 0 16284 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1667941163
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_193
timestamp 1667941163
transform 1 0 18860 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_199
timestamp 1667941163
transform 1 0 19412 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_209
timestamp 1667941163
transform 1 0 20332 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1667941163
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_230
timestamp 1667941163
transform 1 0 22264 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_242
timestamp 1667941163
transform 1 0 23368 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_246
timestamp 1667941163
transform 1 0 23736 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_253
timestamp 1667941163
transform 1 0 24380 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_257
timestamp 1667941163
transform 1 0 24748 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_266
timestamp 1667941163
transform 1 0 25576 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_278
timestamp 1667941163
transform 1 0 26680 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_286
timestamp 1667941163
transform 1 0 27416 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_293
timestamp 1667941163
transform 1 0 28060 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_300
timestamp 1667941163
transform 1 0 28704 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_316
timestamp 1667941163
transform 1 0 30176 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_328
timestamp 1667941163
transform 1 0 31280 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1667941163
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1667941163
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_376
timestamp 1667941163
transform 1 0 35696 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_388
timestamp 1667941163
transform 1 0 36800 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1667941163
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1667941163
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1667941163
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_65
timestamp 1667941163
transform 1 0 7084 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_74
timestamp 1667941163
transform 1 0 7912 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_48_81
timestamp 1667941163
transform 1 0 8556 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_100
timestamp 1667941163
transform 1 0 10304 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_107
timestamp 1667941163
transform 1 0 10948 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_119
timestamp 1667941163
transform 1 0 12052 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_125
timestamp 1667941163
transform 1 0 12604 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_134
timestamp 1667941163
transform 1 0 13432 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_145
timestamp 1667941163
transform 1 0 14444 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_149
timestamp 1667941163
transform 1 0 14812 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_156
timestamp 1667941163
transform 1 0 15456 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_163
timestamp 1667941163
transform 1 0 16100 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_175
timestamp 1667941163
transform 1 0 17204 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_187
timestamp 1667941163
transform 1 0 18308 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1667941163
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_203
timestamp 1667941163
transform 1 0 19780 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_207
timestamp 1667941163
transform 1 0 20148 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_219
timestamp 1667941163
transform 1 0 21252 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_231
timestamp 1667941163
transform 1 0 22356 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_243
timestamp 1667941163
transform 1 0 23460 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1667941163
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1667941163
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1667941163
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1667941163
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_301
timestamp 1667941163
transform 1 0 28796 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_305
timestamp 1667941163
transform 1 0 29164 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_321
timestamp 1667941163
transform 1 0 30636 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_328
timestamp 1667941163
transform 1 0 31280 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_340
timestamp 1667941163
transform 1 0 32384 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_352
timestamp 1667941163
transform 1 0 33488 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1667941163
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1667941163
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_8
timestamp 1667941163
transform 1 0 1840 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_20
timestamp 1667941163
transform 1 0 2944 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_32
timestamp 1667941163
transform 1 0 4048 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_44
timestamp 1667941163
transform 1 0 5152 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_69
timestamp 1667941163
transform 1 0 7452 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_83
timestamp 1667941163
transform 1 0 8740 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_95
timestamp 1667941163
transform 1 0 9844 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_99
timestamp 1667941163
transform 1 0 10212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1667941163
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_120
timestamp 1667941163
transform 1 0 12144 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_132
timestamp 1667941163
transform 1 0 13248 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_144
timestamp 1667941163
transform 1 0 14352 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_153
timestamp 1667941163
transform 1 0 15180 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_165
timestamp 1667941163
transform 1 0 16284 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_181
timestamp 1667941163
transform 1 0 17756 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_188
timestamp 1667941163
transform 1 0 18400 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_196
timestamp 1667941163
transform 1 0 19136 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_200
timestamp 1667941163
transform 1 0 19504 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_207
timestamp 1667941163
transform 1 0 20148 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_213
timestamp 1667941163
transform 1 0 20700 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1667941163
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1667941163
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1667941163
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1667941163
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1667941163
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1667941163
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1667941163
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1667941163
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1667941163
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1667941163
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1667941163
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1667941163
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1667941163
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1667941163
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_401
timestamp 1667941163
transform 1 0 37996 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1667941163
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1667941163
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1667941163
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_41
timestamp 1667941163
transform 1 0 4876 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_46
timestamp 1667941163
transform 1 0 5336 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_58
timestamp 1667941163
transform 1 0 6440 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_69
timestamp 1667941163
transform 1 0 7452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_81
timestamp 1667941163
transform 1 0 8556 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_93
timestamp 1667941163
transform 1 0 9660 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_105
timestamp 1667941163
transform 1 0 10764 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_112
timestamp 1667941163
transform 1 0 11408 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_125
timestamp 1667941163
transform 1 0 12604 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_137
timestamp 1667941163
transform 1 0 13708 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_155
timestamp 1667941163
transform 1 0 15364 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_162
timestamp 1667941163
transform 1 0 16008 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_174
timestamp 1667941163
transform 1 0 17112 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_182
timestamp 1667941163
transform 1 0 17848 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_193
timestamp 1667941163
transform 1 0 18860 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_201
timestamp 1667941163
transform 1 0 19596 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_210
timestamp 1667941163
transform 1 0 20424 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_216
timestamp 1667941163
transform 1 0 20976 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1667941163
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1667941163
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1667941163
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1667941163
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_260
timestamp 1667941163
transform 1 0 25024 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_272
timestamp 1667941163
transform 1 0 26128 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_284
timestamp 1667941163
transform 1 0 27232 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_292
timestamp 1667941163
transform 1 0 27968 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_296
timestamp 1667941163
transform 1 0 28336 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1667941163
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1667941163
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1667941163
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1667941163
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1667941163
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1667941163
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1667941163
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_401
timestamp 1667941163
transform 1 0 37996 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1667941163
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1667941163
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1667941163
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1667941163
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1667941163
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_73
timestamp 1667941163
transform 1 0 7820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_85
timestamp 1667941163
transform 1 0 8924 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_97
timestamp 1667941163
transform 1 0 10028 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_101
timestamp 1667941163
transform 1 0 10396 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1667941163
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1667941163
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_121
timestamp 1667941163
transform 1 0 12236 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_126
timestamp 1667941163
transform 1 0 12696 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_138
timestamp 1667941163
transform 1 0 13800 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_145
timestamp 1667941163
transform 1 0 14444 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_152
timestamp 1667941163
transform 1 0 15088 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_164
timestamp 1667941163
transform 1 0 16192 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_174
timestamp 1667941163
transform 1 0 17112 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_186
timestamp 1667941163
transform 1 0 18216 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_198
timestamp 1667941163
transform 1 0 19320 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_203
timestamp 1667941163
transform 1 0 19780 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_215
timestamp 1667941163
transform 1 0 20884 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1667941163
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_237
timestamp 1667941163
transform 1 0 22908 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_242
timestamp 1667941163
transform 1 0 23368 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_254
timestamp 1667941163
transform 1 0 24472 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_266
timestamp 1667941163
transform 1 0 25576 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_278
timestamp 1667941163
transform 1 0 26680 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_293
timestamp 1667941163
transform 1 0 28060 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_304
timestamp 1667941163
transform 1 0 29072 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_316
timestamp 1667941163
transform 1 0 30176 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_328
timestamp 1667941163
transform 1 0 31280 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_354
timestamp 1667941163
transform 1 0 33672 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_366
timestamp 1667941163
transform 1 0 34776 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_378
timestamp 1667941163
transform 1 0 35880 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_390
timestamp 1667941163
transform 1 0 36984 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1667941163
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1667941163
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1667941163
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1667941163
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1667941163
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1667941163
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1667941163
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1667941163
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_97
timestamp 1667941163
transform 1 0 10028 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_105
timestamp 1667941163
transform 1 0 10764 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_111
timestamp 1667941163
transform 1 0 11316 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_118
timestamp 1667941163
transform 1 0 11960 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_130
timestamp 1667941163
transform 1 0 13064 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1667941163
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_146
timestamp 1667941163
transform 1 0 14536 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_158
timestamp 1667941163
transform 1 0 15640 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_170
timestamp 1667941163
transform 1 0 16744 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_179
timestamp 1667941163
transform 1 0 17572 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_183
timestamp 1667941163
transform 1 0 17940 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_187
timestamp 1667941163
transform 1 0 18308 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1667941163
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_208
timestamp 1667941163
transform 1 0 20240 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_220
timestamp 1667941163
transform 1 0 21344 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_232
timestamp 1667941163
transform 1 0 22448 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_236
timestamp 1667941163
transform 1 0 22816 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_249
timestamp 1667941163
transform 1 0 24012 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1667941163
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1667941163
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1667941163
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1667941163
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1667941163
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1667941163
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1667941163
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_345
timestamp 1667941163
transform 1 0 32844 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_349
timestamp 1667941163
transform 1 0 33212 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_353
timestamp 1667941163
transform 1 0 33580 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_361
timestamp 1667941163
transform 1 0 34316 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1667941163
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1667941163
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_401
timestamp 1667941163
transform 1 0 37996 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1667941163
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1667941163
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1667941163
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1667941163
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1667941163
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1667941163
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1667941163
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1667941163
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1667941163
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1667941163
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1667941163
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1667941163
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_149
timestamp 1667941163
transform 1 0 14812 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_155
timestamp 1667941163
transform 1 0 15364 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_162
timestamp 1667941163
transform 1 0 16008 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1667941163
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_193
timestamp 1667941163
transform 1 0 18860 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_199
timestamp 1667941163
transform 1 0 19412 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_203
timestamp 1667941163
transform 1 0 19780 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_210
timestamp 1667941163
transform 1 0 20424 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1667941163
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1667941163
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_261
timestamp 1667941163
transform 1 0 25116 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_269
timestamp 1667941163
transform 1 0 25852 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1667941163
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1667941163
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1667941163
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1667941163
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_317
timestamp 1667941163
transform 1 0 30268 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_323
timestamp 1667941163
transform 1 0 30820 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1667941163
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1667941163
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1667941163
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1667941163
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1667941163
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1667941163
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1667941163
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1667941163
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1667941163
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1667941163
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1667941163
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1667941163
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1667941163
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1667941163
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_93
timestamp 1667941163
transform 1 0 9660 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_99
timestamp 1667941163
transform 1 0 10212 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_111
timestamp 1667941163
transform 1 0 11316 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_123
timestamp 1667941163
transform 1 0 12420 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_135
timestamp 1667941163
transform 1 0 13524 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1667941163
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_165
timestamp 1667941163
transform 1 0 16284 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_174
timestamp 1667941163
transform 1 0 17112 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_186
timestamp 1667941163
transform 1 0 18216 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_194
timestamp 1667941163
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1667941163
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1667941163
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1667941163
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1667941163
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1667941163
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1667941163
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_277
timestamp 1667941163
transform 1 0 26588 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_282
timestamp 1667941163
transform 1 0 27048 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_294
timestamp 1667941163
transform 1 0 28152 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_306
timestamp 1667941163
transform 1 0 29256 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_316
timestamp 1667941163
transform 1 0 30176 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_328
timestamp 1667941163
transform 1 0 31280 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_340
timestamp 1667941163
transform 1 0 32384 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_352
timestamp 1667941163
transform 1 0 33488 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1667941163
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_401
timestamp 1667941163
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_8
timestamp 1667941163
transform 1 0 1840 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_20
timestamp 1667941163
transform 1 0 2944 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_32
timestamp 1667941163
transform 1 0 4048 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_36
timestamp 1667941163
transform 1 0 4416 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_48
timestamp 1667941163
transform 1 0 5520 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1667941163
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1667941163
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1667941163
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1667941163
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1667941163
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_118
timestamp 1667941163
transform 1 0 11960 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_130
timestamp 1667941163
transform 1 0 13064 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_142
timestamp 1667941163
transform 1 0 14168 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_154
timestamp 1667941163
transform 1 0 15272 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_166
timestamp 1667941163
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_177
timestamp 1667941163
transform 1 0 17388 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1667941163
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1667941163
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1667941163
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1667941163
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1667941163
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1667941163
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1667941163
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1667941163
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1667941163
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1667941163
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_293
timestamp 1667941163
transform 1 0 28060 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_302
timestamp 1667941163
transform 1 0 28888 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_314
timestamp 1667941163
transform 1 0 29992 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_326
timestamp 1667941163
transform 1 0 31096 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_334
timestamp 1667941163
transform 1 0 31832 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1667941163
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1667941163
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1667941163
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1667941163
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1667941163
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1667941163
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1667941163
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1667941163
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1667941163
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1667941163
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1667941163
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1667941163
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_109
timestamp 1667941163
transform 1 0 11132 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_120
timestamp 1667941163
transform 1 0 12144 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_132
timestamp 1667941163
transform 1 0 13248 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1667941163
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1667941163
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1667941163
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1667941163
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1667941163
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1667941163
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1667941163
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1667941163
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1667941163
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1667941163
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1667941163
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1667941163
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1667941163
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1667941163
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_325
timestamp 1667941163
transform 1 0 31004 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_329
timestamp 1667941163
transform 1 0 31372 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_341
timestamp 1667941163
transform 1 0 32476 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_347
timestamp 1667941163
transform 1 0 33028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_359
timestamp 1667941163
transform 1 0 34132 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1667941163
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1667941163
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_401
timestamp 1667941163
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_8
timestamp 1667941163
transform 1 0 1840 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_20
timestamp 1667941163
transform 1 0 2944 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_32
timestamp 1667941163
transform 1 0 4048 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_44
timestamp 1667941163
transform 1 0 5152 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1667941163
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1667941163
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1667941163
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1667941163
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1667941163
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1667941163
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1667941163
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1667941163
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1667941163
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1667941163
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1667941163
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1667941163
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1667941163
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1667941163
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1667941163
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1667941163
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1667941163
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1667941163
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1667941163
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1667941163
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1667941163
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1667941163
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1667941163
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1667941163
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1667941163
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_401
timestamp 1667941163
transform 1 0 37996 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1667941163
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1667941163
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1667941163
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1667941163
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1667941163
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1667941163
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1667941163
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1667941163
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1667941163
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1667941163
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1667941163
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1667941163
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1667941163
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1667941163
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1667941163
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1667941163
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1667941163
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1667941163
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1667941163
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1667941163
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1667941163
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1667941163
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1667941163
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1667941163
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1667941163
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1667941163
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1667941163
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1667941163
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1667941163
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1667941163
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 1667941163
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1667941163
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1667941163
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1667941163
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1667941163
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1667941163
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1667941163
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1667941163
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1667941163
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1667941163
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1667941163
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1667941163
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1667941163
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1667941163
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1667941163
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1667941163
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1667941163
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1667941163
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1667941163
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1667941163
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1667941163
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1667941163
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1667941163
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1667941163
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1667941163
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1667941163
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1667941163
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1667941163
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_329
timestamp 1667941163
transform 1 0 31372 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_59_333
timestamp 1667941163
transform 1 0 31740 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_343
timestamp 1667941163
transform 1 0 32660 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_355
timestamp 1667941163
transform 1 0 33764 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_367
timestamp 1667941163
transform 1 0 34868 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_379
timestamp 1667941163
transform 1 0 35972 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1667941163
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1667941163
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1667941163
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1667941163
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1667941163
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_53
timestamp 1667941163
transform 1 0 5980 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_61
timestamp 1667941163
transform 1 0 6716 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_67
timestamp 1667941163
transform 1 0 7268 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_79
timestamp 1667941163
transform 1 0 8372 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1667941163
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1667941163
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1667941163
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1667941163
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1667941163
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1667941163
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1667941163
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1667941163
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1667941163
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1667941163
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1667941163
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1667941163
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1667941163
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1667941163
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1667941163
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1667941163
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1667941163
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1667941163
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1667941163
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1667941163
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1667941163
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1667941163
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1667941163
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1667941163
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1667941163
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1667941163
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_405
timestamp 1667941163
transform 1 0 38364 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1667941163
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1667941163
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1667941163
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1667941163
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1667941163
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1667941163
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1667941163
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1667941163
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1667941163
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1667941163
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1667941163
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1667941163
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1667941163
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1667941163
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1667941163
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1667941163
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1667941163
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1667941163
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1667941163
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1667941163
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1667941163
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1667941163
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1667941163
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1667941163
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1667941163
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1667941163
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1667941163
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1667941163
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1667941163
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1667941163
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1667941163
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1667941163
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1667941163
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1667941163
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1667941163
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1667941163
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1667941163
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1667941163
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1667941163
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1667941163
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1667941163
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1667941163
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1667941163
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1667941163
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1667941163
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1667941163
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1667941163
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1667941163
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1667941163
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1667941163
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1667941163
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1667941163
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1667941163
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1667941163
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1667941163
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1667941163
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1667941163
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1667941163
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1667941163
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1667941163
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1667941163
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1667941163
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1667941163
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_401
timestamp 1667941163
transform 1 0 37996 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_405
timestamp 1667941163
transform 1 0 38364 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_9
timestamp 1667941163
transform 1 0 1932 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_21
timestamp 1667941163
transform 1 0 3036 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_33
timestamp 1667941163
transform 1 0 4140 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_45
timestamp 1667941163
transform 1 0 5244 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_53
timestamp 1667941163
transform 1 0 5980 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1667941163
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1667941163
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1667941163
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1667941163
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1667941163
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1667941163
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1667941163
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1667941163
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1667941163
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1667941163
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1667941163
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1667941163
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1667941163
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1667941163
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1667941163
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1667941163
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1667941163
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1667941163
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1667941163
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1667941163
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1667941163
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1667941163
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1667941163
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1667941163
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1667941163
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1667941163
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1667941163
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1667941163
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_385
timestamp 1667941163
transform 1 0 36524 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_390
timestamp 1667941163
transform 1 0 36984 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1667941163
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_9
timestamp 1667941163
transform 1 0 1932 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_16
timestamp 1667941163
transform 1 0 2576 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_23
timestamp 1667941163
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1667941163
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_34
timestamp 1667941163
transform 1 0 4232 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1667941163
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_53
timestamp 1667941163
transform 1 0 5980 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_63
timestamp 1667941163
transform 1 0 6900 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_71
timestamp 1667941163
transform 1 0 7636 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1667941163
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1667941163
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_90
timestamp 1667941163
transform 1 0 9384 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_98
timestamp 1667941163
transform 1 0 10120 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_105
timestamp 1667941163
transform 1 0 10764 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_111
timestamp 1667941163
transform 1 0 11316 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_121
timestamp 1667941163
transform 1 0 12236 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_126
timestamp 1667941163
transform 1 0 12696 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_138
timestamp 1667941163
transform 1 0 13800 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_146
timestamp 1667941163
transform 1 0 14536 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_154
timestamp 1667941163
transform 1 0 15272 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_161
timestamp 1667941163
transform 1 0 15916 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_167
timestamp 1667941163
transform 1 0 16468 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_175
timestamp 1667941163
transform 1 0 17204 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_183
timestamp 1667941163
transform 1 0 17940 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_188
timestamp 1667941163
transform 1 0 18400 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_205
timestamp 1667941163
transform 1 0 19964 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_210
timestamp 1667941163
transform 1 0 20424 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_222
timestamp 1667941163
transform 1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_231
timestamp 1667941163
transform 1 0 22356 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_238
timestamp 1667941163
transform 1 0 23000 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_250
timestamp 1667941163
transform 1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_258
timestamp 1667941163
transform 1 0 24840 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_266
timestamp 1667941163
transform 1 0 25576 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_272
timestamp 1667941163
transform 1 0 26128 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_289
timestamp 1667941163
transform 1 0 27692 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_294
timestamp 1667941163
transform 1 0 28152 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_306
timestamp 1667941163
transform 1 0 29256 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_315
timestamp 1667941163
transform 1 0 30084 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_322
timestamp 1667941163
transform 1 0 30728 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_334
timestamp 1667941163
transform 1 0 31832 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_342
timestamp 1667941163
transform 1 0 32568 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_350
timestamp 1667941163
transform 1 0 33304 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_356
timestamp 1667941163
transform 1 0 33856 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_371
timestamp 1667941163
transform 1 0 35236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_383
timestamp 1667941163
transform 1 0 36340 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_390
timestamp 1667941163
transform 1 0 36984 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_393
timestamp 1667941163
transform 1 0 37260 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_405
timestamp 1667941163
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0404_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 9936 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0405_
timestamp 1667941163
transform 1 0 7176 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0406_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 8280 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0407_
timestamp 1667941163
transform 1 0 8188 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0408_
timestamp 1667941163
transform 1 0 11040 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0409_
timestamp 1667941163
transform 1 0 11684 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0410_
timestamp 1667941163
transform 1 0 12052 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0411_
timestamp 1667941163
transform 1 0 22632 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0412_
timestamp 1667941163
transform 1 0 25852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0413_
timestamp 1667941163
transform 1 0 25208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0414_
timestamp 1667941163
transform 1 0 12052 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0415_
timestamp 1667941163
transform 1 0 12052 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0416_
timestamp 1667941163
transform 1 0 24564 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0417_
timestamp 1667941163
transform 1 0 21252 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0418_
timestamp 1667941163
transform 1 0 12052 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0419_
timestamp 1667941163
transform 1 0 12144 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0420_
timestamp 1667941163
transform 1 0 28520 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0421_
timestamp 1667941163
transform 1 0 27876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0422_
timestamp 1667941163
transform 1 0 20792 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0423_
timestamp 1667941163
transform 1 0 28704 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0424_
timestamp 1667941163
transform 1 0 29716 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0425_
timestamp 1667941163
transform 1 0 28704 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0426_
timestamp 1667941163
transform 1 0 4692 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0427_
timestamp 1667941163
transform 1 0 4508 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0428_
timestamp 1667941163
transform 1 0 23552 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0429_
timestamp 1667941163
transform 1 0 4048 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0430_
timestamp 1667941163
transform 1 0 8372 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0431_
timestamp 1667941163
transform 1 0 9844 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0432_
timestamp 1667941163
transform 1 0 24564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0433_
timestamp 1667941163
transform 1 0 25208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0434_
timestamp 1667941163
transform 1 0 15640 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0435_
timestamp 1667941163
transform 1 0 28428 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0436_
timestamp 1667941163
transform 1 0 27140 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0437_
timestamp 1667941163
transform 1 0 27140 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0438_
timestamp 1667941163
transform 1 0 8648 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0439_
timestamp 1667941163
transform 1 0 8280 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0440_
timestamp 1667941163
transform 1 0 11960 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0441_
timestamp 1667941163
transform 1 0 20700 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0442_
timestamp 1667941163
transform 1 0 19780 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0443_
timestamp 1667941163
transform 1 0 19688 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0444_
timestamp 1667941163
transform 1 0 15824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0445_
timestamp 1667941163
transform 1 0 15180 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0446_
timestamp 1667941163
transform 1 0 24564 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0447_
timestamp 1667941163
transform 1 0 9108 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0448_
timestamp 1667941163
transform 1 0 12788 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0449_
timestamp 1667941163
transform 1 0 18492 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0450_
timestamp 1667941163
transform 1 0 27140 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0451_
timestamp 1667941163
transform 1 0 28796 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0452_
timestamp 1667941163
transform 1 0 5336 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0453_
timestamp 1667941163
transform 1 0 5152 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0454_
timestamp 1667941163
transform 1 0 24472 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0455_
timestamp 1667941163
transform 1 0 23276 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0456_
timestamp 1667941163
transform 1 0 26312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0457_
timestamp 1667941163
transform 1 0 27784 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0458_
timestamp 1667941163
transform 1 0 25116 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0459_
timestamp 1667941163
transform 1 0 25760 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0460_
timestamp 1667941163
transform 1 0 29716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0461_
timestamp 1667941163
transform 1 0 24564 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0462_
timestamp 1667941163
transform 1 0 27140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0463_
timestamp 1667941163
transform 1 0 29348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0464_
timestamp 1667941163
transform 1 0 31004 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0465_
timestamp 1667941163
transform 1 0 31556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0466_
timestamp 1667941163
transform 1 0 19412 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0467_
timestamp 1667941163
transform 1 0 27968 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0468_
timestamp 1667941163
transform 1 0 31648 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0469_
timestamp 1667941163
transform 1 0 31924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0470_
timestamp 1667941163
transform 1 0 17112 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0471_
timestamp 1667941163
transform 1 0 16100 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0472_
timestamp 1667941163
transform 1 0 17940 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0473_
timestamp 1667941163
transform 1 0 22264 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0474_
timestamp 1667941163
transform 1 0 23920 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0475_
timestamp 1667941163
transform 1 0 29532 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0476_
timestamp 1667941163
transform 1 0 18860 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0477_
timestamp 1667941163
transform 1 0 19136 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0478_
timestamp 1667941163
transform 1 0 13524 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0479_
timestamp 1667941163
transform 1 0 4692 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0480_
timestamp 1667941163
transform 1 0 5520 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0481_
timestamp 1667941163
transform 1 0 6072 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0482_
timestamp 1667941163
transform 1 0 25116 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0483_
timestamp 1667941163
transform 1 0 28888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0484_
timestamp 1667941163
transform 1 0 25576 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0485_
timestamp 1667941163
transform 1 0 11132 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0486_
timestamp 1667941163
transform 1 0 10856 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0487_
timestamp 1667941163
transform 1 0 9752 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0488_
timestamp 1667941163
transform 1 0 28428 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0489_
timestamp 1667941163
transform 1 0 29716 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0490_
timestamp 1667941163
transform 1 0 21988 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0491_
timestamp 1667941163
transform 1 0 30268 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0492_
timestamp 1667941163
transform 1 0 28520 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0493_
timestamp 1667941163
transform 1 0 30360 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0494_
timestamp 1667941163
transform 1 0 20148 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0495_
timestamp 1667941163
transform 1 0 20148 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0496_
timestamp 1667941163
transform 1 0 18676 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0497_
timestamp 1667941163
transform 1 0 12972 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0498_
timestamp 1667941163
transform 1 0 12328 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0499_
timestamp 1667941163
transform 1 0 13432 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0500_
timestamp 1667941163
transform 1 0 23276 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0501_
timestamp 1667941163
transform 1 0 23920 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0502_
timestamp 1667941163
transform 1 0 9660 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0503_
timestamp 1667941163
transform 1 0 5796 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0504_
timestamp 1667941163
transform 1 0 18676 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0505_
timestamp 1667941163
transform 1 0 18032 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0506_
timestamp 1667941163
transform 1 0 9752 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0507_
timestamp 1667941163
transform 1 0 9844 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0508_
timestamp 1667941163
transform 1 0 16008 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0509_
timestamp 1667941163
transform 1 0 13248 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0510_
timestamp 1667941163
transform 1 0 13064 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0511_
timestamp 1667941163
transform 1 0 15732 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0512_
timestamp 1667941163
transform 1 0 22540 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0513_
timestamp 1667941163
transform 1 0 24932 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0514_
timestamp 1667941163
transform 1 0 25392 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0515_
timestamp 1667941163
transform 1 0 15088 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0516_
timestamp 1667941163
transform 1 0 15732 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0517_
timestamp 1667941163
transform 1 0 19228 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0518_
timestamp 1667941163
transform 1 0 19504 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0519_
timestamp 1667941163
transform 1 0 19504 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0520_
timestamp 1667941163
transform 1 0 28612 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0521_
timestamp 1667941163
transform 1 0 25760 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0522_
timestamp 1667941163
transform 1 0 16928 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0523_
timestamp 1667941163
transform 1 0 15916 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0524_
timestamp 1667941163
transform 1 0 29164 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0525_
timestamp 1667941163
transform 1 0 29808 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0526_
timestamp 1667941163
transform 1 0 29716 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0527_
timestamp 1667941163
transform 1 0 29992 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0528_
timestamp 1667941163
transform 1 0 31280 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0529_
timestamp 1667941163
transform 1 0 23092 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0530_
timestamp 1667941163
transform 1 0 22448 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0531_
timestamp 1667941163
transform 1 0 23460 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0532_
timestamp 1667941163
transform 1 0 25024 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0533_
timestamp 1667941163
transform 1 0 20792 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0534_
timestamp 1667941163
transform 1 0 20976 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0535_
timestamp 1667941163
transform 1 0 14444 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0536_
timestamp 1667941163
transform 1 0 17572 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0537_
timestamp 1667941163
transform 1 0 17204 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0538_
timestamp 1667941163
transform 1 0 7176 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0539_
timestamp 1667941163
transform 1 0 5796 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0540_
timestamp 1667941163
transform 1 0 6992 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0541_
timestamp 1667941163
transform 1 0 7636 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0542_
timestamp 1667941163
transform 1 0 23092 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0543_
timestamp 1667941163
transform 1 0 23736 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0544_
timestamp 1667941163
transform 1 0 23828 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0545_
timestamp 1667941163
transform 1 0 29532 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0546_
timestamp 1667941163
transform 1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0547_
timestamp 1667941163
transform 1 0 16100 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0548_
timestamp 1667941163
transform 1 0 9108 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0549_
timestamp 1667941163
transform 1 0 20332 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0550_
timestamp 1667941163
transform 1 0 21988 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0551_
timestamp 1667941163
transform 1 0 16744 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0552_
timestamp 1667941163
transform 1 0 15456 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0553_
timestamp 1667941163
transform 1 0 16100 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0554_
timestamp 1667941163
transform 1 0 12696 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0555_
timestamp 1667941163
transform 1 0 12052 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0556_
timestamp 1667941163
transform 1 0 25760 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0557_
timestamp 1667941163
transform 1 0 29716 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0558_
timestamp 1667941163
transform 1 0 23460 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0559_
timestamp 1667941163
transform 1 0 24104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0560_
timestamp 1667941163
transform 1 0 24932 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0561_
timestamp 1667941163
transform 1 0 26128 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0562_
timestamp 1667941163
transform 1 0 27140 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0563_
timestamp 1667941163
transform 1 0 27784 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0564_
timestamp 1667941163
transform 1 0 27140 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0565_
timestamp 1667941163
transform 1 0 11040 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0566_
timestamp 1667941163
transform 1 0 16744 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0567_
timestamp 1667941163
transform 1 0 21988 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0568_
timestamp 1667941163
transform 1 0 22632 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0569_
timestamp 1667941163
transform 1 0 10948 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0570_
timestamp 1667941163
transform 1 0 11776 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0571_
timestamp 1667941163
transform 1 0 13248 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0572_
timestamp 1667941163
transform 1 0 13432 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0573_
timestamp 1667941163
transform 1 0 12788 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0574_
timestamp 1667941163
transform 1 0 27508 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0575_
timestamp 1667941163
transform 1 0 30084 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0576_
timestamp 1667941163
transform 1 0 29992 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0577_
timestamp 1667941163
transform 1 0 29992 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0578_
timestamp 1667941163
transform 1 0 27968 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0579_
timestamp 1667941163
transform 1 0 28244 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0580_
timestamp 1667941163
transform 1 0 26772 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0581_
timestamp 1667941163
transform 1 0 28428 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0582_
timestamp 1667941163
transform 1 0 28060 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0583_
timestamp 1667941163
transform 1 0 6532 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0584_
timestamp 1667941163
transform 1 0 4416 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0585_
timestamp 1667941163
transform 1 0 5428 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0586_
timestamp 1667941163
transform 1 0 5336 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0587_
timestamp 1667941163
transform 1 0 6992 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0588_
timestamp 1667941163
transform 1 0 7084 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0589_
timestamp 1667941163
transform 1 0 12696 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0590_
timestamp 1667941163
transform 1 0 10948 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0591_
timestamp 1667941163
transform 1 0 10856 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0592_
timestamp 1667941163
transform 1 0 25668 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0593_
timestamp 1667941163
transform 1 0 23828 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0594_
timestamp 1667941163
transform 1 0 21804 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0595_
timestamp 1667941163
transform 1 0 21344 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0596_
timestamp 1667941163
transform 1 0 25760 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0597_
timestamp 1667941163
transform 1 0 27140 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0598_
timestamp 1667941163
transform 1 0 24840 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0599_
timestamp 1667941163
transform 1 0 26036 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0600_
timestamp 1667941163
transform 1 0 27140 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0601_
timestamp 1667941163
transform 1 0 14260 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0602_
timestamp 1667941163
transform 1 0 22448 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0603_
timestamp 1667941163
transform 1 0 14260 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0604_
timestamp 1667941163
transform 1 0 14904 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0605_
timestamp 1667941163
transform 1 0 16284 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0606_
timestamp 1667941163
transform 1 0 19228 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0607_
timestamp 1667941163
transform 1 0 31372 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0608_
timestamp 1667941163
transform 1 0 31004 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0609_
timestamp 1667941163
transform 1 0 30820 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0610_
timestamp 1667941163
transform 1 0 20884 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0611_
timestamp 1667941163
transform 1 0 21252 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0612_
timestamp 1667941163
transform 1 0 20240 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0613_
timestamp 1667941163
transform 1 0 20608 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0614_
timestamp 1667941163
transform 1 0 21252 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0615_
timestamp 1667941163
transform 1 0 21620 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0616_
timestamp 1667941163
transform 1 0 28704 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0617_
timestamp 1667941163
transform 1 0 27600 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0618_
timestamp 1667941163
transform 1 0 28244 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0619_
timestamp 1667941163
transform 1 0 14260 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0620_
timestamp 1667941163
transform 1 0 16100 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0621_
timestamp 1667941163
transform 1 0 14352 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0622_
timestamp 1667941163
transform 1 0 14444 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0623_
timestamp 1667941163
transform 1 0 15088 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0624_
timestamp 1667941163
transform 1 0 14812 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0625_
timestamp 1667941163
transform 1 0 7820 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0626_
timestamp 1667941163
transform 1 0 11500 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0627_
timestamp 1667941163
transform 1 0 10948 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0628_
timestamp 1667941163
transform 1 0 23552 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0629_
timestamp 1667941163
transform 1 0 25208 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0630_
timestamp 1667941163
transform 1 0 24840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0631_
timestamp 1667941163
transform 1 0 25484 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0632_
timestamp 1667941163
transform 1 0 23276 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0633_
timestamp 1667941163
transform 1 0 23644 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0634_
timestamp 1667941163
transform 1 0 9108 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0635_
timestamp 1667941163
transform 1 0 6900 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0636_
timestamp 1667941163
transform 1 0 7636 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0637_
timestamp 1667941163
transform 1 0 27784 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0638_
timestamp 1667941163
transform 1 0 26496 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0639_
timestamp 1667941163
transform 1 0 26772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0640_
timestamp 1667941163
transform 1 0 27324 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0641_
timestamp 1667941163
transform 1 0 28244 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0642_
timestamp 1667941163
transform 1 0 29256 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0643_
timestamp 1667941163
transform 1 0 24656 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0644_
timestamp 1667941163
transform 1 0 25392 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0645_
timestamp 1667941163
transform 1 0 26036 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0646_
timestamp 1667941163
transform 1 0 11684 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0647_
timestamp 1667941163
transform 1 0 10120 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0648_
timestamp 1667941163
transform 1 0 10764 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0649_
timestamp 1667941163
transform 1 0 10028 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0650_
timestamp 1667941163
transform 1 0 9108 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0651_
timestamp 1667941163
transform 1 0 8924 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0652_
timestamp 1667941163
transform 1 0 8188 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0653_
timestamp 1667941163
transform 1 0 6532 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0654_
timestamp 1667941163
transform 1 0 7820 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0655_
timestamp 1667941163
transform 1 0 24564 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0656_
timestamp 1667941163
transform 1 0 21252 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0657_
timestamp 1667941163
transform 1 0 14352 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0658_
timestamp 1667941163
transform 1 0 13524 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0659_
timestamp 1667941163
transform 1 0 25668 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0660_
timestamp 1667941163
transform 1 0 26312 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0661_
timestamp 1667941163
transform 1 0 28796 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0662_
timestamp 1667941163
transform 1 0 33028 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0663_
timestamp 1667941163
transform 1 0 32384 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1667941163
transform 1 0 29164 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0665_
timestamp 1667941163
transform 1 0 29164 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0666_
timestamp 1667941163
transform 1 0 27140 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0667_
timestamp 1667941163
transform 1 0 27784 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0668_
timestamp 1667941163
transform 1 0 29808 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0669_
timestamp 1667941163
transform 1 0 30820 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0670_
timestamp 1667941163
transform 1 0 31924 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0671_
timestamp 1667941163
transform 1 0 31188 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0672_
timestamp 1667941163
transform 1 0 32292 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0673_
timestamp 1667941163
transform 1 0 25852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1667941163
transform 1 0 26588 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0675_
timestamp 1667941163
transform 1 0 26680 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0676_
timestamp 1667941163
transform 1 0 27140 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 1667941163
transform 1 0 11960 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0678_
timestamp 1667941163
transform 1 0 18492 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0679_
timestamp 1667941163
transform 1 0 18492 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0680_
timestamp 1667941163
transform 1 0 28796 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0681_
timestamp 1667941163
transform 1 0 28152 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1667941163
transform 1 0 3220 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0683_
timestamp 1667941163
transform 1 0 10948 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0684_
timestamp 1667941163
transform 1 0 17848 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0685_
timestamp 1667941163
transform 1 0 17204 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0686_
timestamp 1667941163
transform 1 0 17112 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0687_
timestamp 1667941163
transform 1 0 2300 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0688_
timestamp 1667941163
transform 1 0 2116 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1667941163
transform 1 0 34868 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0690_
timestamp 1667941163
transform 1 0 18124 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1667941163
transform 1 0 1840 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0692_
timestamp 1667941163
transform 1 0 1932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1667941163
transform 1 0 32384 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0694_
timestamp 1667941163
transform 1 0 28428 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0695_
timestamp 1667941163
transform 1 0 1840 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0696_
timestamp 1667941163
transform 1 0 30360 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0697_
timestamp 1667941163
transform 1 0 33304 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0698_
timestamp 1667941163
transform 1 0 28060 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1667941163
transform 1 0 28704 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0700_
timestamp 1667941163
transform 1 0 11132 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0701_
timestamp 1667941163
transform 1 0 5704 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0702_
timestamp 1667941163
transform 1 0 30176 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0703_
timestamp 1667941163
transform 1 0 27232 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0704_
timestamp 1667941163
transform 1 0 8924 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1667941163
transform 1 0 25116 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0706_
timestamp 1667941163
transform 1 0 32844 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0707_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1840 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0708_
timestamp 1667941163
transform 1 0 1932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0709_
timestamp 1667941163
transform 1 0 31096 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0710_
timestamp 1667941163
transform 1 0 14996 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0711_
timestamp 1667941163
transform 1 0 6256 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0712_
timestamp 1667941163
transform 1 0 21068 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1667941163
transform 1 0 5060 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0714_
timestamp 1667941163
transform 1 0 28244 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1667941163
transform 1 0 6164 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1667941163
transform 1 0 33396 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1667941163
transform 1 0 31280 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1667941163
transform 1 0 26588 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0719_
timestamp 1667941163
transform 1 0 4140 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1667941163
transform 1 0 2392 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1667941163
transform 1 0 3128 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0722_
timestamp 1667941163
transform 1 0 27232 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0723_
timestamp 1667941163
transform 1 0 32200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0724_
timestamp 1667941163
transform 1 0 2024 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0725_
timestamp 1667941163
transform 1 0 17940 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1667941163
transform 1 0 28428 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1667941163
transform 1 0 31004 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1667941163
transform 1 0 24748 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0729_
timestamp 1667941163
transform 1 0 28796 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1667941163
transform 1 0 4876 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1667941163
transform 1 0 1840 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1667941163
transform 1 0 19044 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0733_
timestamp 1667941163
transform 1 0 5336 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1667941163
transform 1 0 28980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1667941163
transform 1 0 28796 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0736_
timestamp 1667941163
transform 1 0 8280 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1667941163
transform 1 0 7636 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1667941163
transform 1 0 30544 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1667941163
transform 1 0 22908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0740_
timestamp 1667941163
transform 1 0 30452 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1667941163
transform 1 0 14168 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1667941163
transform 1 0 29900 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1667941163
transform 1 0 2760 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1667941163
transform 1 0 5336 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1667941163
transform 1 0 28888 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1667941163
transform 1 0 10672 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1667941163
transform 1 0 19872 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1667941163
transform 1 0 31648 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1667941163
transform 1 0 31372 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1667941163
transform 1 0 28796 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1667941163
transform 1 0 7176 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1667941163
transform 1 0 33304 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0753_
timestamp 1667941163
transform 1 0 6900 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1667941163
transform 1 0 1840 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0755_
timestamp 1667941163
transform 1 0 17296 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0756_
timestamp 1667941163
transform 1 0 30912 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1667941163
transform 1 0 14812 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 1667941163
transform 1 0 32752 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0759_
timestamp 1667941163
transform 1 0 25852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0760_
timestamp 1667941163
transform 1 0 25852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1667941163
transform 1 0 23920 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0762_
timestamp 1667941163
transform 1 0 27968 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1667941163
transform 1 0 30360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 1667941163
transform 1 0 7544 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1667941163
transform 1 0 25944 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0766_
timestamp 1667941163
transform 1 0 12420 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1667941163
transform 1 0 23092 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1667941163
transform 1 0 30820 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0769_
timestamp 1667941163
transform 1 0 9108 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1667941163
transform 1 0 30636 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1667941163
transform 1 0 28336 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1667941163
transform 1 0 16836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1667941163
transform 1 0 1932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1667941163
transform 1 0 21988 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0775_
timestamp 1667941163
transform 1 0 2300 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1667941163
transform 1 0 29716 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 1667941163
transform 1 0 25024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1667941163
transform 1 0 23184 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1667941163
transform 1 0 10488 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0780_
timestamp 1667941163
transform 1 0 22172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1667941163
transform 1 0 16836 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1667941163
transform 1 0 5060 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0783_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 22448 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0784_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 22356 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0785_
timestamp 1667941163
transform 1 0 10304 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0786_
timestamp 1667941163
transform 1 0 6532 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1667941163
transform 1 0 20516 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 1667941163
transform 1 0 21160 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1667941163
transform 1 0 23460 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0790_
timestamp 1667941163
transform 1 0 21252 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0791_
timestamp 1667941163
transform 1 0 20884 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 1667941163
transform 1 0 21252 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1667941163
transform 1 0 3864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0794_
timestamp 1667941163
transform 1 0 8004 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0795_
timestamp 1667941163
transform 1 0 21988 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1667941163
transform 1 0 22632 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0797_
timestamp 1667941163
transform 1 0 22908 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1667941163
transform 1 0 21988 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0799_
timestamp 1667941163
transform 1 0 22632 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1667941163
transform 1 0 22540 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1667941163
transform 1 0 22356 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0802_
timestamp 1667941163
transform 1 0 21804 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0803_
timestamp 1667941163
transform 1 0 21160 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0804_
timestamp 1667941163
transform 1 0 21988 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0805_
timestamp 1667941163
transform 1 0 21068 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0806_
timestamp 1667941163
transform 1 0 20792 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0807_
timestamp 1667941163
transform 1 0 19872 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1667941163
transform 1 0 20148 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0809_
timestamp 1667941163
transform 1 0 11316 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0810_
timestamp 1667941163
transform 1 0 21988 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0811_
timestamp 1667941163
transform 1 0 20424 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1667941163
transform 1 0 14996 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0813_
timestamp 1667941163
transform 1 0 10488 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0814_
timestamp 1667941163
transform 1 0 20056 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0815_
timestamp 1667941163
transform 1 0 21068 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1667941163
transform 1 0 21988 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0817_
timestamp 1667941163
transform 1 0 21528 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0818_
timestamp 1667941163
transform 1 0 17848 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1667941163
transform 1 0 20332 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1667941163
transform 1 0 21988 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0821_
timestamp 1667941163
transform 1 0 21436 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1667941163
transform 1 0 21620 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0823_
timestamp 1667941163
transform 1 0 21252 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0824_
timestamp 1667941163
transform 1 0 20516 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0825_
timestamp 1667941163
transform 1 0 22356 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0826_
timestamp 1667941163
transform 1 0 20608 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0827_
timestamp 1667941163
transform 1 0 21712 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0828_
timestamp 1667941163
transform 1 0 22540 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0829_
timestamp 1667941163
transform 1 0 21988 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1667941163
transform 1 0 14260 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1667941163
transform 1 0 21160 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0832_
timestamp 1667941163
transform 1 0 22632 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1667941163
transform 1 0 21988 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1667941163
transform 1 0 21344 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1667941163
transform 1 0 21712 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1667941163
transform 1 0 21068 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1667941163
transform 1 0 21252 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0838_
timestamp 1667941163
transform 1 0 22632 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0839_
timestamp 1667941163
transform 1 0 22356 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0840_
timestamp 1667941163
transform 1 0 23460 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1667941163
transform 1 0 23276 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1667941163
transform 1 0 23552 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0843_
timestamp 1667941163
transform 1 0 23460 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0844_
timestamp 1667941163
transform 1 0 20516 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0845_
timestamp 1667941163
transform 1 0 17480 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0846_
timestamp 1667941163
transform 1 0 18676 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0847_
timestamp 1667941163
transform 1 0 20424 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0848_
timestamp 1667941163
transform 1 0 23276 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0849_
timestamp 1667941163
transform 1 0 24564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0850_
timestamp 1667941163
transform 1 0 22540 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0851_
timestamp 1667941163
transform 1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0852_
timestamp 1667941163
transform 1 0 21988 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0853_
timestamp 1667941163
transform 1 0 22172 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0854_
timestamp 1667941163
transform 1 0 22264 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0855_
timestamp 1667941163
transform 1 0 19872 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0856_
timestamp 1667941163
transform 1 0 24196 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0857_
timestamp 1667941163
transform 1 0 17756 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0858_
timestamp 1667941163
transform 1 0 17112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0859_
timestamp 1667941163
transform 1 0 16836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0860_
timestamp 1667941163
transform 1 0 18124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0861_
timestamp 1667941163
transform 1 0 21344 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0862_
timestamp 1667941163
transform 1 0 22080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0863_
timestamp 1667941163
transform 1 0 21160 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0864_
timestamp 1667941163
transform 1 0 20976 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _0865_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14260 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0866_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 8648 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0867_
timestamp 1667941163
transform 1 0 4968 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0868_
timestamp 1667941163
transform 1 0 9108 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0869_
timestamp 1667941163
transform 1 0 9844 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0870_
timestamp 1667941163
transform 1 0 17940 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0871_
timestamp 1667941163
transform 1 0 14444 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0872_
timestamp 1667941163
transform 1 0 12236 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0873_
timestamp 1667941163
transform 1 0 9568 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0874_
timestamp 1667941163
transform 1 0 3496 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0875_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 12604 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0876_
timestamp 1667941163
transform 1 0 7636 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0877_
timestamp 1667941163
transform 1 0 3956 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0878_
timestamp 1667941163
transform 1 0 14260 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0879_
timestamp 1667941163
transform 1 0 4508 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0880_
timestamp 1667941163
transform 1 0 4048 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0881_
timestamp 1667941163
transform 1 0 15824 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0882_
timestamp 1667941163
transform 1 0 15272 0 1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0883_
timestamp 1667941163
transform 1 0 8188 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0884_
timestamp 1667941163
transform 1 0 18308 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0885_
timestamp 1667941163
transform 1 0 18032 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0886_
timestamp 1667941163
transform 1 0 14076 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0887_
timestamp 1667941163
transform 1 0 11684 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0888_
timestamp 1667941163
transform 1 0 3680 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0889_
timestamp 1667941163
transform 1 0 14260 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0890_
timestamp 1667941163
transform 1 0 9108 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0891_
timestamp 1667941163
transform 1 0 4232 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0892_
timestamp 1667941163
transform 1 0 16100 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0893_
timestamp 1667941163
transform 1 0 14444 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0894_
timestamp 1667941163
transform 1 0 11316 0 1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0895_
timestamp 1667941163
transform 1 0 3588 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0896_
timestamp 1667941163
transform 1 0 18124 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0897_
timestamp 1667941163
transform 1 0 3956 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0898_
timestamp 1667941163
transform 1 0 3956 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0899_
timestamp 1667941163
transform 1 0 11132 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0900_
timestamp 1667941163
transform 1 0 3956 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0901_
timestamp 1667941163
transform 1 0 17112 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0902_
timestamp 1667941163
transform 1 0 18216 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0903_
timestamp 1667941163
transform 1 0 12144 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0904_
timestamp 1667941163
transform 1 0 16560 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0905_
timestamp 1667941163
transform 1 0 9200 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0906_
timestamp 1667941163
transform 1 0 3956 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0907_
timestamp 1667941163
transform 1 0 6716 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0908_
timestamp 1667941163
transform 1 0 3956 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0909_
timestamp 1667941163
transform 1 0 14260 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0910_
timestamp 1667941163
transform 1 0 8740 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0911_
timestamp 1667941163
transform 1 0 11040 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0912_
timestamp 1667941163
transform 1 0 9108 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0913_
timestamp 1667941163
transform 1 0 6532 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0914_
timestamp 1667941163
transform 1 0 3956 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0915_
timestamp 1667941163
transform 1 0 18216 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0916_
timestamp 1667941163
transform 1 0 17940 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0917_
timestamp 1667941163
transform 1 0 19412 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0918_
timestamp 1667941163
transform 1 0 13984 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0919_
timestamp 1667941163
transform 1 0 6072 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0920_
timestamp 1667941163
transform 1 0 12696 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0921_
timestamp 1667941163
transform 1 0 13984 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0922_
timestamp 1667941163
transform 1 0 7544 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0923_
timestamp 1667941163
transform 1 0 4140 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0924_
timestamp 1667941163
transform 1 0 3680 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0925_
timestamp 1667941163
transform 1 0 16836 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0926_
timestamp 1667941163
transform 1 0 17388 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0927_
timestamp 1667941163
transform 1 0 18400 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0928_
timestamp 1667941163
transform 1 0 13524 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0929_
timestamp 1667941163
transform 1 0 3956 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0930_
timestamp 1667941163
transform 1 0 8648 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0931_
timestamp 1667941163
transform 1 0 17756 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0932_
timestamp 1667941163
transform 1 0 11684 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0933_
timestamp 1667941163
transform 1 0 6900 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0934_
timestamp 1667941163
transform 1 0 18860 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0935_
timestamp 1667941163
transform 1 0 11408 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0936_
timestamp 1667941163
transform 1 0 10488 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0937_
timestamp 1667941163
transform 1 0 7360 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0938_
timestamp 1667941163
transform 1 0 6716 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _0976_
timestamp 1667941163
transform 1 0 33304 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0977_
timestamp 1667941163
transform 1 0 7544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0978_
timestamp 1667941163
transform 1 0 27876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0979_
timestamp 1667941163
transform 1 0 14260 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0980_
timestamp 1667941163
transform 1 0 16836 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0981_
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0982_
timestamp 1667941163
transform 1 0 33764 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0983_
timestamp 1667941163
transform 1 0 18032 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0984_
timestamp 1667941163
transform 1 0 33396 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0985_
timestamp 1667941163
transform 1 0 7084 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0986_
timestamp 1667941163
transform 1 0 20792 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0987_
timestamp 1667941163
transform 1 0 31464 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0988_
timestamp 1667941163
transform 1 0 35420 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0989_
timestamp 1667941163
transform 1 0 31004 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0990_
timestamp 1667941163
transform 1 0 11684 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0991_
timestamp 1667941163
transform 1 0 28612 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0992_
timestamp 1667941163
transform 1 0 31280 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0993_
timestamp 1667941163
transform 1 0 30360 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0994_
timestamp 1667941163
transform 1 0 1748 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0995_
timestamp 1667941163
transform 1 0 1748 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0996_
timestamp 1667941163
transform 1 0 17480 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0997_
timestamp 1667941163
transform 1 0 9936 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0998_
timestamp 1667941163
transform 1 0 26404 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0999_
timestamp 1667941163
transform 1 0 2300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1000_
timestamp 1667941163
transform 1 0 16928 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1001_
timestamp 1667941163
transform 1 0 7084 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1002_
timestamp 1667941163
transform 1 0 11868 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1003_
timestamp 1667941163
transform 1 0 26772 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1004_
timestamp 1667941163
transform 1 0 6992 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1005_
timestamp 1667941163
transform 1 0 32292 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1006_
timestamp 1667941163
transform 1 0 32752 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1007_
timestamp 1667941163
transform 1 0 18492 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1008_
timestamp 1667941163
transform 1 0 25944 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1009_
timestamp 1667941163
transform 1 0 32384 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1010_
timestamp 1667941163
transform 1 0 2760 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1011_
timestamp 1667941163
transform 1 0 3128 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1012_
timestamp 1667941163
transform 1 0 4140 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1013_
timestamp 1667941163
transform 1 0 32292 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1014_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6624 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1015_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3956 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1015__100 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3220 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1016_
timestamp 1667941163
transform 1 0 17020 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1017_
timestamp 1667941163
transform 1 0 10396 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1018_
timestamp 1667941163
transform 1 0 17756 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1019_
timestamp 1667941163
transform 1 0 2392 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1020_
timestamp 1667941163
transform 1 0 26128 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1021_
timestamp 1667941163
transform 1 0 18492 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1021__101
timestamp 1667941163
transform 1 0 18676 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1022_
timestamp 1667941163
transform 1 0 24656 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1023_
timestamp 1667941163
transform 1 0 25852 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1024_
timestamp 1667941163
transform 1 0 11776 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1025_
timestamp 1667941163
transform 1 0 25944 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1026_
timestamp 1667941163
transform 1 0 30452 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1027__102
timestamp 1667941163
transform 1 0 30452 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1027_
timestamp 1667941163
transform 1 0 31096 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1028_
timestamp 1667941163
transform 1 0 28244 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1029_
timestamp 1667941163
transform 1 0 29716 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1030_
timestamp 1667941163
transform 1 0 31740 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1031_
timestamp 1667941163
transform 1 0 29716 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1032_
timestamp 1667941163
transform 1 0 25576 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1033__103
timestamp 1667941163
transform 1 0 31924 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1033_
timestamp 1667941163
transform 1 0 32292 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1034_
timestamp 1667941163
transform 1 0 13156 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1035_
timestamp 1667941163
transform 1 0 25300 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1036_
timestamp 1667941163
transform 1 0 28980 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1037_
timestamp 1667941163
transform 1 0 21988 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1038_
timestamp 1667941163
transform 1 0 9108 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1039__104
timestamp 1667941163
transform 1 0 7268 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1039_
timestamp 1667941163
transform 1 0 7268 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1040_
timestamp 1667941163
transform 1 0 9844 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1041_
timestamp 1667941163
transform 1 0 10120 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1042_
timestamp 1667941163
transform 1 0 7084 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1043_
timestamp 1667941163
transform 1 0 11224 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1044_
timestamp 1667941163
transform 1 0 28060 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1045_
timestamp 1667941163
transform 1 0 25668 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1045__105
timestamp 1667941163
transform 1 0 25852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1046_
timestamp 1667941163
transform 1 0 27140 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1047_
timestamp 1667941163
transform 1 0 28244 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1048_
timestamp 1667941163
transform 1 0 24932 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1049_
timestamp 1667941163
transform 1 0 26956 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1050_
timestamp 1667941163
transform 1 0 23184 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1051__106
timestamp 1667941163
transform 1 0 9200 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1051_
timestamp 1667941163
transform 1 0 9108 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1052_
timestamp 1667941163
transform 1 0 22816 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1053_
timestamp 1667941163
transform 1 0 23276 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1054_
timestamp 1667941163
transform 1 0 5888 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1055_
timestamp 1667941163
transform 1 0 23828 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1056_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14260 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _1057_
timestamp 1667941163
transform 1 0 10488 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1057__107
timestamp 1667941163
transform 1 0 10488 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1058_
timestamp 1667941163
transform 1 0 15180 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1059_
timestamp 1667941163
transform 1 0 17112 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _1060_
timestamp 1667941163
transform 1 0 7544 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1061_
timestamp 1667941163
transform 1 0 16836 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1062_
timestamp 1667941163
transform 1 0 21896 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1063__108
timestamp 1667941163
transform 1 0 28060 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1063_
timestamp 1667941163
transform 1 0 28060 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1064_
timestamp 1667941163
transform 1 0 20148 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1065_
timestamp 1667941163
transform 1 0 21988 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1066_
timestamp 1667941163
transform 1 0 28428 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1067_
timestamp 1667941163
transform 1 0 20792 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1068_
timestamp 1667941163
transform 1 0 20608 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1069__109
timestamp 1667941163
transform 1 0 30176 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1069_
timestamp 1667941163
transform 1 0 30176 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1070_
timestamp 1667941163
transform 1 0 16376 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1071_
timestamp 1667941163
transform 1 0 13984 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1072_
timestamp 1667941163
transform 1 0 30176 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1073_
timestamp 1667941163
transform 1 0 21988 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1074_
timestamp 1667941163
transform 1 0 25392 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1075_
timestamp 1667941163
transform 1 0 25024 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1075__110
timestamp 1667941163
transform 1 0 25116 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1076_
timestamp 1667941163
transform 1 0 20516 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1077_
timestamp 1667941163
transform 1 0 24472 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1078_
timestamp 1667941163
transform 1 0 24564 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1079_
timestamp 1667941163
transform 1 0 24564 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1080_
timestamp 1667941163
transform 1 0 6900 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1081__111
timestamp 1667941163
transform 1 0 10212 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1081_
timestamp 1667941163
transform 1 0 10120 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1082_
timestamp 1667941163
transform 1 0 4232 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1083_
timestamp 1667941163
transform 1 0 4968 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1084_
timestamp 1667941163
transform 1 0 13248 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1085_
timestamp 1667941163
transform 1 0 2760 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1086_
timestamp 1667941163
transform 1 0 28244 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1087__112
timestamp 1667941163
transform 1 0 29072 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1087_
timestamp 1667941163
transform 1 0 27968 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1088_
timestamp 1667941163
transform 1 0 30636 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1089_
timestamp 1667941163
transform 1 0 27140 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1090_
timestamp 1667941163
transform 1 0 27324 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1091_
timestamp 1667941163
transform 1 0 30452 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1092_
timestamp 1667941163
transform 1 0 12696 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1093_
timestamp 1667941163
transform 1 0 12144 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1093__113
timestamp 1667941163
transform 1 0 12144 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1094_
timestamp 1667941163
transform 1 0 24104 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1095_
timestamp 1667941163
transform 1 0 11868 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1096_
timestamp 1667941163
transform 1 0 12972 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1097_
timestamp 1667941163
transform 1 0 17388 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1098_
timestamp 1667941163
transform 1 0 27416 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1099__114
timestamp 1667941163
transform 1 0 26404 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1099_
timestamp 1667941163
transform 1 0 25944 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1100_
timestamp 1667941163
transform 1 0 24840 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1101_
timestamp 1667941163
transform 1 0 26404 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1102_
timestamp 1667941163
transform 1 0 27140 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1103_
timestamp 1667941163
transform 1 0 29440 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1104_
timestamp 1667941163
transform 1 0 15364 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1105__115
timestamp 1667941163
transform 1 0 12788 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1105_
timestamp 1667941163
transform 1 0 12696 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1106_
timestamp 1667941163
transform 1 0 22448 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1107_
timestamp 1667941163
transform 1 0 16836 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1108_
timestamp 1667941163
transform 1 0 15824 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1109_
timestamp 1667941163
transform 1 0 8648 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1110_
timestamp 1667941163
transform 1 0 24564 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1111__116
timestamp 1667941163
transform 1 0 26496 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1111_
timestamp 1667941163
transform 1 0 27140 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1112_
timestamp 1667941163
transform 1 0 10672 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1113_
timestamp 1667941163
transform 1 0 8280 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _1114_
timestamp 1667941163
transform 1 0 24656 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1115_
timestamp 1667941163
transform 1 0 6900 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1116_
timestamp 1667941163
transform 1 0 20792 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1117__117
timestamp 1667941163
transform 1 0 16100 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1117_
timestamp 1667941163
transform 1 0 16468 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1118_
timestamp 1667941163
transform 1 0 24564 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1119_
timestamp 1667941163
transform 1 0 23460 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1120_
timestamp 1667941163
transform 1 0 14720 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1121_
timestamp 1667941163
transform 1 0 23460 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1122_
timestamp 1667941163
transform 1 0 29808 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1123_
timestamp 1667941163
transform 1 0 29808 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1123__118
timestamp 1667941163
transform 1 0 29900 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1124_
timestamp 1667941163
transform 1 0 14720 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1125_
timestamp 1667941163
transform 1 0 28612 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1126_
timestamp 1667941163
transform 1 0 28060 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1127_
timestamp 1667941163
transform 1 0 24564 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1128_
timestamp 1667941163
transform 1 0 14628 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1129__119
timestamp 1667941163
transform 1 0 20148 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1129_
timestamp 1667941163
transform 1 0 19504 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1130_
timestamp 1667941163
transform 1 0 23368 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1131_
timestamp 1667941163
transform 1 0 14444 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1132_
timestamp 1667941163
transform 1 0 19688 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1133_
timestamp 1667941163
transform 1 0 23184 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1134_
timestamp 1667941163
transform 1 0 9660 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1135_
timestamp 1667941163
transform 1 0 12512 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1135__120
timestamp 1667941163
transform 1 0 11868 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1136_
timestamp 1667941163
transform 1 0 17756 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1137_
timestamp 1667941163
transform 1 0 8004 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1138_
timestamp 1667941163
transform 1 0 15640 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1139_
timestamp 1667941163
transform 1 0 5244 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1140__121
timestamp 1667941163
transform 1 0 23092 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1140_
timestamp 1667941163
transform 1 0 22908 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1141_
timestamp 1667941163
transform 1 0 11684 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1142_
timestamp 1667941163
transform 1 0 19412 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1143_
timestamp 1667941163
transform 1 0 16744 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1144__122
timestamp 1667941163
transform 1 0 19872 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1144_
timestamp 1667941163
transform 1 0 19504 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1145_
timestamp 1667941163
transform 1 0 30360 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1146_
timestamp 1667941163
transform 1 0 22448 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1147_
timestamp 1667941163
transform 1 0 30452 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1148_
timestamp 1667941163
transform 1 0 30728 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1148__123
timestamp 1667941163
transform 1 0 30912 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1149_
timestamp 1667941163
transform 1 0 8832 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1150_
timestamp 1667941163
transform 1 0 27140 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1151_
timestamp 1667941163
transform 1 0 19504 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1152__124
timestamp 1667941163
transform 1 0 32292 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1152_
timestamp 1667941163
transform 1 0 32292 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1153_
timestamp 1667941163
transform 1 0 5244 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1154_
timestamp 1667941163
transform 1 0 13984 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1155_
timestamp 1667941163
transform 1 0 5704 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1156_
timestamp 1667941163
transform 1 0 18032 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1156__125
timestamp 1667941163
transform 1 0 18124 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1157_
timestamp 1667941163
transform 1 0 29808 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1158_
timestamp 1667941163
transform 1 0 18124 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1159_
timestamp 1667941163
transform 1 0 22172 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1160__126
timestamp 1667941163
transform 1 0 14536 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1160_
timestamp 1667941163
transform 1 0 14352 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1161_
timestamp 1667941163
transform 1 0 31188 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1162_
timestamp 1667941163
transform 1 0 17296 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1163_
timestamp 1667941163
transform 1 0 27600 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1164__127
timestamp 1667941163
transform 1 0 30728 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1164_
timestamp 1667941163
transform 1 0 29808 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1165_
timestamp 1667941163
transform 1 0 25484 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1166_
timestamp 1667941163
transform 1 0 28612 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1167_
timestamp 1667941163
transform 1 0 22356 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1168__128
timestamp 1667941163
transform 1 0 25208 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1168_
timestamp 1667941163
transform 1 0 23368 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1169_
timestamp 1667941163
transform 1 0 27876 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1170_
timestamp 1667941163
transform 1 0 25208 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1171_
timestamp 1667941163
transform 1 0 17940 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1172_
timestamp 1667941163
transform 1 0 28336 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1172__129
timestamp 1667941163
transform 1 0 28152 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1173_
timestamp 1667941163
transform 1 0 19688 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1174_
timestamp 1667941163
transform 1 0 25116 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1175_
timestamp 1667941163
transform 1 0 8556 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1176__130
timestamp 1667941163
transform 1 0 12696 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1176_
timestamp 1667941163
transform 1 0 12604 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1177_
timestamp 1667941163
transform 1 0 19688 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1178_
timestamp 1667941163
transform 1 0 12696 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1179_
timestamp 1667941163
transform 1 0 20700 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1180__131
timestamp 1667941163
transform 1 0 7912 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1180_
timestamp 1667941163
transform 1 0 7820 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1181_
timestamp 1667941163
transform 1 0 26772 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1182_
timestamp 1667941163
transform 1 0 14996 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1183_
timestamp 1667941163
transform 1 0 29164 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1184__132
timestamp 1667941163
transform 1 0 20976 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1184_
timestamp 1667941163
transform 1 0 20792 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1185_
timestamp 1667941163
transform 1 0 11776 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1186_
timestamp 1667941163
transform 1 0 23460 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1187_
timestamp 1667941163
transform 1 0 6440 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1188__133
timestamp 1667941163
transform 1 0 6808 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1188_
timestamp 1667941163
transform 1 0 6624 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1189_
timestamp 1667941163
transform 1 0 28336 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1190_
timestamp 1667941163
transform 1 0 21988 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1191_
timestamp 1667941163
transform 1 0 28980 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1192__134
timestamp 1667941163
transform 1 0 28520 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1192_
timestamp 1667941163
transform 1 0 27140 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1193_
timestamp 1667941163
transform 1 0 11684 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1194_
timestamp 1667941163
transform 1 0 23920 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1195_
timestamp 1667941163
transform 1 0 23276 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1196_
timestamp 1667941163
transform 1 0 11684 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1196__135
timestamp 1667941163
transform 1 0 11500 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1197_
timestamp 1667941163
transform 1 0 23000 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1198_
timestamp 1667941163
transform 1 0 10396 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1199_
timestamp 1667941163
transform 1 0 21988 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1200_
timestamp 1667941163
transform 1 0 11776 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1200__136
timestamp 1667941163
transform 1 0 11868 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1201_
timestamp 1667941163
transform 1 0 8004 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1202_
timestamp 1667941163
transform 1 0 9936 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1203_
timestamp 1667941163
transform 1 0 7084 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1667941163
transform 1 0 38088 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1667941163
transform 1 0 38088 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1667941163
transform 1 0 22724 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37444 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1667941163
transform 1 0 1564 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1667941163
transform 1 0 34868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1667941163
transform 1 0 2300 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1667941163
transform 1 0 38088 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1667941163
transform 1 0 31004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1667941163
transform 1 0 2576 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1667941163
transform 1 0 1564 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1667941163
transform 1 0 2944 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1667941163
transform 1 0 3220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1667941163
transform 1 0 1564 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1667941163
transform 1 0 1564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1667941163
transform 1 0 38088 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1667941163
transform 1 0 18124 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1667941163
transform 1 0 33672 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1667941163
transform 1 0 1564 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1667941163
transform 1 0 1564 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1667941163
transform 1 0 1564 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1667941163
transform 1 0 23552 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1667941163
transform 1 0 14904 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1667941163
transform 1 0 36708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1667941163
transform 1 0 1564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1667941163
transform 1 0 38088 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1667941163
transform 1 0 24564 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1667941163
transform 1 0 14260 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1667941163
transform 1 0 36708 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1667941163
transform 1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1667941163
transform 1 0 38088 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1667941163
transform 1 0 1564 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1667941163
transform 1 0 1564 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1667941163
transform 1 0 25852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1667941163
transform 1 0 1564 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1667941163
transform 1 0 33028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1667941163
transform 1 0 33580 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1667941163
transform 1 0 1564 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1667941163
transform 1 0 2576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1667941163
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1667941163
transform 1 0 36156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1667941163
transform 1 0 38088 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1667941163
transform 1 0 38088 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1667941163
transform 1 0 1564 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1667941163
transform 1 0 1564 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1667941163
transform 1 0 38088 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1667941163
transform 1 0 4600 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1667941163
transform 1 0 38088 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1667941163
transform 1 0 38088 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50
timestamp 1667941163
transform 1 0 37444 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1667941163
transform 1 0 14260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1667941163
transform 1 0 1564 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1667941163
transform 1 0 38088 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1667941163
transform 1 0 21252 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1667941163
transform 1 0 32292 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1667941163
transform 1 0 30452 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1667941163
transform 1 0 3956 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1667941163
transform 1 0 9108 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1667941163
transform 1 0 29716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1667941163
transform 1 0 1564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output61 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 10396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1667941163
transform 1 0 1564 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1667941163
transform 1 0 37996 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1667941163
transform 1 0 15548 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1667941163
transform 1 0 37996 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1667941163
transform 1 0 37996 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1667941163
transform 1 0 16836 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1667941163
transform 1 0 10396 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1667941163
transform 1 0 27140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1667941163
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1667941163
transform 1 0 37996 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1667941163
transform 1 0 37996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1667941163
transform 1 0 37996 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1667941163
transform 1 0 29716 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1667941163
transform 1 0 12328 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1667941163
transform 1 0 37996 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1667941163
transform 1 0 37996 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1667941163
transform 1 0 36616 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1667941163
transform 1 0 21988 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1667941163
transform 1 0 1564 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1667941163
transform 1 0 32292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1667941163
transform 1 0 37996 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1667941163
transform 1 0 6532 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1667941163
transform 1 0 1564 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1667941163
transform 1 0 19412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1667941163
transform 1 0 1564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1667941163
transform 1 0 24564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1667941163
transform 1 0 7820 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1667941163
transform 1 0 20056 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1667941163
transform 1 0 1564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1667941163
transform 1 0 1564 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1667941163
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1667941163
transform 1 0 1564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1667941163
transform 1 0 34868 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1667941163
transform 1 0 27784 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1667941163
transform 1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1667941163
transform 1 0 37996 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1667941163
transform 1 0 37996 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1667941163
transform 1 0 1564 0 1 36992
box -38 -48 406 592
<< labels >>
flabel metal3 s 39200 6128 39800 6248 0 FreeSans 480 0 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 0 nsew signal input
flabel metal3 s 39200 33328 39800 33448 0 FreeSans 480 0 0 0 bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 1 nsew signal input
flabel metal2 s 22558 39200 22614 39800 0 FreeSans 224 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 2 nsew signal input
flabel metal3 s 39200 38088 39800 38208 0 FreeSans 480 0 0 0 bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 3 nsew signal input
flabel metal3 s 200 12248 800 12368 0 FreeSans 480 0 0 0 bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_
port 4 nsew signal input
flabel metal2 s 34794 200 34850 800 0 FreeSans 224 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_
port 5 nsew signal input
flabel metal3 s 200 36728 800 36848 0 FreeSans 480 0 0 0 bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_
port 6 nsew signal input
flabel metal2 s 38014 39200 38070 39800 0 FreeSans 224 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_
port 7 nsew signal input
flabel metal2 s 28998 200 29054 800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
port 8 nsew signal input
flabel metal3 s 200 7488 800 7608 0 FreeSans 480 0 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
port 9 nsew signal input
flabel metal3 s 200 30608 800 30728 0 FreeSans 480 0 0 0 ccff_head
port 10 nsew signal input
flabel metal2 s 10322 200 10378 800 0 FreeSans 224 90 0 0 ccff_tail
port 11 nsew signal tristate
flabel metal3 s 200 38088 800 38208 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 12 nsew signal input
flabel metal2 s 4526 200 4582 800 0 FreeSans 224 90 0 0 chanx_right_in[10]
port 13 nsew signal input
flabel metal3 s 200 20408 800 20528 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 14 nsew signal input
flabel metal3 s 200 17688 800 17808 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 15 nsew signal input
flabel metal3 s 39200 28568 39800 28688 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 16 nsew signal input
flabel metal2 s 18050 39200 18106 39800 0 FreeSans 224 90 0 0 chanx_right_in[14]
port 17 nsew signal input
flabel metal2 s 33506 200 33562 800 0 FreeSans 224 90 0 0 chanx_right_in[15]
port 18 nsew signal input
flabel metal3 s 200 25168 800 25288 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 19 nsew signal input
flabel metal3 s 200 31968 800 32088 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 20 nsew signal input
flabel metal3 s 200 27208 800 27328 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 21 nsew signal input
flabel metal2 s 22558 200 22614 800 0 FreeSans 224 90 0 0 chanx_right_in[1]
port 22 nsew signal input
flabel metal2 s 14830 200 14886 800 0 FreeSans 224 90 0 0 chanx_right_in[2]
port 23 nsew signal input
flabel metal2 s 39302 200 39358 800 0 FreeSans 224 90 0 0 chanx_right_in[3]
port 24 nsew signal input
flabel metal3 s 200 1368 800 1488 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 25 nsew signal input
flabel metal3 s 39200 20408 39800 20528 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 26 nsew signal input
flabel metal2 s 24490 39200 24546 39800 0 FreeSans 224 90 0 0 chanx_right_in[6]
port 27 nsew signal input
flabel metal2 s 13542 39200 13598 39800 0 FreeSans 224 90 0 0 chanx_right_in[7]
port 28 nsew signal input
flabel metal3 s 39200 36728 39800 36848 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 29 nsew signal input
flabel metal2 s 16762 200 16818 800 0 FreeSans 224 90 0 0 chanx_right_in[9]
port 30 nsew signal input
flabel metal3 s 200 15648 800 15768 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 31 nsew signal tristate
flabel metal3 s 39200 34688 39800 34808 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 32 nsew signal tristate
flabel metal2 s 15474 39200 15530 39800 0 FreeSans 224 90 0 0 chanx_right_out[11]
port 33 nsew signal tristate
flabel metal3 s 39200 8848 39800 8968 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 34 nsew signal tristate
flabel metal3 s 39200 12248 39800 12368 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 35 nsew signal tristate
flabel metal2 s 16762 39200 16818 39800 0 FreeSans 224 90 0 0 chanx_right_out[14]
port 36 nsew signal tristate
flabel metal2 s 10322 39200 10378 39800 0 FreeSans 224 90 0 0 chanx_right_out[15]
port 37 nsew signal tristate
flabel metal2 s 25778 200 25834 800 0 FreeSans 224 90 0 0 chanx_right_out[16]
port 38 nsew signal tristate
flabel metal2 s 9034 200 9090 800 0 FreeSans 224 90 0 0 chanx_right_out[17]
port 39 nsew signal tristate
flabel metal3 s 39200 29928 39800 30048 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 40 nsew signal tristate
flabel metal2 s 38014 200 38070 800 0 FreeSans 224 90 0 0 chanx_right_out[1]
port 41 nsew signal tristate
flabel metal3 s 39200 15648 39800 15768 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 42 nsew signal tristate
flabel metal2 s 28998 39200 29054 39800 0 FreeSans 224 90 0 0 chanx_right_out[3]
port 43 nsew signal tristate
flabel metal2 s 12254 39200 12310 39800 0 FreeSans 224 90 0 0 chanx_right_out[4]
port 44 nsew signal tristate
flabel metal3 s 39200 1368 39800 1488 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 45 nsew signal tristate
flabel metal3 s 39200 31968 39800 32088 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 46 nsew signal tristate
flabel metal2 s 36726 39200 36782 39800 0 FreeSans 224 90 0 0 chanx_right_out[7]
port 47 nsew signal tristate
flabel metal2 s 21270 39200 21326 39800 0 FreeSans 224 90 0 0 chanx_right_out[8]
port 48 nsew signal tristate
flabel metal3 s 200 19048 800 19168 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 49 nsew signal tristate
flabel metal3 s 39200 7488 39800 7608 0 FreeSans 480 0 0 0 chany_bottom_in[0]
port 50 nsew signal input
flabel metal3 s 200 22448 800 22568 0 FreeSans 480 0 0 0 chany_bottom_in[10]
port 51 nsew signal input
flabel metal3 s 200 2728 800 2848 0 FreeSans 480 0 0 0 chany_bottom_in[11]
port 52 nsew signal input
flabel metal2 s 25778 39200 25834 39800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 53 nsew signal input
flabel metal3 s 200 28568 800 28688 0 FreeSans 480 0 0 0 chany_bottom_in[13]
port 54 nsew signal input
flabel metal2 s 30286 200 30342 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 55 nsew signal input
flabel metal2 s 33506 39200 33562 39800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 56 nsew signal input
flabel metal3 s 200 9528 800 9648 0 FreeSans 480 0 0 0 chany_bottom_in[16]
port 57 nsew signal input
flabel metal2 s 2594 200 2650 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 58 nsew signal input
flabel metal2 s 11610 200 11666 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 59 nsew signal input
flabel metal2 s 36082 200 36138 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 60 nsew signal input
flabel metal3 s 39200 17008 39800 17128 0 FreeSans 480 0 0 0 chany_bottom_in[2]
port 61 nsew signal input
flabel metal3 s 39200 10888 39800 11008 0 FreeSans 480 0 0 0 chany_bottom_in[3]
port 62 nsew signal input
flabel metal3 s 200 6128 800 6248 0 FreeSans 480 0 0 0 chany_bottom_in[4]
port 63 nsew signal input
flabel metal3 s 200 33328 800 33448 0 FreeSans 480 0 0 0 chany_bottom_in[5]
port 64 nsew signal input
flabel metal3 s 39200 2728 39800 2848 0 FreeSans 480 0 0 0 chany_bottom_in[6]
port 65 nsew signal input
flabel metal2 s 4526 39200 4582 39800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 66 nsew signal input
flabel metal3 s 39200 14288 39800 14408 0 FreeSans 480 0 0 0 chany_bottom_in[8]
port 67 nsew signal input
flabel metal3 s 39200 25168 39800 25288 0 FreeSans 480 0 0 0 chany_bottom_in[9]
port 68 nsew signal input
flabel metal2 s 31574 200 31630 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 69 nsew signal tristate
flabel metal3 s 39200 27208 39800 27328 0 FreeSans 480 0 0 0 chany_bottom_out[10]
port 70 nsew signal tristate
flabel metal2 s 5814 39200 5870 39800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 71 nsew signal tristate
flabel metal3 s 200 23808 800 23928 0 FreeSans 480 0 0 0 chany_bottom_out[12]
port 72 nsew signal tristate
flabel metal2 s 19338 200 19394 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 73 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 74 nsew signal tristate
flabel metal2 s 23846 200 23902 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 75 nsew signal tristate
flabel metal2 s 7746 39200 7802 39800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 76 nsew signal tristate
flabel metal2 s 19982 39200 20038 39800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 77 nsew signal tristate
flabel metal3 s 200 4768 800 4888 0 FreeSans 480 0 0 0 chany_bottom_out[18]
port 78 nsew signal tristate
flabel metal2 s 18 39200 74 39800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 79 nsew signal tristate
flabel metal2 s 5814 200 5870 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 80 nsew signal tristate
flabel metal2 s 1306 200 1362 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 81 nsew signal tristate
flabel metal2 s 34794 39200 34850 39800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 82 nsew signal tristate
flabel metal2 s 27710 39200 27766 39800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 83 nsew signal tristate
flabel metal2 s 18050 200 18106 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 84 nsew signal tristate
flabel metal2 s 39302 39200 39358 39800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 85 nsew signal tristate
flabel metal3 s 39200 4088 39800 4208 0 FreeSans 480 0 0 0 chany_bottom_out[8]
port 86 nsew signal tristate
flabel metal2 s 1306 39200 1362 39800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 87 nsew signal tristate
flabel metal3 s 39200 21768 39800 21888 0 FreeSans 480 0 0 0 pReset
port 88 nsew signal input
flabel metal2 s 7102 200 7158 800 0 FreeSans 224 90 0 0 prog_clk
port 89 nsew signal input
flabel metal2 s 13542 200 13598 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 90 nsew signal input
flabel metal3 s 200 14288 800 14408 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 91 nsew signal input
flabel metal3 s 39200 23808 39800 23928 0 FreeSans 480 0 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 92 nsew signal input
flabel metal2 s 21270 200 21326 800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
port 93 nsew signal input
flabel metal2 s 32218 39200 32274 39800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
port 94 nsew signal input
flabel metal2 s 30286 39200 30342 39800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
port 95 nsew signal input
flabel metal2 s 3238 39200 3294 39800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_
port 96 nsew signal input
flabel metal2 s 9034 39200 9090 39800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_
port 97 nsew signal input
flabel metal2 s 27066 200 27122 800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_
port 98 nsew signal input
flabel metal3 s 200 10888 800 11008 0 FreeSans 480 0 0 0 right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_
port 99 nsew signal input
flabel metal3 s 200 35368 800 35488 0 FreeSans 480 0 0 0 vccd1
port 100 nsew signal bidirectional
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 100 nsew signal bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 100 nsew signal bidirectional
flabel metal3 s 39200 19048 39800 19168 0 FreeSans 480 0 0 0 vssd1
port 101 nsew signal bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 101 nsew signal bidirectional
rlabel metal1 19964 37536 19964 37536 0 vccd1
rlabel metal1 19964 36992 19964 36992 0 vssd1
rlabel metal2 20746 4369 20746 4369 0 _0000_
rlabel metal2 21574 8432 21574 8432 0 _0001_
rlabel metal1 12558 7895 12558 7895 0 _0002_
rlabel metal1 21114 3094 21114 3094 0 _0003_
rlabel metal1 20424 9622 20424 9622 0 _0004_
rlabel metal1 20891 11798 20891 11798 0 _0005_
rlabel metal1 20102 18598 20102 18598 0 _0006_
rlabel metal1 20976 8058 20976 8058 0 _0007_
rlabel metal2 17710 4505 17710 4505 0 _0008_
rlabel metal1 5382 12281 5382 12281 0 _0009_
rlabel metal1 21298 13804 21298 13804 0 _0010_
rlabel metal2 12742 13294 12742 13294 0 _0011_
rlabel metal1 17211 13294 17211 13294 0 _0012_
rlabel metal1 19412 10166 19412 10166 0 _0013_
rlabel metal1 13761 13226 13761 13226 0 _0014_
rlabel metal1 20286 13158 20286 13158 0 _0015_
rlabel metal1 21344 5338 21344 5338 0 _0016_
rlabel metal1 14214 5780 14214 5780 0 _0017_
rlabel metal1 19642 9513 19642 9513 0 _0018_
rlabel metal2 20654 5406 20654 5406 0 _0019_
rlabel metal2 23690 8024 23690 8024 0 _0020_
rlabel metal2 18170 9316 18170 9316 0 _0021_
rlabel metal2 16606 6664 16606 6664 0 _0022_
rlabel metal2 17618 4318 17618 4318 0 _0023_
rlabel metal1 18676 7718 18676 7718 0 _0024_
rlabel metal2 9338 8670 9338 8670 0 _0025_
rlabel metal2 17986 2346 17986 2346 0 _0026_
rlabel metal1 8786 5304 8786 5304 0 _0027_
rlabel metal1 21988 12070 21988 12070 0 _0028_
rlabel metal1 20523 12886 20523 12886 0 _0029_
rlabel metal1 21160 14586 21160 14586 0 _0030_
rlabel metal2 18538 14382 18538 14382 0 _0031_
rlabel metal1 7406 2414 7406 2414 0 _0032_
rlabel metal1 23138 6392 23138 6392 0 _0033_
rlabel metal1 18216 3706 18216 3706 0 _0034_
rlabel metal2 17250 3264 17250 3264 0 _0035_
rlabel metal1 14398 4760 14398 4760 0 _0036_
rlabel metal1 18945 3094 18945 3094 0 _0037_
rlabel metal1 21068 4726 21068 4726 0 _0038_
rlabel metal2 19366 4862 19366 4862 0 _0039_
rlabel metal1 21298 9656 21298 9656 0 _0040_
rlabel metal2 21114 8874 21114 8874 0 _0041_
rlabel metal1 13064 10166 13064 10166 0 _0042_
rlabel metal2 9430 14654 9430 14654 0 _0043_
rlabel metal1 7459 3502 7459 3502 0 _0044_
rlabel metal1 13386 2856 13386 2856 0 _0045_
rlabel metal1 22494 6664 22494 6664 0 _0046_
rlabel metal1 20431 7446 20431 7446 0 _0047_
rlabel metal1 20838 15878 20838 15878 0 _0048_
rlabel metal1 18354 13498 18354 13498 0 _0049_
rlabel metal1 7636 16966 7636 16966 0 _0050_
rlabel metal1 7360 18666 7360 18666 0 _0051_
rlabel metal2 14030 10438 14030 10438 0 _0052_
rlabel metal2 20746 14586 20746 14586 0 _0053_
rlabel metal1 18078 6188 18078 6188 0 _0054_
rlabel metal1 18630 7480 18630 7480 0 _0055_
rlabel metal1 20102 16150 20102 16150 0 _0056_
rlabel metal2 20746 11050 20746 11050 0 _0057_
rlabel metal1 19649 14314 19649 14314 0 _0058_
rlabel metal1 17671 15470 17671 15470 0 _0059_
rlabel metal1 14122 7412 14122 7412 0 _0060_
rlabel metal1 20930 14246 20930 14246 0 _0061_
rlabel metal2 20010 7395 20010 7395 0 _0062_
rlabel metal1 19182 2618 19182 2618 0 _0063_
rlabel metal1 11684 9010 11684 9010 0 _0064_
rlabel metal2 8142 8704 8142 8704 0 _0065_
rlabel metal1 18177 4522 18177 4522 0 _0066_
rlabel metal2 10534 9078 10534 9078 0 _0067_
rlabel metal1 9292 10778 9292 10778 0 _0068_
rlabel metal2 20194 4828 20194 4828 0 _0069_
rlabel metal1 19504 12614 19504 12614 0 _0070_
rlabel metal2 20838 14824 20838 14824 0 _0071_
rlabel metal1 17434 18326 17434 18326 0 _0072_
rlabel metal2 20470 15198 20470 15198 0 _0073_
rlabel metal2 8418 28220 8418 28220 0 _0074_
rlabel metal1 11914 30668 11914 30668 0 _0075_
rlabel metal1 25668 5338 25668 5338 0 _0076_
rlabel metal1 12190 20026 12190 20026 0 _0077_
rlabel metal1 12236 16762 12236 16762 0 _0078_
rlabel metal1 28336 2618 28336 2618 0 _0079_
rlabel metal1 29302 13294 29302 13294 0 _0080_
rlabel metal2 4738 16966 4738 16966 0 _0081_
rlabel metal1 9246 17850 9246 17850 0 _0082_
rlabel metal1 25438 7888 25438 7888 0 _0083_
rlabel metal2 27370 19788 27370 19788 0 _0084_
rlabel metal2 8694 21828 8694 21828 0 _0085_
rlabel metal1 19918 22746 19918 22746 0 _0086_
rlabel metal1 15640 28526 15640 28526 0 _0087_
rlabel metal2 18722 15402 18722 15402 0 _0088_
rlabel metal1 28106 5338 28106 5338 0 _0089_
rlabel metal2 5382 16966 5382 16966 0 _0090_
rlabel metal1 27186 4794 27186 4794 0 _0091_
rlabel metal1 25990 4080 25990 4080 0 _0092_
rlabel metal1 29486 4114 29486 4114 0 _0093_
rlabel metal2 31050 3332 31050 3332 0 _0094_
rlabel metal2 32154 12852 32154 12852 0 _0095_
rlabel metal1 16974 23290 16974 23290 0 _0096_
rlabel metal1 29578 16082 29578 16082 0 _0097_
rlabel metal1 19136 26010 19136 26010 0 _0098_
rlabel metal1 5934 16218 5934 16218 0 _0099_
rlabel metal2 29118 11322 29118 11322 0 _0100_
rlabel metal1 10442 24922 10442 24922 0 _0101_
rlabel metal1 29210 12682 29210 12682 0 _0102_
rlabel metal1 30498 7854 30498 7854 0 _0103_
rlabel metal1 20286 26010 20286 26010 0 _0104_
rlabel metal2 13662 25398 13662 25398 0 _0105_
rlabel metal1 24150 26996 24150 26996 0 _0106_
rlabel metal1 18492 22610 18492 22610 0 _0107_
rlabel metal1 9936 20026 9936 20026 0 _0108_
rlabel metal2 13294 22202 13294 22202 0 _0109_
rlabel metal1 25300 20570 25300 20570 0 _0110_
rlabel metal1 15962 31280 15962 31280 0 _0111_
rlabel metal1 19504 30362 19504 30362 0 _0112_
rlabel metal2 16974 23324 16974 23324 0 _0113_
rlabel metal2 30038 10234 30038 10234 0 _0114_
rlabel metal1 31510 19788 31510 19788 0 _0115_
rlabel metal1 24380 10234 24380 10234 0 _0116_
rlabel metal1 21022 26010 21022 26010 0 _0117_
rlabel metal2 17618 26758 17618 26758 0 _0118_
rlabel metal1 7866 17136 7866 17136 0 _0119_
rlabel metal1 23966 11152 23966 11152 0 _0120_
rlabel metal1 29348 8466 29348 8466 0 _0121_
rlabel metal1 20792 23290 20792 23290 0 _0122_
rlabel metal1 15686 25296 15686 25296 0 _0123_
rlabel metal1 12351 26350 12351 26350 0 _0124_
rlabel metal1 24334 28084 24334 28084 0 _0125_
rlabel metal2 26358 26180 26358 26180 0 _0126_
rlabel metal1 27370 27982 27370 27982 0 _0127_
rlabel metal1 22034 27064 22034 27064 0 _0128_
rlabel metal1 12006 19380 12006 19380 0 _0129_
rlabel metal1 13248 24174 13248 24174 0 _0130_
rlabel metal2 30038 6086 30038 6086 0 _0131_
rlabel metal2 28474 8636 28474 8636 0 _0132_
rlabel metal2 28474 18564 28474 18564 0 _0133_
rlabel metal2 5474 18598 5474 18598 0 _0134_
rlabel metal2 7038 21318 7038 21318 0 _0135_
rlabel metal1 11040 20570 11040 20570 0 _0136_
rlabel metal1 21712 17850 21712 17850 0 _0137_
rlabel metal2 27370 16252 27370 16252 0 _0138_
rlabel metal1 27370 15028 27370 15028 0 _0139_
rlabel metal1 14720 18938 14720 18938 0 _0140_
rlabel metal2 19458 19516 19458 19516 0 _0141_
rlabel metal2 31050 17850 31050 17850 0 _0142_
rlabel metal2 20286 21386 20286 21386 0 _0143_
rlabel metal2 21298 22916 21298 22916 0 _0144_
rlabel metal1 28474 20944 28474 20944 0 _0145_
rlabel metal2 14674 20604 14674 20604 0 _0146_
rlabel metal1 15088 22746 15088 22746 0 _0147_
rlabel metal2 11546 25670 11546 25670 0 _0148_
rlabel metal1 25714 15436 25714 15436 0 _0149_
rlabel metal2 23322 16388 23322 16388 0 _0150_
rlabel metal1 7866 17680 7866 17680 0 _0151_
rlabel metal1 27186 14586 27186 14586 0 _0152_
rlabel metal1 28888 14586 28888 14586 0 _0153_
rlabel metal1 26266 23120 26266 23120 0 _0154_
rlabel metal1 10534 26826 10534 26826 0 _0155_
rlabel metal2 9154 27132 9154 27132 0 _0156_
rlabel metal1 6578 27540 6578 27540 0 _0157_
rlabel metal2 14398 26180 14398 26180 0 _0158_
rlabel metal1 26542 20400 26542 20400 0 _0159_
rlabel metal1 33074 16490 33074 16490 0 _0160_
rlabel metal1 28014 22576 28014 22576 0 _0161_
rlabel metal1 30452 21658 30452 21658 0 _0162_
rlabel metal2 32522 23494 32522 23494 0 _0163_
rlabel metal2 27370 7548 27370 7548 0 _0164_
rlabel metal1 18630 16762 18630 16762 0 _0165_
rlabel metal1 28612 15470 28612 15470 0 _0166_
rlabel metal1 17296 18394 17296 18394 0 _0167_
rlabel metal2 2346 17204 2346 17204 0 _0168_
rlabel metal2 22034 8789 22034 8789 0 _0169_
rlabel metal1 20838 16082 20838 16082 0 _0170_
rlabel metal1 21114 14416 21114 14416 0 _0171_
rlabel metal2 20148 2652 20148 2652 0 _0172_
rlabel metal1 20746 18734 20746 18734 0 _0173_
rlabel metal1 21298 5236 21298 5236 0 _0174_
rlabel metal1 18400 7854 18400 7854 0 _0175_
rlabel metal1 21942 12818 21942 12818 0 _0176_
rlabel metal2 6854 14926 6854 14926 0 _0177_
rlabel metal1 2162 17748 2162 17748 0 _0178_
rlabel metal1 17204 19482 17204 19482 0 _0179_
rlabel metal1 11132 14586 11132 14586 0 _0180_
rlabel metal2 17986 17986 17986 17986 0 _0181_
rlabel metal2 3358 16830 3358 16830 0 _0182_
rlabel metal1 26910 13294 26910 13294 0 _0183_
rlabel metal1 18630 17306 18630 17306 0 _0184_
rlabel metal1 24886 7480 24886 7480 0 _0185_
rlabel metal1 26082 8058 26082 8058 0 _0186_
rlabel metal2 12006 8670 12006 8670 0 _0187_
rlabel metal2 26726 11764 26726 11764 0 _0188_
rlabel metal1 30774 22202 30774 22202 0 _0189_
rlabel metal1 32338 23596 32338 23596 0 _0190_
rlabel metal1 28106 22746 28106 22746 0 _0191_
rlabel metal2 29302 21828 29302 21828 0 _0192_
rlabel metal1 32016 24378 32016 24378 0 _0193_
rlabel metal1 29624 23154 29624 23154 0 _0194_
rlabel metal1 25852 19754 25852 19754 0 _0195_
rlabel metal1 32476 16762 32476 16762 0 _0196_
rlabel metal2 13570 26792 13570 26792 0 _0197_
rlabel metal1 25116 24038 25116 24038 0 _0198_
rlabel metal2 29210 11934 29210 11934 0 _0199_
rlabel metal2 22218 24344 22218 24344 0 _0200_
rlabel metal2 9338 26588 9338 26588 0 _0201_
rlabel metal1 7682 25874 7682 25874 0 _0202_
rlabel metal2 10074 28220 10074 28220 0 _0203_
rlabel metal1 11822 27064 11822 27064 0 _0204_
rlabel metal1 7820 26894 7820 26894 0 _0205_
rlabel metal1 10856 27098 10856 27098 0 _0206_
rlabel metal1 28290 15096 28290 15096 0 _0207_
rlabel metal2 25898 22814 25898 22814 0 _0208_
rlabel metal2 27370 14620 27370 14620 0 _0209_
rlabel metal1 28198 12954 28198 12954 0 _0210_
rlabel metal1 24978 24378 24978 24378 0 _0211_
rlabel metal1 26910 22202 26910 22202 0 _0212_
rlabel metal2 23690 17000 23690 17000 0 _0213_
rlabel metal1 8832 17578 8832 17578 0 _0214_
rlabel metal1 23368 14450 23368 14450 0 _0215_
rlabel metal1 23598 15130 23598 15130 0 _0216_
rlabel metal1 7866 13158 7866 13158 0 _0217_
rlabel metal2 24058 14076 24058 14076 0 _0218_
rlabel metal2 14490 23256 14490 23256 0 _0219_
rlabel metal1 10856 23698 10856 23698 0 _0220_
rlabel metal2 15410 19754 15410 19754 0 _0221_
rlabel metal1 17158 18666 17158 18666 0 _0222_
rlabel metal1 7866 23290 7866 23290 0 _0223_
rlabel metal1 16652 17170 16652 17170 0 _0224_
rlabel metal1 21896 22950 21896 22950 0 _0225_
rlabel metal2 28290 21284 28290 21284 0 _0226_
rlabel metal2 20378 20026 20378 20026 0 _0227_
rlabel metal2 22218 21726 22218 21726 0 _0228_
rlabel metal1 28750 22202 28750 22202 0 _0229_
rlabel metal2 21390 20196 21390 20196 0 _0230_
rlabel metal1 20792 17238 20792 17238 0 _0231_
rlabel metal2 30406 17068 30406 17068 0 _0232_
rlabel metal2 16606 18836 16606 18836 0 _0233_
rlabel metal1 14306 17850 14306 17850 0 _0234_
rlabel metal1 30958 15674 30958 15674 0 _0235_
rlabel metal1 22402 17850 22402 17850 0 _0236_
rlabel metal1 25622 16184 25622 16184 0 _0237_
rlabel metal2 25254 14348 25254 14348 0 _0238_
rlabel metal1 21068 18258 21068 18258 0 _0239_
rlabel metal1 25254 18326 25254 18326 0 _0240_
rlabel metal1 24886 12750 24886 12750 0 _0241_
rlabel metal1 24380 18394 24380 18394 0 _0242_
rlabel metal2 7130 21794 7130 21794 0 _0243_
rlabel metal2 10902 21828 10902 21828 0 _0244_
rlabel metal1 4922 19278 4922 19278 0 _0245_
rlabel metal2 5198 19992 5198 19992 0 _0246_
rlabel metal1 13156 20026 13156 20026 0 _0247_
rlabel metal1 4600 18938 4600 18938 0 _0248_
rlabel metal2 28474 8024 28474 8024 0 _0249_
rlabel metal1 28152 17714 28152 17714 0 _0250_
rlabel metal1 30866 6188 30866 6188 0 _0251_
rlabel metal2 27646 6120 27646 6120 0 _0252_
rlabel metal1 27232 17850 27232 17850 0 _0253_
rlabel metal2 30682 3740 30682 3740 0 _0254_
rlabel metal2 12926 18904 12926 18904 0 _0255_
rlabel metal2 12374 23868 12374 23868 0 _0256_
rlabel metal2 24334 26384 24334 26384 0 _0257_
rlabel metal1 12098 18632 12098 18632 0 _0258_
rlabel metal2 13386 24276 13386 24276 0 _0259_
rlabel metal1 17618 27336 17618 27336 0 _0260_
rlabel metal1 26864 26010 26864 26010 0 _0261_
rlabel metal1 26680 26418 26680 26418 0 _0262_
rlabel metal1 25070 27948 25070 27948 0 _0263_
rlabel metal1 26266 27098 26266 27098 0 _0264_
rlabel metal1 27324 24922 27324 24922 0 _0265_
rlabel metal1 29762 27642 29762 27642 0 _0266_
rlabel metal2 15502 25704 15502 25704 0 _0267_
rlabel metal2 12926 25942 12926 25942 0 _0268_
rlabel metal2 22678 23902 22678 23902 0 _0269_
rlabel metal1 16652 22746 16652 22746 0 _0270_
rlabel metal1 16146 22202 16146 22202 0 _0271_
rlabel metal1 9062 22202 9062 22202 0 _0272_
rlabel metal2 24794 10472 24794 10472 0 _0273_
rlabel metal1 28152 8398 28152 8398 0 _0274_
rlabel metal1 9292 17306 9292 17306 0 _0275_
rlabel metal1 7360 16558 7360 16558 0 _0276_
rlabel metal1 24426 8058 24426 8058 0 _0277_
rlabel metal1 6532 17306 6532 17306 0 _0278_
rlabel metal2 21022 26520 21022 26520 0 _0279_
rlabel metal2 16698 26588 16698 26588 0 _0280_
rlabel metal2 25070 10948 25070 10948 0 _0281_
rlabel metal1 23460 22066 23460 22066 0 _0282_
rlabel metal1 14766 26554 14766 26554 0 _0283_
rlabel metal1 23138 12750 23138 12750 0 _0284_
rlabel metal1 29900 10234 29900 10234 0 _0285_
rlabel metal1 30682 19278 30682 19278 0 _0286_
rlabel metal1 15456 24378 15456 24378 0 _0287_
rlabel metal2 28750 9316 28750 9316 0 _0288_
rlabel metal1 28658 20434 28658 20434 0 _0289_
rlabel metal1 24794 8840 24794 8840 0 _0290_
rlabel metal1 15088 29682 15088 29682 0 _0291_
rlabel metal2 19734 30940 19734 30940 0 _0292_
rlabel metal1 24518 20502 24518 20502 0 _0293_
rlabel metal1 15272 29138 15272 29138 0 _0294_
rlabel metal2 19366 29444 19366 29444 0 _0295_
rlabel metal1 23414 30600 23414 30600 0 _0296_
rlabel metal2 9890 21352 9890 21352 0 _0297_
rlabel metal2 13110 21148 13110 21148 0 _0298_
rlabel metal1 18032 22406 18032 22406 0 _0299_
rlabel metal2 9798 19992 9798 19992 0 _0300_
rlabel metal1 16008 18938 16008 18938 0 _0301_
rlabel metal1 5612 22678 5612 22678 0 _0302_
rlabel metal1 23552 25942 23552 25942 0 _0303_
rlabel metal1 11914 25738 11914 25738 0 _0304_
rlabel metal1 19642 25160 19642 25160 0 _0305_
rlabel metal1 15042 21114 15042 21114 0 _0306_
rlabel metal1 20148 26554 20148 26554 0 _0307_
rlabel metal1 30498 8058 30498 8058 0 _0308_
rlabel metal1 22402 19482 22402 19482 0 _0309_
rlabel metal1 30544 12410 30544 12410 0 _0310_
rlabel metal2 30958 13022 30958 13022 0 _0311_
rlabel metal2 9798 25704 9798 25704 0 _0312_
rlabel metal1 27370 17272 27370 17272 0 _0313_
rlabel metal1 16054 24072 16054 24072 0 _0314_
rlabel metal2 32522 11560 32522 11560 0 _0315_
rlabel metal1 5796 17510 5796 17510 0 _0316_
rlabel metal2 13662 18632 13662 18632 0 _0317_
rlabel metal2 4830 17442 4830 17442 0 _0318_
rlabel metal1 18722 27098 18722 27098 0 _0319_
rlabel metal2 30038 15640 30038 15640 0 _0320_
rlabel metal1 18216 23290 18216 23290 0 _0321_
rlabel metal2 22402 20808 22402 20808 0 _0322_
rlabel metal2 16146 26792 16146 26792 0 _0323_
rlabel metal1 31878 13498 31878 13498 0 _0324_
rlabel metal1 17526 20808 17526 20808 0 _0325_
rlabel metal2 28106 11730 28106 11730 0 _0326_
rlabel metal1 30820 3094 30820 3094 0 _0327_
rlabel metal1 27554 3570 27554 3570 0 _0328_
rlabel metal2 28842 3230 28842 3230 0 _0329_
rlabel metal1 24012 5814 24012 5814 0 _0330_
rlabel metal2 25806 4352 25806 4352 0 _0331_
rlabel metal2 28106 4828 28106 4828 0 _0332_
rlabel metal1 24656 4114 24656 4114 0 _0333_
rlabel metal1 18170 6188 18170 6188 0 _0334_
rlabel metal2 28842 6120 28842 6120 0 _0335_
rlabel metal1 19274 15674 19274 15674 0 _0336_
rlabel metal1 25024 4522 25024 4522 0 _0337_
rlabel metal1 9154 16762 9154 16762 0 _0338_
rlabel metal1 14030 27982 14030 27982 0 _0339_
rlabel metal1 20010 21590 20010 21590 0 _0340_
rlabel metal2 12926 28356 12926 28356 0 _0341_
rlabel metal1 20884 24378 20884 24378 0 _0342_
rlabel metal2 8326 21352 8326 21352 0 _0343_
rlabel metal2 27186 19618 27186 19618 0 _0344_
rlabel metal1 15502 20026 15502 20026 0 _0345_
rlabel metal1 28980 20026 28980 20026 0 _0346_
rlabel via1 21482 7429 21482 7429 0 _0347_
rlabel metal2 12006 17816 12006 17816 0 _0348_
rlabel metal2 23690 10200 23690 10200 0 _0349_
rlabel metal1 4462 16422 4462 16422 0 _0350_
rlabel metal1 5566 17034 5566 17034 0 _0351_
rlabel metal1 28658 13498 28658 13498 0 _0352_
rlabel metal2 22218 7582 22218 7582 0 _0353_
rlabel metal1 29026 6834 29026 6834 0 _0354_
rlabel metal1 27646 3026 27646 3026 0 _0355_
rlabel metal1 12052 16966 12052 16966 0 _0356_
rlabel metal2 24150 3196 24150 3196 0 _0357_
rlabel metal2 23506 3706 23506 3706 0 _0358_
rlabel metal1 12006 21658 12006 21658 0 _0359_
rlabel metal1 24242 5882 24242 5882 0 _0360_
rlabel metal2 12190 19074 12190 19074 0 _0361_
rlabel metal2 22218 3502 22218 3502 0 _0362_
rlabel metal2 12006 30056 12006 30056 0 _0363_
rlabel metal2 8234 28628 8234 28628 0 _0364_
rlabel metal1 10120 29274 10120 29274 0 _0365_
rlabel metal2 7314 29988 7314 29988 0 _0366_
rlabel metal2 38318 6239 38318 6239 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 38318 33439 38318 33439 0 bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 22770 37230 22770 37230 0 bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 37490 37723 37490 37723 0 bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal3 1234 12308 1234 12308 0 bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal2 34822 1588 34822 1588 0 bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_
rlabel metal3 1740 36788 1740 36788 0 bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal1 38180 36142 38180 36142 0 bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_
rlabel metal2 29026 1554 29026 1554 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
rlabel metal2 2806 7701 2806 7701 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
rlabel metal3 1142 30668 1142 30668 0 ccff_head
rlabel metal2 10350 1520 10350 1520 0 ccff_tail
rlabel metal3 1924 38148 1924 38148 0 chanx_right_in[0]
rlabel metal2 4554 1520 4554 1520 0 chanx_right_in[10]
rlabel metal3 1234 20468 1234 20468 0 chanx_right_in[11]
rlabel metal3 1234 17748 1234 17748 0 chanx_right_in[12]
rlabel metal2 38318 28883 38318 28883 0 chanx_right_in[13]
rlabel metal1 18216 37230 18216 37230 0 chanx_right_in[14]
rlabel metal2 33534 1588 33534 1588 0 chanx_right_in[15]
rlabel metal3 1234 25228 1234 25228 0 chanx_right_in[16]
rlabel metal3 1234 32028 1234 32028 0 chanx_right_in[17]
rlabel metal3 1234 27268 1234 27268 0 chanx_right_in[18]
rlabel metal2 22586 1554 22586 1554 0 chanx_right_in[1]
rlabel metal2 14858 1588 14858 1588 0 chanx_right_in[2]
rlabel metal2 39330 1860 39330 1860 0 chanx_right_in[3]
rlabel metal3 1740 1428 1740 1428 0 chanx_right_in[4]
rlabel metal2 38318 20689 38318 20689 0 chanx_right_in[5]
rlabel metal1 24656 37230 24656 37230 0 chanx_right_in[6]
rlabel metal1 14030 37230 14030 37230 0 chanx_right_in[7]
rlabel via2 36938 36771 36938 36771 0 chanx_right_in[8]
rlabel metal2 16790 1588 16790 1588 0 chanx_right_in[9]
rlabel metal3 1234 15708 1234 15708 0 chanx_right_out[0]
rlabel metal2 38226 34833 38226 34833 0 chanx_right_out[10]
rlabel metal1 15640 37094 15640 37094 0 chanx_right_out[11]
rlabel metal2 38226 8857 38226 8857 0 chanx_right_out[12]
rlabel metal2 38226 12461 38226 12461 0 chanx_right_out[13]
rlabel metal1 16928 37094 16928 37094 0 chanx_right_out[14]
rlabel metal1 10488 37094 10488 37094 0 chanx_right_out[15]
rlabel metal2 25806 823 25806 823 0 chanx_right_out[16]
rlabel metal2 9062 1520 9062 1520 0 chanx_right_out[17]
rlabel via2 38226 30005 38226 30005 0 chanx_right_out[18]
rlabel metal2 38042 1520 38042 1520 0 chanx_right_out[1]
rlabel metal2 38226 15793 38226 15793 0 chanx_right_out[2]
rlabel metal1 29486 37094 29486 37094 0 chanx_right_out[3]
rlabel metal1 12512 37094 12512 37094 0 chanx_right_out[4]
rlabel metal2 38226 2125 38226 2125 0 chanx_right_out[5]
rlabel metal2 38226 32113 38226 32113 0 chanx_right_out[6]
rlabel metal1 36800 37094 36800 37094 0 chanx_right_out[7]
rlabel metal1 21758 37094 21758 37094 0 chanx_right_out[8]
rlabel metal3 1234 19108 1234 19108 0 chanx_right_out[9]
rlabel metal2 38318 7701 38318 7701 0 chany_bottom_in[0]
rlabel metal3 1234 22508 1234 22508 0 chany_bottom_in[10]
rlabel metal3 1234 2788 1234 2788 0 chany_bottom_in[11]
rlabel metal1 25944 37230 25944 37230 0 chany_bottom_in[12]
rlabel metal3 1234 28628 1234 28628 0 chany_bottom_in[13]
rlabel metal2 31786 2652 31786 2652 0 chany_bottom_in[14]
rlabel metal1 33672 37230 33672 37230 0 chany_bottom_in[15]
rlabel metal3 1234 9588 1234 9588 0 chany_bottom_in[16]
rlabel metal2 2622 1588 2622 1588 0 chany_bottom_in[17]
rlabel metal2 11638 1588 11638 1588 0 chany_bottom_in[18]
rlabel metal2 36110 1588 36110 1588 0 chany_bottom_in[1]
rlabel metal2 38318 17119 38318 17119 0 chany_bottom_in[2]
rlabel metal2 38318 11033 38318 11033 0 chany_bottom_in[3]
rlabel metal3 1234 6188 1234 6188 0 chany_bottom_in[4]
rlabel metal3 1234 33388 1234 33388 0 chany_bottom_in[5]
rlabel metal2 38318 3145 38318 3145 0 chany_bottom_in[6]
rlabel metal1 4738 37230 4738 37230 0 chany_bottom_in[7]
rlabel via2 38318 14365 38318 14365 0 chany_bottom_in[8]
rlabel via2 38318 25245 38318 25245 0 chany_bottom_in[9]
rlabel metal2 31602 1520 31602 1520 0 chany_bottom_out[0]
rlabel via2 38226 27285 38226 27285 0 chany_bottom_out[10]
rlabel metal1 6302 37094 6302 37094 0 chany_bottom_out[11]
rlabel metal3 1234 23868 1234 23868 0 chany_bottom_out[12]
rlabel metal2 19366 1520 19366 1520 0 chany_bottom_out[13]
rlabel metal2 46 1792 46 1792 0 chany_bottom_out[14]
rlabel metal2 23874 1520 23874 1520 0 chany_bottom_out[15]
rlabel metal1 7912 37094 7912 37094 0 chany_bottom_out[16]
rlabel metal1 20148 37094 20148 37094 0 chany_bottom_out[17]
rlabel metal3 1234 4828 1234 4828 0 chany_bottom_out[18]
rlabel metal1 920 36890 920 36890 0 chany_bottom_out[1]
rlabel metal2 5842 1520 5842 1520 0 chany_bottom_out[2]
rlabel metal2 1334 1520 1334 1520 0 chany_bottom_out[3]
rlabel metal1 34960 37094 34960 37094 0 chany_bottom_out[4]
rlabel metal1 27876 37094 27876 37094 0 chany_bottom_out[5]
rlabel metal2 18078 1520 18078 1520 0 chany_bottom_out[6]
rlabel metal1 38778 36890 38778 36890 0 chany_bottom_out[7]
rlabel metal2 38226 4301 38226 4301 0 chany_bottom_out[8]
rlabel metal1 1564 37094 1564 37094 0 chany_bottom_out[9]
rlabel metal2 20838 13940 20838 13940 0 mem_bottom_track_1.DFFR_0_.D
rlabel metal2 13018 16932 13018 16932 0 mem_bottom_track_1.DFFR_0_.Q
rlabel metal2 14030 4522 14030 4522 0 mem_bottom_track_1.DFFR_1_.Q
rlabel metal1 18298 14790 18298 14790 0 mem_bottom_track_11.DFFR_0_.D
rlabel metal2 13386 14756 13386 14756 0 mem_bottom_track_11.DFFR_0_.Q
rlabel metal2 16146 22372 16146 22372 0 mem_bottom_track_11.DFFR_1_.Q
rlabel metal1 5934 17170 5934 17170 0 mem_bottom_track_13.DFFR_0_.Q
rlabel metal2 17250 12206 17250 12206 0 mem_bottom_track_13.DFFR_1_.Q
rlabel metal2 14950 15028 14950 15028 0 mem_bottom_track_15.DFFR_0_.Q
rlabel metal1 18446 11662 18446 11662 0 mem_bottom_track_15.DFFR_1_.Q
rlabel metal1 19504 22066 19504 22066 0 mem_bottom_track_17.DFFR_0_.Q
rlabel metal2 16882 8738 16882 8738 0 mem_bottom_track_17.DFFR_1_.Q
rlabel metal2 19274 29682 19274 29682 0 mem_bottom_track_19.DFFR_0_.Q
rlabel metal1 14766 15130 14766 15130 0 mem_bottom_track_19.DFFR_1_.Q
rlabel metal1 18170 10574 18170 10574 0 mem_bottom_track_23.DFFR_0_.Q
rlabel metal1 13931 13702 13931 13702 0 mem_bottom_track_23.DFFR_1_.Q
rlabel metal2 18722 15929 18722 15929 0 mem_bottom_track_25.DFFR_0_.Q
rlabel metal1 15824 19822 15824 19822 0 mem_bottom_track_25.DFFR_1_.Q
rlabel metal1 8924 2618 8924 2618 0 mem_bottom_track_27.DFFR_0_.Q
rlabel metal1 9522 2074 9522 2074 0 mem_bottom_track_27.DFFR_1_.Q
rlabel metal1 17986 4046 17986 4046 0 mem_bottom_track_29.DFFR_0_.Q
rlabel metal2 13570 13634 13570 13634 0 mem_bottom_track_29.DFFR_1_.Q
rlabel metal1 5796 17646 5796 17646 0 mem_bottom_track_3.DFFR_0_.Q
rlabel metal1 7452 20910 7452 20910 0 mem_bottom_track_3.DFFR_1_.Q
rlabel metal1 19320 3162 19320 3162 0 mem_bottom_track_31.DFFR_0_.Q
rlabel metal2 24610 3417 24610 3417 0 mem_bottom_track_31.DFFR_1_.Q
rlabel metal2 17250 4352 17250 4352 0 mem_bottom_track_33.DFFR_0_.Q
rlabel metal2 12098 17527 12098 17527 0 mem_bottom_track_33.DFFR_1_.Q
rlabel metal1 7866 29614 7866 29614 0 mem_bottom_track_35.DFFR_0_.Q
rlabel metal1 10626 29138 10626 29138 0 mem_bottom_track_35.DFFR_1_.Q
rlabel metal2 14858 18938 14858 18938 0 mem_bottom_track_37.DFFR_0_.Q
rlabel metal1 14536 4522 14536 4522 0 mem_bottom_track_5.DFFR_0_.Q
rlabel metal1 19083 5882 19083 5882 0 mem_bottom_track_5.DFFR_1_.Q
rlabel via2 18170 5627 18170 5627 0 mem_bottom_track_7.DFFR_0_.Q
rlabel metal1 11592 15402 11592 15402 0 mem_bottom_track_7.DFFR_1_.Q
rlabel metal1 13938 15538 13938 15538 0 mem_bottom_track_9.DFFR_0_.Q
rlabel metal1 12834 7752 12834 7752 0 mem_right_track_0.DFFR_0_.Q
rlabel metal1 10672 14382 10672 14382 0 mem_right_track_0.DFFR_1_.Q
rlabel metal1 11638 26962 11638 26962 0 mem_right_track_10.DFFR_0_.D
rlabel metal2 13478 14212 13478 14212 0 mem_right_track_10.DFFR_0_.Q
rlabel metal2 14398 10268 14398 10268 0 mem_right_track_10.DFFR_1_.Q
rlabel via2 12650 12597 12650 12597 0 mem_right_track_12.DFFR_0_.Q
rlabel metal2 17066 11356 17066 11356 0 mem_right_track_12.DFFR_1_.Q
rlabel metal2 11730 24276 11730 24276 0 mem_right_track_14.DFFR_0_.Q
rlabel metal1 14306 19754 14306 19754 0 mem_right_track_14.DFFR_1_.Q
rlabel metal1 17250 15402 17250 15402 0 mem_right_track_16.DFFR_0_.Q
rlabel metal1 20976 21998 20976 21998 0 mem_right_track_16.DFFR_1_.Q
rlabel metal1 14536 16694 14536 16694 0 mem_right_track_18.DFFR_0_.Q
rlabel metal1 14076 17646 14076 17646 0 mem_right_track_18.DFFR_1_.Q
rlabel metal2 18722 16354 18722 16354 0 mem_right_track_2.DFFR_0_.Q
rlabel metal2 18262 7038 18262 7038 0 mem_right_track_2.DFFR_1_.Q
rlabel metal1 12742 20910 12742 20910 0 mem_right_track_20.DFFR_0_.Q
rlabel metal2 17986 16252 17986 16252 0 mem_right_track_20.DFFR_1_.Q
rlabel metal1 14204 13498 14204 13498 0 mem_right_track_22.DFFR_0_.Q
rlabel metal2 20654 17017 20654 17017 0 mem_right_track_22.DFFR_1_.Q
rlabel metal1 10994 24174 10994 24174 0 mem_right_track_24.DFFR_0_.Q
rlabel metal1 15778 12852 15778 12852 0 mem_right_track_24.DFFR_1_.Q
rlabel metal1 5244 16082 5244 16082 0 mem_right_track_26.DFFR_0_.Q
rlabel metal1 13570 17578 13570 17578 0 mem_right_track_26.DFFR_1_.Q
rlabel metal1 18860 9486 18860 9486 0 mem_right_track_28.DFFR_0_.Q
rlabel metal2 20516 17204 20516 17204 0 mem_right_track_28.DFFR_1_.Q
rlabel metal2 31878 11696 31878 11696 0 mem_right_track_30.DFFR_0_.Q
rlabel metal2 19458 20740 19458 20740 0 mem_right_track_30.DFFR_1_.Q
rlabel metal1 14582 3910 14582 3910 0 mem_right_track_32.DFFR_0_.Q
rlabel metal2 7866 5032 7866 5032 0 mem_right_track_32.DFFR_1_.Q
rlabel metal1 14306 5304 14306 5304 0 mem_right_track_34.DFFR_0_.Q
rlabel metal2 15778 3944 15778 3944 0 mem_right_track_34.DFFR_1_.Q
rlabel metal1 22034 17680 22034 17680 0 mem_right_track_36.DFFR_0_.Q
rlabel metal1 19964 7310 19964 7310 0 mem_right_track_4.DFFR_0_.Q
rlabel metal1 14076 12750 14076 12750 0 mem_right_track_4.DFFR_1_.Q
rlabel metal2 33258 14416 33258 14416 0 mem_right_track_6.DFFR_0_.Q
rlabel metal2 16238 18258 16238 18258 0 mem_right_track_6.DFFR_1_.Q
rlabel metal2 6762 27234 6762 27234 0 mem_right_track_8.DFFR_0_.Q
rlabel metal1 8050 24582 8050 24582 0 mux_bottom_track_1.INVTX1_0_.out
rlabel metal1 19826 17544 19826 17544 0 mux_bottom_track_1.INVTX1_1_.out
rlabel metal1 19458 17714 19458 17714 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 29762 6358 29762 6358 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 31510 2618 31510 2618 0 mux_bottom_track_1.out
rlabel metal1 7406 22542 7406 22542 0 mux_bottom_track_11.INVTX1_0_.out
rlabel metal1 28566 16014 28566 16014 0 mux_bottom_track_11.INVTX1_1_.out
rlabel metal1 15870 23018 15870 23018 0 mux_bottom_track_11.INVTX1_2_.out
rlabel metal2 9430 22950 9430 22950 0 mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 15870 25806 15870 25806 0 mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 16376 25874 16376 25874 0 mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 25530 29818 25530 29818 0 mux_bottom_track_11.out
rlabel metal1 6256 18394 6256 18394 0 mux_bottom_track_13.INVTX1_0_.out
rlabel metal1 23138 6188 23138 6188 0 mux_bottom_track_13.INVTX1_2_.out
rlabel metal1 9752 18190 9752 18190 0 mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 25070 9214 25070 9214 0 mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 21942 9503 21942 9503 0 mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel via1 18722 3500 18722 3500 0 mux_bottom_track_13.out
rlabel metal1 18400 13158 18400 13158 0 mux_bottom_track_15.INVTX1_0_.out
rlabel metal2 8050 28866 8050 28866 0 mux_bottom_track_15.INVTX1_2_.out
rlabel metal2 25484 16116 25484 16116 0 mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 19044 26418 19044 26418 0 mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 24794 28322 24794 28322 0 mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 32982 31586 32982 31586 0 mux_bottom_track_15.out
rlabel metal1 23414 2618 23414 2618 0 mux_bottom_track_17.INVTX1_0_.out
rlabel metal1 18883 20434 18883 20434 0 mux_bottom_track_17.INVTX1_2_.out
rlabel metal1 15732 8602 15732 8602 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 30314 19346 30314 19346 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 30590 9690 30590 9690 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 32522 8636 32522 8636 0 mux_bottom_track_17.out
rlabel metal1 28796 31858 28796 31858 0 mux_bottom_track_19.INVTX1_0_.out
rlabel metal1 14490 29172 14490 29172 0 mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 19274 29750 19274 29750 0 mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 14628 29818 14628 29818 0 mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 10672 35054 10672 35054 0 mux_bottom_track_19.out
rlabel metal2 23230 29002 23230 29002 0 mux_bottom_track_23.INVTX1_0_.out
rlabel metal2 19826 21114 19826 21114 0 mux_bottom_track_23.INVTX1_1_.out
rlabel metal1 20562 21590 20562 21590 0 mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 12788 28730 12788 28730 0 mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 12328 32878 12328 32878 0 mux_bottom_track_23.out
rlabel metal2 30774 20196 30774 20196 0 mux_bottom_track_25.INVTX1_0_.out
rlabel metal1 27324 19890 27324 19890 0 mux_bottom_track_25.INVTX1_1_.out
rlabel metal1 18630 20910 18630 20910 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 14053 21046 14053 21046 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 8280 23698 8280 23698 0 mux_bottom_track_25.out
rlabel metal2 6118 8738 6118 8738 0 mux_bottom_track_27.INVTX1_0_.out
rlabel metal1 13248 24786 13248 24786 0 mux_bottom_track_27.INVTX1_1_.out
rlabel metal2 13662 10200 13662 10200 0 mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 21574 4811 21574 4811 0 mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 17066 4250 17066 4250 0 mux_bottom_track_27.out
rlabel metal1 29486 5338 29486 5338 0 mux_bottom_track_29.INVTX1_0_.out
rlabel metal1 29210 16014 29210 16014 0 mux_bottom_track_29.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 2346 5270 2346 5270 0 mux_bottom_track_29.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 2530 4012 2530 4012 0 mux_bottom_track_29.out
rlabel metal1 3036 20434 3036 20434 0 mux_bottom_track_3.INVTX1_0_.out
rlabel metal2 3450 16694 3450 16694 0 mux_bottom_track_3.INVTX1_1_.out
rlabel metal2 5106 20060 5106 20060 0 mux_bottom_track_3.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 11500 21862 11500 21862 0 mux_bottom_track_3.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 4186 24140 4186 24140 0 mux_bottom_track_3.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 4462 24378 4462 24378 0 mux_bottom_track_3.out
rlabel metal1 23368 3162 23368 3162 0 mux_bottom_track_31.INVTX1_0_.out
rlabel metal2 14950 10472 14950 10472 0 mux_bottom_track_31.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 25070 3094 25070 3094 0 mux_bottom_track_31.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 25668 3094 25668 3094 0 mux_bottom_track_31.out
rlabel metal1 22172 2618 22172 2618 0 mux_bottom_track_33.INVTX1_0_.out
rlabel metal2 10534 18768 10534 18768 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 12052 22542 12052 22542 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 10626 31042 10626 31042 0 mux_bottom_track_33.out
rlabel metal2 5198 29988 5198 29988 0 mux_bottom_track_35.INVTX1_0_.out
rlabel metal2 8694 29648 8694 29648 0 mux_bottom_track_35.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 14674 29750 14674 29750 0 mux_bottom_track_35.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 17342 32402 17342 32402 0 mux_bottom_track_35.out
rlabel metal2 5382 23630 5382 23630 0 mux_bottom_track_37.INVTX1_0_.out
rlabel metal1 7038 22474 7038 22474 0 mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 14628 20298 14628 20298 0 mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 8694 18224 8694 18224 0 mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 2898 15130 2898 15130 0 mux_bottom_track_37.out
rlabel metal1 30498 3468 30498 3468 0 mux_bottom_track_5.INVTX1_0_.out
rlabel metal1 29302 6426 29302 6426 0 mux_bottom_track_5.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 28336 17782 28336 17782 0 mux_bottom_track_5.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 27830 4828 27830 4828 0 mux_bottom_track_5.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 3358 2975 3358 2975 0 mux_bottom_track_5.out
rlabel metal2 17526 27234 17526 27234 0 mux_bottom_track_7.INVTX1_0_.out
rlabel metal2 18170 24725 18170 24725 0 mux_bottom_track_7.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 12834 24208 12834 24208 0 mux_bottom_track_7.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 2254 6800 2254 6800 0 mux_bottom_track_7.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 2668 6766 2668 6766 0 mux_bottom_track_7.out
rlabel metal2 29486 28220 29486 28220 0 mux_bottom_track_9.INVTX1_0_.out
rlabel metal1 26864 27506 26864 27506 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 27048 26350 27048 26350 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 27830 26928 27830 26928 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 30590 34510 30590 34510 0 mux_bottom_track_9.out
rlabel metal2 19274 18972 19274 18972 0 mux_right_track_0.INVTX1_0_.out
rlabel metal1 17756 19890 17756 19890 0 mux_right_track_0.INVTX1_1_.out
rlabel metal1 2254 17102 2254 17102 0 mux_right_track_0.INVTX1_2_.out
rlabel metal1 17710 19754 17710 19754 0 mux_right_track_0.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 4646 15130 4646 15130 0 mux_right_track_0.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 1886 12240 1886 12240 0 mux_right_track_0.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 1978 13158 1978 13158 0 mux_right_track_0.out
rlabel metal2 9890 27812 9890 27812 0 mux_right_track_10.INVTX1_0_.out
rlabel metal1 27186 13940 27186 13940 0 mux_right_track_10.INVTX1_1_.out
rlabel metal2 25070 26044 25070 26044 0 mux_right_track_10.INVTX1_2_.out
rlabel metal1 28106 13838 28106 13838 0 mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 28106 15062 28106 15062 0 mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 29532 13838 29532 13838 0 mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 31234 6188 31234 6188 0 mux_right_track_10.out
rlabel metal2 21482 17136 21482 17136 0 mux_right_track_12.INVTX1_1_.out
rlabel metal2 6026 8398 6026 8398 0 mux_right_track_12.INVTX1_2_.out
rlabel metal1 23644 14586 23644 14586 0 mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 16790 17034 16790 17034 0 mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 32890 27404 32890 27404 0 mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 33074 27574 33074 27574 0 mux_right_track_12.out
rlabel metal1 18676 20366 18676 20366 0 mux_right_track_14.INVTX1_1_.out
rlabel metal1 6992 24174 6992 24174 0 mux_right_track_14.INVTX1_2_.out
rlabel metal1 17158 18802 17158 18802 0 mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 9706 23834 9706 23834 0 mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 18400 18802 18400 18802 0 mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 31464 33082 31464 33082 0 mux_right_track_14.out
rlabel metal2 16422 18190 16422 18190 0 mux_right_track_16.INVTX1_1_.out
rlabel metal2 28474 23324 28474 23324 0 mux_right_track_16.INVTX1_2_.out
rlabel metal2 21206 19856 21206 19856 0 mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 22034 21794 22034 21794 0 mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 21850 21726 21850 21726 0 mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 21022 29308 21022 29308 0 mux_right_track_16.out
rlabel metal2 33534 15776 33534 15776 0 mux_right_track_18.INVTX1_2_.out
rlabel metal1 17112 17850 17112 17850 0 mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 30590 16864 30590 16864 0 mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 14812 18190 14812 18190 0 mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 7314 18972 7314 18972 0 mux_right_track_18.out
rlabel metal2 31878 18190 31878 18190 0 mux_right_track_2.INVTX1_1_.out
rlabel metal2 8602 8602 8602 8602 0 mux_right_track_2.INVTX1_2_.out
rlabel metal1 26404 13430 26404 13430 0 mux_right_track_2.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 18906 18156 18906 18156 0 mux_right_track_2.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 26542 6800 26542 6800 0 mux_right_track_2.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 30590 5168 30590 5168 0 mux_right_track_2.out
rlabel metal1 11270 28390 11270 28390 0 mux_right_track_20.INVTX1_1_.out
rlabel metal1 17664 22066 17664 22066 0 mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 23874 25874 23874 25874 0 mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 33626 29478 33626 29478 0 mux_right_track_20.out
rlabel metal2 31786 8228 31786 8228 0 mux_right_track_22.INVTX1_1_.out
rlabel metal1 30820 13430 30820 13430 0 mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 20056 29138 20056 29138 0 mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 20010 29988 20010 29988 0 mux_right_track_22.out
rlabel metal2 28290 25228 28290 25228 0 mux_right_track_24.INVTX1_0_.out
rlabel metal1 8142 27370 8142 27370 0 mux_right_track_24.INVTX1_1_.out
rlabel metal1 11822 25840 11822 25840 0 mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 31142 14892 31142 14892 0 mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 33534 10642 33534 10642 0 mux_right_track_24.out
rlabel metal2 6854 27744 6854 27744 0 mux_right_track_26.INVTX1_0_.out
rlabel metal1 3680 10574 3680 10574 0 mux_right_track_26.INVTX1_1_.out
rlabel metal2 14122 19618 14122 19618 0 mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 33028 12206 33028 12206 0 mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 34730 12206 34730 12206 0 mux_right_track_26.out
rlabel metal2 31050 14790 31050 14790 0 mux_right_track_28.INVTX1_1_.out
rlabel metal1 18262 24276 18262 24276 0 mux_right_track_28.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 18860 29546 18860 29546 0 mux_right_track_28.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 17250 30906 17250 30906 0 mux_right_track_28.out
rlabel metal2 32890 14892 32890 14892 0 mux_right_track_30.INVTX1_1_.out
rlabel metal2 31970 13328 31970 13328 0 mux_right_track_30.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 17802 21046 17802 21046 0 mux_right_track_30.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 14720 30362 14720 30362 0 mux_right_track_30.out
rlabel metal1 25714 2618 25714 2618 0 mux_right_track_32.INVTX1_1_.out
rlabel metal1 25806 3706 25806 3706 0 mux_right_track_32.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 29026 2924 29026 2924 0 mux_right_track_32.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 27600 2346 27600 2346 0 mux_right_track_32.out
rlabel metal2 27922 4420 27922 4420 0 mux_right_track_34.INVTX1_1_.out
rlabel metal2 18630 5950 18630 5950 0 mux_right_track_34.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 24840 4726 24840 4726 0 mux_right_track_34.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 7774 2176 7774 2176 0 mux_right_track_34.out
rlabel metal1 25622 12818 25622 12818 0 mux_right_track_36.INVTX1_2_.out
rlabel metal1 24932 18598 24932 18598 0 mux_right_track_36.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 25622 14042 25622 14042 0 mux_right_track_36.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 25622 18190 25622 18190 0 mux_right_track_36.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 33534 23868 33534 23868 0 mux_right_track_36.out
rlabel metal1 32614 30566 32614 30566 0 mux_right_track_4.INVTX1_2_.out
rlabel metal1 29532 23222 29532 23222 0 mux_right_track_4.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 31970 23834 31970 23834 0 mux_right_track_4.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 30406 22304 30406 22304 0 mux_right_track_4.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 31510 18428 31510 18428 0 mux_right_track_4.out
rlabel metal1 29072 4114 29072 4114 0 mux_right_track_6.INVTX1_2_.out
rlabel metal2 20838 25534 20838 25534 0 mux_right_track_6.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 32660 17102 32660 17102 0 mux_right_track_6.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 26358 20985 26358 20985 0 mux_right_track_6.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 28520 29818 28520 29818 0 mux_right_track_6.out
rlabel metal2 5842 27132 5842 27132 0 mux_right_track_8.INVTX1_2_.out
rlabel metal1 10166 27540 10166 27540 0 mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 7866 26010 7866 26010 0 mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 10810 28526 10810 28526 0 mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 11592 29818 11592 29818 0 mux_right_track_8.out
rlabel metal2 38134 5882 38134 5882 0 net1
rlabel metal1 2530 8058 2530 8058 0 net10
rlabel metal1 3634 17646 3634 17646 0 net100
rlabel metal1 18676 17714 18676 17714 0 net101
rlabel metal1 30820 23630 30820 23630 0 net102
rlabel metal2 32430 17374 32430 17374 0 net103
rlabel metal2 7314 26044 7314 26044 0 net104
rlabel metal1 25852 22066 25852 22066 0 net105
rlabel metal2 9246 18156 9246 18156 0 net106
rlabel metal2 10534 23868 10534 23868 0 net107
rlabel metal2 28106 21692 28106 21692 0 net108
rlabel metal2 30222 16864 30222 16864 0 net109
rlabel metal2 1886 21692 1886 21692 0 net11
rlabel metal1 25116 13362 25116 13362 0 net110
rlabel metal1 10212 22542 10212 22542 0 net111
rlabel metal1 28566 17646 28566 17646 0 net112
rlabel metal2 12190 23392 12190 23392 0 net113
rlabel metal2 25990 26656 25990 26656 0 net114
rlabel metal2 12742 25568 12742 25568 0 net115
rlabel metal2 27186 8636 27186 8636 0 net116
rlabel metal2 16514 26656 16514 26656 0 net117
rlabel metal1 29900 18802 29900 18802 0 net118
rlabel metal2 19550 31008 19550 31008 0 net119
rlabel metal1 4048 29614 4048 29614 0 net12
rlabel metal1 12236 20366 12236 20366 0 net120
rlabel metal2 23046 26078 23046 26078 0 net121
rlabel metal1 19642 28152 19642 28152 0 net122
rlabel metal1 30912 12274 30912 12274 0 net123
rlabel metal2 32430 11934 32430 11934 0 net124
rlabel metal2 18170 29410 18170 29410 0 net125
rlabel metal2 14490 28254 14490 28254 0 net126
rlabel metal1 30360 2958 30360 2958 0 net127
rlabel metal2 23414 4896 23414 4896 0 net128
rlabel metal2 28198 5984 28198 5984 0 net129
rlabel metal1 5336 2618 5336 2618 0 net13
rlabel metal1 12696 27506 12696 27506 0 net130
rlabel metal2 7958 21216 7958 21216 0 net131
rlabel metal2 20930 5916 20930 5916 0 net132
rlabel metal2 6762 10846 6762 10846 0 net133
rlabel metal1 27186 3060 27186 3060 0 net134
rlabel metal1 11684 22066 11684 22066 0 net135
rlabel metal2 11914 29410 11914 29410 0 net136
rlabel metal2 5382 19516 5382 19516 0 net14
rlabel metal2 3818 19652 3818 19652 0 net15
rlabel metal2 34546 28764 34546 28764 0 net16
rlabel metal1 18078 37094 18078 37094 0 net17
rlabel metal2 33718 3060 33718 3060 0 net18
rlabel metal2 3174 23868 3174 23868 0 net19
rlabel metal2 38134 29376 38134 29376 0 net2
rlabel metal1 3956 32198 3956 32198 0 net20
rlabel metal1 3496 27302 3496 27302 0 net21
rlabel metal1 22402 2448 22402 2448 0 net22
rlabel metal2 16698 2414 16698 2414 0 net23
rlabel metal2 36754 4216 36754 4216 0 net24
rlabel metal1 1656 3978 1656 3978 0 net25
rlabel metal2 34546 20332 34546 20332 0 net26
rlabel metal1 23874 37094 23874 37094 0 net27
rlabel metal1 21390 31858 21390 31858 0 net28
rlabel metal2 36754 34170 36754 34170 0 net29
rlabel metal1 22402 28050 22402 28050 0 net3
rlabel metal1 22724 2414 22724 2414 0 net30
rlabel metal1 37720 7718 37720 7718 0 net31
rlabel metal1 3726 22474 3726 22474 0 net32
rlabel metal1 1748 3706 1748 3706 0 net33
rlabel metal1 25530 37094 25530 37094 0 net34
rlabel metal2 5750 28220 5750 28220 0 net35
rlabel metal1 32384 2550 32384 2550 0 net36
rlabel metal1 33488 37094 33488 37094 0 net37
rlabel metal2 1886 9418 1886 9418 0 net38
rlabel metal1 2530 2618 2530 2618 0 net39
rlabel metal2 37766 31790 37766 31790 0 net4
rlabel metal2 11730 2142 11730 2142 0 net40
rlabel metal1 26082 2380 26082 2380 0 net41
rlabel metal1 37030 16966 37030 16966 0 net42
rlabel metal2 38134 12614 38134 12614 0 net43
rlabel metal1 1748 10642 1748 10642 0 net44
rlabel metal2 7222 30362 7222 30362 0 net45
rlabel metal1 35604 3706 35604 3706 0 net46
rlabel metal2 4646 36992 4646 36992 0 net47
rlabel metal2 34638 15028 34638 15028 0 net48
rlabel metal2 38134 24684 38134 24684 0 net49
rlabel metal2 1610 13124 1610 13124 0 net5
rlabel metal2 37766 15708 37766 15708 0 net50
rlabel metal1 14674 2618 14674 2618 0 net51
rlabel metal2 5106 16762 5106 16762 0 net52
rlabel metal2 37030 23562 37030 23562 0 net53
rlabel metal1 21252 2278 21252 2278 0 net54
rlabel metal1 32384 37094 32384 37094 0 net55
rlabel metal1 29716 37162 29716 37162 0 net56
rlabel metal2 4002 32572 4002 32572 0 net57
rlabel metal1 9062 37094 9062 37094 0 net58
rlabel metal1 28520 4522 28520 4522 0 net59
rlabel metal1 34040 2550 34040 2550 0 net6
rlabel metal1 1794 11254 1794 11254 0 net60
rlabel metal1 10212 19346 10212 19346 0 net61
rlabel metal1 1702 14042 1702 14042 0 net62
rlabel metal2 33442 32572 33442 32572 0 net63
rlabel metal2 15594 37060 15594 37060 0 net64
rlabel metal2 34822 9690 34822 9690 0 net65
rlabel metal2 36754 12614 36754 12614 0 net66
rlabel metal2 16882 34612 16882 34612 0 net67
rlabel metal1 12098 37162 12098 37162 0 net68
rlabel metal1 27554 2414 27554 2414 0 net69
rlabel metal2 2346 36958 2346 36958 0 net7
rlabel metal1 9154 2380 9154 2380 0 net70
rlabel metal1 36961 30226 36961 30226 0 net71
rlabel metal1 38042 2448 38042 2448 0 net72
rlabel metal1 36961 16082 36961 16082 0 net73
rlabel metal1 29210 37230 29210 37230 0 net74
rlabel metal1 12052 37230 12052 37230 0 net75
rlabel metal1 38042 3060 38042 3060 0 net76
rlabel metal2 35466 30294 35466 30294 0 net77
rlabel metal1 36271 37230 36271 37230 0 net78
rlabel metal1 21436 29274 21436 29274 0 net79
rlabel metal1 37720 36006 37720 36006 0 net8
rlabel metal1 1610 19380 1610 19380 0 net80
rlabel metal2 32338 2618 32338 2618 0 net81
rlabel metal1 36961 27438 36961 27438 0 net82
rlabel metal1 6739 37230 6739 37230 0 net83
rlabel metal2 1610 24004 1610 24004 0 net84
rlabel viali 19458 2415 19458 2415 0 net85
rlabel metal1 1978 3026 1978 3026 0 net86
rlabel metal1 25024 2414 25024 2414 0 net87
rlabel metal1 8924 31994 8924 31994 0 net88
rlabel metal1 18814 37162 18814 37162 0 net89
rlabel metal1 29256 2278 29256 2278 0 net9
rlabel metal1 1564 5202 1564 5202 0 net90
rlabel metal1 3128 36754 3128 36754 0 net91
rlabel metal1 6210 2414 6210 2414 0 net92
rlabel metal1 2254 2482 2254 2482 0 net93
rlabel metal1 34408 37230 34408 37230 0 net94
rlabel metal1 26910 31450 26910 31450 0 net95
rlabel metal1 18354 3366 18354 3366 0 net96
rlabel metal1 37536 36754 37536 36754 0 net97
rlabel metal1 36248 4590 36248 4590 0 net98
rlabel metal1 2852 37162 2852 37162 0 net99
rlabel metal2 37490 21913 37490 21913 0 pReset
rlabel metal1 18032 14994 18032 14994 0 prog_clk
rlabel metal2 13570 1588 13570 1588 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel metal3 1234 14348 1234 14348 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal2 38318 24021 38318 24021 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 21298 1588 21298 1588 0 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 32384 37230 32384 37230 0 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 30544 37230 30544 37230 0 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 3726 37230 3726 37230 0 right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal1 9200 37230 9200 37230 0 right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_
rlabel metal2 27094 1095 27094 1095 0 right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal3 1234 10948 1234 10948 0 right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
